module TauswortheUniform(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h2ec82d18 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h3536544e : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'hf64f2de : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_1(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h26ce5c2f : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h28cb727d : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h13c77c0e : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Trigonometric(
  input         clock,
  input         reset,
  input         io_theta_valid,
  input  [31:0] io_theta_bits,
  output        io_result_valid,
  output [31:0] io_result_bits_sine,
  output [31:0] io_result_bits_cosine
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
`endif // RANDOMIZE_REG_INIT
  reg  result_v; // @[Valid.scala 127:22]
  reg [31:0] result_b_z; // @[Reg.scala 16:16]
  reg  result_v_1; // @[Valid.scala 127:22]
  wire [31:0] result_nx = 32'sh26dd3b6a - 32'sh0; // @[Trigonometric.scala 67:54]
  wire [31:0] result_nz = $signed(result_b_z) - 32'sh3243f6a8; // @[Trigonometric.scala 71:51]
  wire  result_ns = $signed(result_nz) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_3 = 32'sh0 - $signed(result_nz); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_4 = $signed(result_nz) < 32'sh0 ? $signed(_result_improved_T_3) : $signed(result_nz); // @[Trigonometric.scala 79:15]
  wire  result_improved = $signed(_result_improved_T_4) < 32'sh40000000; // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_z; // @[Reg.scala 16:16]
  wire [31:0] _result_nx_T_11 = $signed(result_nextPipe_bits_x) - 32'sh136e9db5; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_15 = $signed(result_nextPipe_bits_x) + 32'sh136e9db5; // @[Trigonometric.scala 67:94]
  wire [30:0] _result_ny_T_8 = result_nextPipe_bits_x[31:1]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_264 = {{1{_result_ny_T_8[30]}},_result_ny_T_8}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_11 = 32'sh26dd3b6a + $signed(_GEN_264); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_15 = 32'sh26dd3b6a - $signed(_GEN_264); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_8 = $signed(result_nextPipe_bits_z) - 32'sh1dac6705; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_11 = $signed(result_nextPipe_bits_z) + 32'sh1dac6705; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_1 = result_nextPipe_bits_sigma ? $signed(_result_nz_T_8) : $signed(_result_nz_T_11); // @[Trigonometric.scala 71:21]
  wire  result_ns_1 = $signed(result_nz_1) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_1; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_1_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_1_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_1_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_1_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_13 = 32'sh0 - $signed(result_nz_1); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_14 = $signed(result_nz_1) < 32'sh0 ? $signed(_result_improved_T_13) : $signed(
    result_nz_1); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_18 = 32'sh0 - $signed(result_nextBestPipe_bits_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_19 = $signed(result_nextBestPipe_bits_z) < 32'sh0 ? $signed(_result_improved_T_18) :
    $signed(result_nextBestPipe_bits_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_1 = $signed(_result_improved_T_14) < $signed(_result_improved_T_19); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_1; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_1_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_1_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_1_z; // @[Reg.scala 16:16]
  wire [29:0] _result_nx_T_16 = result_nextPipe_bits_1_y[31:2]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_266 = {{2{_result_nx_T_16[29]}},_result_nx_T_16}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_19 = $signed(result_nextPipe_bits_1_x) - $signed(_GEN_266); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_23 = $signed(result_nextPipe_bits_1_x) + $signed(_GEN_266); // @[Trigonometric.scala 67:94]
  wire [29:0] _result_ny_T_16 = result_nextPipe_bits_1_x[31:2]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_268 = {{2{_result_ny_T_16[29]}},_result_ny_T_16}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_19 = $signed(result_nextPipe_bits_1_y) + $signed(_GEN_268); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_23 = $signed(result_nextPipe_bits_1_y) - $signed(_GEN_268); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_14 = $signed(result_nextPipe_bits_1_z) - 32'shfadbafc; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_17 = $signed(result_nextPipe_bits_1_z) + 32'shfadbafc; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_2 = result_nextPipe_bits_1_sigma ? $signed(_result_nz_T_14) : $signed(_result_nz_T_17); // @[Trigonometric.scala 71:21]
  wire  result_ns_2 = $signed(result_nz_2) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_2; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_2_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_2_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_2_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_2_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_23 = 32'sh0 - $signed(result_nz_2); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_24 = $signed(result_nz_2) < 32'sh0 ? $signed(_result_improved_T_23) : $signed(
    result_nz_2); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_28 = 32'sh0 - $signed(result_nextBestPipe_bits_1_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_29 = $signed(result_nextBestPipe_bits_1_z) < 32'sh0 ? $signed(_result_improved_T_28) :
    $signed(result_nextBestPipe_bits_1_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_2 = $signed(_result_improved_T_24) < $signed(_result_improved_T_29); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_2; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_2_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_2_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_2_z; // @[Reg.scala 16:16]
  wire [28:0] _result_nx_T_24 = result_nextPipe_bits_2_y[31:3]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_270 = {{3{_result_nx_T_24[28]}},_result_nx_T_24}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_27 = $signed(result_nextPipe_bits_2_x) - $signed(_GEN_270); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_31 = $signed(result_nextPipe_bits_2_x) + $signed(_GEN_270); // @[Trigonometric.scala 67:94]
  wire [28:0] _result_ny_T_24 = result_nextPipe_bits_2_x[31:3]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_272 = {{3{_result_ny_T_24[28]}},_result_ny_T_24}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_27 = $signed(result_nextPipe_bits_2_y) + $signed(_GEN_272); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_31 = $signed(result_nextPipe_bits_2_y) - $signed(_GEN_272); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_20 = $signed(result_nextPipe_bits_2_z) - 32'sh7f56ea6; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_23 = $signed(result_nextPipe_bits_2_z) + 32'sh7f56ea6; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_3 = result_nextPipe_bits_2_sigma ? $signed(_result_nz_T_20) : $signed(_result_nz_T_23); // @[Trigonometric.scala 71:21]
  wire  result_ns_3 = $signed(result_nz_3) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_3; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_3_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_3_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_3_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_3_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_33 = 32'sh0 - $signed(result_nz_3); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_34 = $signed(result_nz_3) < 32'sh0 ? $signed(_result_improved_T_33) : $signed(
    result_nz_3); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_38 = 32'sh0 - $signed(result_nextBestPipe_bits_2_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_39 = $signed(result_nextBestPipe_bits_2_z) < 32'sh0 ? $signed(_result_improved_T_38) :
    $signed(result_nextBestPipe_bits_2_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_3 = $signed(_result_improved_T_34) < $signed(_result_improved_T_39); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_3; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_3_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_3_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_3_z; // @[Reg.scala 16:16]
  wire [27:0] _result_nx_T_32 = result_nextPipe_bits_3_y[31:4]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_274 = {{4{_result_nx_T_32[27]}},_result_nx_T_32}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_35 = $signed(result_nextPipe_bits_3_x) - $signed(_GEN_274); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_39 = $signed(result_nextPipe_bits_3_x) + $signed(_GEN_274); // @[Trigonometric.scala 67:94]
  wire [27:0] _result_ny_T_32 = result_nextPipe_bits_3_x[31:4]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_276 = {{4{_result_ny_T_32[27]}},_result_ny_T_32}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_35 = $signed(result_nextPipe_bits_3_y) + $signed(_GEN_276); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_39 = $signed(result_nextPipe_bits_3_y) - $signed(_GEN_276); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_26 = $signed(result_nextPipe_bits_3_z) - 32'sh3feab76; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_29 = $signed(result_nextPipe_bits_3_z) + 32'sh3feab76; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_4 = result_nextPipe_bits_3_sigma ? $signed(_result_nz_T_26) : $signed(_result_nz_T_29); // @[Trigonometric.scala 71:21]
  wire  result_ns_4 = $signed(result_nz_4) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_4; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_4_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_4_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_4_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_4_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_43 = 32'sh0 - $signed(result_nz_4); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_44 = $signed(result_nz_4) < 32'sh0 ? $signed(_result_improved_T_43) : $signed(
    result_nz_4); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_48 = 32'sh0 - $signed(result_nextBestPipe_bits_3_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_49 = $signed(result_nextBestPipe_bits_3_z) < 32'sh0 ? $signed(_result_improved_T_48) :
    $signed(result_nextBestPipe_bits_3_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_4 = $signed(_result_improved_T_44) < $signed(_result_improved_T_49); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_4; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_4_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_4_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_4_z; // @[Reg.scala 16:16]
  wire [26:0] _result_nx_T_40 = result_nextPipe_bits_4_y[31:5]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_278 = {{5{_result_nx_T_40[26]}},_result_nx_T_40}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_43 = $signed(result_nextPipe_bits_4_x) - $signed(_GEN_278); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_47 = $signed(result_nextPipe_bits_4_x) + $signed(_GEN_278); // @[Trigonometric.scala 67:94]
  wire [26:0] _result_ny_T_40 = result_nextPipe_bits_4_x[31:5]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_280 = {{5{_result_ny_T_40[26]}},_result_ny_T_40}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_43 = $signed(result_nextPipe_bits_4_y) + $signed(_GEN_280); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_47 = $signed(result_nextPipe_bits_4_y) - $signed(_GEN_280); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_32 = $signed(result_nextPipe_bits_4_z) - 32'sh1ffd55b; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_35 = $signed(result_nextPipe_bits_4_z) + 32'sh1ffd55b; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_5 = result_nextPipe_bits_4_sigma ? $signed(_result_nz_T_32) : $signed(_result_nz_T_35); // @[Trigonometric.scala 71:21]
  wire  result_ns_5 = $signed(result_nz_5) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_5; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_5_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_5_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_5_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_5_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_53 = 32'sh0 - $signed(result_nz_5); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_54 = $signed(result_nz_5) < 32'sh0 ? $signed(_result_improved_T_53) : $signed(
    result_nz_5); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_58 = 32'sh0 - $signed(result_nextBestPipe_bits_4_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_59 = $signed(result_nextBestPipe_bits_4_z) < 32'sh0 ? $signed(_result_improved_T_58) :
    $signed(result_nextBestPipe_bits_4_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_5 = $signed(_result_improved_T_54) < $signed(_result_improved_T_59); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_5; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_5_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_5_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_5_z; // @[Reg.scala 16:16]
  wire [25:0] _result_nx_T_48 = result_nextPipe_bits_5_y[31:6]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_282 = {{6{_result_nx_T_48[25]}},_result_nx_T_48}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_51 = $signed(result_nextPipe_bits_5_x) - $signed(_GEN_282); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_55 = $signed(result_nextPipe_bits_5_x) + $signed(_GEN_282); // @[Trigonometric.scala 67:94]
  wire [25:0] _result_ny_T_48 = result_nextPipe_bits_5_x[31:6]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_284 = {{6{_result_ny_T_48[25]}},_result_ny_T_48}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_51 = $signed(result_nextPipe_bits_5_y) + $signed(_GEN_284); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_55 = $signed(result_nextPipe_bits_5_y) - $signed(_GEN_284); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_38 = $signed(result_nextPipe_bits_5_z) - 32'shfffaaa; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_41 = $signed(result_nextPipe_bits_5_z) + 32'shfffaaa; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_6 = result_nextPipe_bits_5_sigma ? $signed(_result_nz_T_38) : $signed(_result_nz_T_41); // @[Trigonometric.scala 71:21]
  wire  result_ns_6 = $signed(result_nz_6) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_6; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_6_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_6_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_6_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_6_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_63 = 32'sh0 - $signed(result_nz_6); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_64 = $signed(result_nz_6) < 32'sh0 ? $signed(_result_improved_T_63) : $signed(
    result_nz_6); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_68 = 32'sh0 - $signed(result_nextBestPipe_bits_5_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_69 = $signed(result_nextBestPipe_bits_5_z) < 32'sh0 ? $signed(_result_improved_T_68) :
    $signed(result_nextBestPipe_bits_5_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_6 = $signed(_result_improved_T_64) < $signed(_result_improved_T_69); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_6; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_6_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_6_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_6_z; // @[Reg.scala 16:16]
  wire [24:0] _result_nx_T_56 = result_nextPipe_bits_6_y[31:7]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_286 = {{7{_result_nx_T_56[24]}},_result_nx_T_56}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_59 = $signed(result_nextPipe_bits_6_x) - $signed(_GEN_286); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_63 = $signed(result_nextPipe_bits_6_x) + $signed(_GEN_286); // @[Trigonometric.scala 67:94]
  wire [24:0] _result_ny_T_56 = result_nextPipe_bits_6_x[31:7]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_288 = {{7{_result_ny_T_56[24]}},_result_ny_T_56}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_59 = $signed(result_nextPipe_bits_6_y) + $signed(_GEN_288); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_63 = $signed(result_nextPipe_bits_6_y) - $signed(_GEN_288); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_44 = $signed(result_nextPipe_bits_6_z) - 32'sh7fff55; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_47 = $signed(result_nextPipe_bits_6_z) + 32'sh7fff55; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_7 = result_nextPipe_bits_6_sigma ? $signed(_result_nz_T_44) : $signed(_result_nz_T_47); // @[Trigonometric.scala 71:21]
  wire  result_ns_7 = $signed(result_nz_7) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_7; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_7_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_7_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_7_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_7_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_73 = 32'sh0 - $signed(result_nz_7); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_74 = $signed(result_nz_7) < 32'sh0 ? $signed(_result_improved_T_73) : $signed(
    result_nz_7); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_78 = 32'sh0 - $signed(result_nextBestPipe_bits_6_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_79 = $signed(result_nextBestPipe_bits_6_z) < 32'sh0 ? $signed(_result_improved_T_78) :
    $signed(result_nextBestPipe_bits_6_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_7 = $signed(_result_improved_T_74) < $signed(_result_improved_T_79); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_7; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_7_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_7_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_7_z; // @[Reg.scala 16:16]
  wire [23:0] _result_nx_T_64 = result_nextPipe_bits_7_y[31:8]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_290 = {{8{_result_nx_T_64[23]}},_result_nx_T_64}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_67 = $signed(result_nextPipe_bits_7_x) - $signed(_GEN_290); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_71 = $signed(result_nextPipe_bits_7_x) + $signed(_GEN_290); // @[Trigonometric.scala 67:94]
  wire [23:0] _result_ny_T_64 = result_nextPipe_bits_7_x[31:8]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_292 = {{8{_result_ny_T_64[23]}},_result_ny_T_64}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_67 = $signed(result_nextPipe_bits_7_y) + $signed(_GEN_292); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_71 = $signed(result_nextPipe_bits_7_y) - $signed(_GEN_292); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_50 = $signed(result_nextPipe_bits_7_z) - 32'sh3fffea; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_53 = $signed(result_nextPipe_bits_7_z) + 32'sh3fffea; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_8 = result_nextPipe_bits_7_sigma ? $signed(_result_nz_T_50) : $signed(_result_nz_T_53); // @[Trigonometric.scala 71:21]
  wire  result_ns_8 = $signed(result_nz_8) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_8; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_8_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_8_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_8_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_8_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_83 = 32'sh0 - $signed(result_nz_8); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_84 = $signed(result_nz_8) < 32'sh0 ? $signed(_result_improved_T_83) : $signed(
    result_nz_8); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_88 = 32'sh0 - $signed(result_nextBestPipe_bits_7_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_89 = $signed(result_nextBestPipe_bits_7_z) < 32'sh0 ? $signed(_result_improved_T_88) :
    $signed(result_nextBestPipe_bits_7_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_8 = $signed(_result_improved_T_84) < $signed(_result_improved_T_89); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_8; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_8_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_8_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_8_z; // @[Reg.scala 16:16]
  wire [22:0] _result_nx_T_72 = result_nextPipe_bits_8_y[31:9]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_294 = {{9{_result_nx_T_72[22]}},_result_nx_T_72}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_75 = $signed(result_nextPipe_bits_8_x) - $signed(_GEN_294); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_79 = $signed(result_nextPipe_bits_8_x) + $signed(_GEN_294); // @[Trigonometric.scala 67:94]
  wire [22:0] _result_ny_T_72 = result_nextPipe_bits_8_x[31:9]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_296 = {{9{_result_ny_T_72[22]}},_result_ny_T_72}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_75 = $signed(result_nextPipe_bits_8_y) + $signed(_GEN_296); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_79 = $signed(result_nextPipe_bits_8_y) - $signed(_GEN_296); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_56 = $signed(result_nextPipe_bits_8_z) - 32'sh1ffffd; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_59 = $signed(result_nextPipe_bits_8_z) + 32'sh1ffffd; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_9 = result_nextPipe_bits_8_sigma ? $signed(_result_nz_T_56) : $signed(_result_nz_T_59); // @[Trigonometric.scala 71:21]
  wire  result_ns_9 = $signed(result_nz_9) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_9; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_9_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_9_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_9_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_9_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_93 = 32'sh0 - $signed(result_nz_9); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_94 = $signed(result_nz_9) < 32'sh0 ? $signed(_result_improved_T_93) : $signed(
    result_nz_9); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_98 = 32'sh0 - $signed(result_nextBestPipe_bits_8_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_99 = $signed(result_nextBestPipe_bits_8_z) < 32'sh0 ? $signed(_result_improved_T_98) :
    $signed(result_nextBestPipe_bits_8_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_9 = $signed(_result_improved_T_94) < $signed(_result_improved_T_99); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_9; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_9_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_9_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_9_z; // @[Reg.scala 16:16]
  wire [21:0] _result_nx_T_80 = result_nextPipe_bits_9_y[31:10]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_298 = {{10{_result_nx_T_80[21]}},_result_nx_T_80}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_83 = $signed(result_nextPipe_bits_9_x) - $signed(_GEN_298); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_87 = $signed(result_nextPipe_bits_9_x) + $signed(_GEN_298); // @[Trigonometric.scala 67:94]
  wire [21:0] _result_ny_T_80 = result_nextPipe_bits_9_x[31:10]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_300 = {{10{_result_ny_T_80[21]}},_result_ny_T_80}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_83 = $signed(result_nextPipe_bits_9_y) + $signed(_GEN_300); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_87 = $signed(result_nextPipe_bits_9_y) - $signed(_GEN_300); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_62 = $signed(result_nextPipe_bits_9_z) - 32'shfffff; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_65 = $signed(result_nextPipe_bits_9_z) + 32'shfffff; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_10 = result_nextPipe_bits_9_sigma ? $signed(_result_nz_T_62) : $signed(_result_nz_T_65); // @[Trigonometric.scala 71:21]
  wire  result_ns_10 = $signed(result_nz_10) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_10; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_10_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_10_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_10_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_10_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_103 = 32'sh0 - $signed(result_nz_10); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_104 = $signed(result_nz_10) < 32'sh0 ? $signed(_result_improved_T_103) : $signed(
    result_nz_10); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_108 = 32'sh0 - $signed(result_nextBestPipe_bits_9_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_109 = $signed(result_nextBestPipe_bits_9_z) < 32'sh0 ? $signed(_result_improved_T_108)
     : $signed(result_nextBestPipe_bits_9_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_10 = $signed(_result_improved_T_104) < $signed(_result_improved_T_109); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_10; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_10_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_10_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_10_z; // @[Reg.scala 16:16]
  wire [20:0] _result_nx_T_88 = result_nextPipe_bits_10_y[31:11]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_302 = {{11{_result_nx_T_88[20]}},_result_nx_T_88}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_91 = $signed(result_nextPipe_bits_10_x) - $signed(_GEN_302); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_95 = $signed(result_nextPipe_bits_10_x) + $signed(_GEN_302); // @[Trigonometric.scala 67:94]
  wire [20:0] _result_ny_T_88 = result_nextPipe_bits_10_x[31:11]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_304 = {{11{_result_ny_T_88[20]}},_result_ny_T_88}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_91 = $signed(result_nextPipe_bits_10_y) + $signed(_GEN_304); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_95 = $signed(result_nextPipe_bits_10_y) - $signed(_GEN_304); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_68 = $signed(result_nextPipe_bits_10_z) - 32'sh7ffff; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_71 = $signed(result_nextPipe_bits_10_z) + 32'sh7ffff; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_11 = result_nextPipe_bits_10_sigma ? $signed(_result_nz_T_68) : $signed(_result_nz_T_71); // @[Trigonometric.scala 71:21]
  wire  result_ns_11 = $signed(result_nz_11) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_11; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_11_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_11_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_11_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_11_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_113 = 32'sh0 - $signed(result_nz_11); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_114 = $signed(result_nz_11) < 32'sh0 ? $signed(_result_improved_T_113) : $signed(
    result_nz_11); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_118 = 32'sh0 - $signed(result_nextBestPipe_bits_10_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_119 = $signed(result_nextBestPipe_bits_10_z) < 32'sh0 ? $signed(_result_improved_T_118)
     : $signed(result_nextBestPipe_bits_10_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_11 = $signed(_result_improved_T_114) < $signed(_result_improved_T_119); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_11; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_11_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_11_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_11_z; // @[Reg.scala 16:16]
  wire [19:0] _result_nx_T_96 = result_nextPipe_bits_11_y[31:12]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_306 = {{12{_result_nx_T_96[19]}},_result_nx_T_96}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_99 = $signed(result_nextPipe_bits_11_x) - $signed(_GEN_306); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_103 = $signed(result_nextPipe_bits_11_x) + $signed(_GEN_306); // @[Trigonometric.scala 67:94]
  wire [19:0] _result_ny_T_96 = result_nextPipe_bits_11_x[31:12]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_308 = {{12{_result_ny_T_96[19]}},_result_ny_T_96}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_99 = $signed(result_nextPipe_bits_11_y) + $signed(_GEN_308); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_103 = $signed(result_nextPipe_bits_11_y) - $signed(_GEN_308); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_74 = $signed(result_nextPipe_bits_11_z) - 32'sh3ffff; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_77 = $signed(result_nextPipe_bits_11_z) + 32'sh3ffff; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_12 = result_nextPipe_bits_11_sigma ? $signed(_result_nz_T_74) : $signed(_result_nz_T_77); // @[Trigonometric.scala 71:21]
  wire  result_ns_12 = $signed(result_nz_12) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_12; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_12_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_12_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_12_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_12_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_123 = 32'sh0 - $signed(result_nz_12); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_124 = $signed(result_nz_12) < 32'sh0 ? $signed(_result_improved_T_123) : $signed(
    result_nz_12); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_128 = 32'sh0 - $signed(result_nextBestPipe_bits_11_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_129 = $signed(result_nextBestPipe_bits_11_z) < 32'sh0 ? $signed(_result_improved_T_128)
     : $signed(result_nextBestPipe_bits_11_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_12 = $signed(_result_improved_T_124) < $signed(_result_improved_T_129); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_12; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_12_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_12_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_12_z; // @[Reg.scala 16:16]
  wire [18:0] _result_nx_T_104 = result_nextPipe_bits_12_y[31:13]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_310 = {{13{_result_nx_T_104[18]}},_result_nx_T_104}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_107 = $signed(result_nextPipe_bits_12_x) - $signed(_GEN_310); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_111 = $signed(result_nextPipe_bits_12_x) + $signed(_GEN_310); // @[Trigonometric.scala 67:94]
  wire [18:0] _result_ny_T_104 = result_nextPipe_bits_12_x[31:13]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_312 = {{13{_result_ny_T_104[18]}},_result_ny_T_104}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_107 = $signed(result_nextPipe_bits_12_y) + $signed(_GEN_312); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_111 = $signed(result_nextPipe_bits_12_y) - $signed(_GEN_312); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_80 = $signed(result_nextPipe_bits_12_z) - 32'sh1ffff; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_83 = $signed(result_nextPipe_bits_12_z) + 32'sh1ffff; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_13 = result_nextPipe_bits_12_sigma ? $signed(_result_nz_T_80) : $signed(_result_nz_T_83); // @[Trigonometric.scala 71:21]
  wire  result_ns_13 = $signed(result_nz_13) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_13; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_13_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_13_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_13_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_13_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_133 = 32'sh0 - $signed(result_nz_13); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_134 = $signed(result_nz_13) < 32'sh0 ? $signed(_result_improved_T_133) : $signed(
    result_nz_13); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_138 = 32'sh0 - $signed(result_nextBestPipe_bits_12_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_139 = $signed(result_nextBestPipe_bits_12_z) < 32'sh0 ? $signed(_result_improved_T_138)
     : $signed(result_nextBestPipe_bits_12_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_13 = $signed(_result_improved_T_134) < $signed(_result_improved_T_139); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_13; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_13_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_13_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_13_z; // @[Reg.scala 16:16]
  wire [17:0] _result_nx_T_112 = result_nextPipe_bits_13_y[31:14]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_314 = {{14{_result_nx_T_112[17]}},_result_nx_T_112}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_115 = $signed(result_nextPipe_bits_13_x) - $signed(_GEN_314); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_119 = $signed(result_nextPipe_bits_13_x) + $signed(_GEN_314); // @[Trigonometric.scala 67:94]
  wire [17:0] _result_ny_T_112 = result_nextPipe_bits_13_x[31:14]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_316 = {{14{_result_ny_T_112[17]}},_result_ny_T_112}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_115 = $signed(result_nextPipe_bits_13_y) + $signed(_GEN_316); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_119 = $signed(result_nextPipe_bits_13_y) - $signed(_GEN_316); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_86 = $signed(result_nextPipe_bits_13_z) - 32'shffff; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_89 = $signed(result_nextPipe_bits_13_z) + 32'shffff; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_14 = result_nextPipe_bits_13_sigma ? $signed(_result_nz_T_86) : $signed(_result_nz_T_89); // @[Trigonometric.scala 71:21]
  wire  result_ns_14 = $signed(result_nz_14) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_14; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_14_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_14_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_14_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_14_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_143 = 32'sh0 - $signed(result_nz_14); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_144 = $signed(result_nz_14) < 32'sh0 ? $signed(_result_improved_T_143) : $signed(
    result_nz_14); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_148 = 32'sh0 - $signed(result_nextBestPipe_bits_13_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_149 = $signed(result_nextBestPipe_bits_13_z) < 32'sh0 ? $signed(_result_improved_T_148)
     : $signed(result_nextBestPipe_bits_13_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_14 = $signed(_result_improved_T_144) < $signed(_result_improved_T_149); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_14; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_14_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_14_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_14_z; // @[Reg.scala 16:16]
  wire [16:0] _result_nx_T_120 = result_nextPipe_bits_14_y[31:15]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_318 = {{15{_result_nx_T_120[16]}},_result_nx_T_120}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_123 = $signed(result_nextPipe_bits_14_x) - $signed(_GEN_318); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_127 = $signed(result_nextPipe_bits_14_x) + $signed(_GEN_318); // @[Trigonometric.scala 67:94]
  wire [16:0] _result_ny_T_120 = result_nextPipe_bits_14_x[31:15]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_320 = {{15{_result_ny_T_120[16]}},_result_ny_T_120}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_123 = $signed(result_nextPipe_bits_14_y) + $signed(_GEN_320); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_127 = $signed(result_nextPipe_bits_14_y) - $signed(_GEN_320); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_92 = $signed(result_nextPipe_bits_14_z) - 32'sh7fff; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_95 = $signed(result_nextPipe_bits_14_z) + 32'sh7fff; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_15 = result_nextPipe_bits_14_sigma ? $signed(_result_nz_T_92) : $signed(_result_nz_T_95); // @[Trigonometric.scala 71:21]
  wire  result_ns_15 = $signed(result_nz_15) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_15; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_15_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_15_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_15_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_15_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_153 = 32'sh0 - $signed(result_nz_15); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_154 = $signed(result_nz_15) < 32'sh0 ? $signed(_result_improved_T_153) : $signed(
    result_nz_15); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_158 = 32'sh0 - $signed(result_nextBestPipe_bits_14_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_159 = $signed(result_nextBestPipe_bits_14_z) < 32'sh0 ? $signed(_result_improved_T_158)
     : $signed(result_nextBestPipe_bits_14_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_15 = $signed(_result_improved_T_154) < $signed(_result_improved_T_159); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_15; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_15_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_15_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_15_z; // @[Reg.scala 16:16]
  wire [15:0] _result_nx_T_128 = result_nextPipe_bits_15_y[31:16]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_322 = {{16{_result_nx_T_128[15]}},_result_nx_T_128}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_131 = $signed(result_nextPipe_bits_15_x) - $signed(_GEN_322); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_135 = $signed(result_nextPipe_bits_15_x) + $signed(_GEN_322); // @[Trigonometric.scala 67:94]
  wire [15:0] _result_ny_T_128 = result_nextPipe_bits_15_x[31:16]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_324 = {{16{_result_ny_T_128[15]}},_result_ny_T_128}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_131 = $signed(result_nextPipe_bits_15_y) + $signed(_GEN_324); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_135 = $signed(result_nextPipe_bits_15_y) - $signed(_GEN_324); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_98 = $signed(result_nextPipe_bits_15_z) - 32'sh3fff; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_101 = $signed(result_nextPipe_bits_15_z) + 32'sh3fff; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_16 = result_nextPipe_bits_15_sigma ? $signed(_result_nz_T_98) : $signed(_result_nz_T_101); // @[Trigonometric.scala 71:21]
  wire  result_ns_16 = $signed(result_nz_16) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_16; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_16_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_16_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_16_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_16_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_163 = 32'sh0 - $signed(result_nz_16); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_164 = $signed(result_nz_16) < 32'sh0 ? $signed(_result_improved_T_163) : $signed(
    result_nz_16); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_168 = 32'sh0 - $signed(result_nextBestPipe_bits_15_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_169 = $signed(result_nextBestPipe_bits_15_z) < 32'sh0 ? $signed(_result_improved_T_168)
     : $signed(result_nextBestPipe_bits_15_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_16 = $signed(_result_improved_T_164) < $signed(_result_improved_T_169); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_16; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_16_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_16_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_16_z; // @[Reg.scala 16:16]
  wire [14:0] _result_nx_T_136 = result_nextPipe_bits_16_y[31:17]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_326 = {{17{_result_nx_T_136[14]}},_result_nx_T_136}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_139 = $signed(result_nextPipe_bits_16_x) - $signed(_GEN_326); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_143 = $signed(result_nextPipe_bits_16_x) + $signed(_GEN_326); // @[Trigonometric.scala 67:94]
  wire [14:0] _result_ny_T_136 = result_nextPipe_bits_16_x[31:17]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_328 = {{17{_result_ny_T_136[14]}},_result_ny_T_136}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_139 = $signed(result_nextPipe_bits_16_y) + $signed(_GEN_328); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_143 = $signed(result_nextPipe_bits_16_y) - $signed(_GEN_328); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_104 = $signed(result_nextPipe_bits_16_z) - 32'sh1fff; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_107 = $signed(result_nextPipe_bits_16_z) + 32'sh1fff; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_17 = result_nextPipe_bits_16_sigma ? $signed(_result_nz_T_104) : $signed(_result_nz_T_107); // @[Trigonometric.scala 71:21]
  wire  result_ns_17 = $signed(result_nz_17) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_17; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_17_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_17_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_17_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_17_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_173 = 32'sh0 - $signed(result_nz_17); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_174 = $signed(result_nz_17) < 32'sh0 ? $signed(_result_improved_T_173) : $signed(
    result_nz_17); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_178 = 32'sh0 - $signed(result_nextBestPipe_bits_16_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_179 = $signed(result_nextBestPipe_bits_16_z) < 32'sh0 ? $signed(_result_improved_T_178)
     : $signed(result_nextBestPipe_bits_16_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_17 = $signed(_result_improved_T_174) < $signed(_result_improved_T_179); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_17; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_17_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_17_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_17_z; // @[Reg.scala 16:16]
  wire [13:0] _result_nx_T_144 = result_nextPipe_bits_17_y[31:18]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_330 = {{18{_result_nx_T_144[13]}},_result_nx_T_144}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_147 = $signed(result_nextPipe_bits_17_x) - $signed(_GEN_330); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_151 = $signed(result_nextPipe_bits_17_x) + $signed(_GEN_330); // @[Trigonometric.scala 67:94]
  wire [13:0] _result_ny_T_144 = result_nextPipe_bits_17_x[31:18]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_332 = {{18{_result_ny_T_144[13]}},_result_ny_T_144}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_147 = $signed(result_nextPipe_bits_17_y) + $signed(_GEN_332); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_151 = $signed(result_nextPipe_bits_17_y) - $signed(_GEN_332); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_110 = $signed(result_nextPipe_bits_17_z) - 32'shfff; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_113 = $signed(result_nextPipe_bits_17_z) + 32'shfff; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_18 = result_nextPipe_bits_17_sigma ? $signed(_result_nz_T_110) : $signed(_result_nz_T_113); // @[Trigonometric.scala 71:21]
  wire  result_ns_18 = $signed(result_nz_18) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_18; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_18_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_18_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_18_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_18_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_183 = 32'sh0 - $signed(result_nz_18); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_184 = $signed(result_nz_18) < 32'sh0 ? $signed(_result_improved_T_183) : $signed(
    result_nz_18); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_188 = 32'sh0 - $signed(result_nextBestPipe_bits_17_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_189 = $signed(result_nextBestPipe_bits_17_z) < 32'sh0 ? $signed(_result_improved_T_188)
     : $signed(result_nextBestPipe_bits_17_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_18 = $signed(_result_improved_T_184) < $signed(_result_improved_T_189); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_18; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_18_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_18_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_18_z; // @[Reg.scala 16:16]
  wire [12:0] _result_nx_T_152 = result_nextPipe_bits_18_y[31:19]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_334 = {{19{_result_nx_T_152[12]}},_result_nx_T_152}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_155 = $signed(result_nextPipe_bits_18_x) - $signed(_GEN_334); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_159 = $signed(result_nextPipe_bits_18_x) + $signed(_GEN_334); // @[Trigonometric.scala 67:94]
  wire [12:0] _result_ny_T_152 = result_nextPipe_bits_18_x[31:19]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_336 = {{19{_result_ny_T_152[12]}},_result_ny_T_152}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_155 = $signed(result_nextPipe_bits_18_y) + $signed(_GEN_336); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_159 = $signed(result_nextPipe_bits_18_y) - $signed(_GEN_336); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_116 = $signed(result_nextPipe_bits_18_z) - 32'sh7ff; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_119 = $signed(result_nextPipe_bits_18_z) + 32'sh7ff; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_19 = result_nextPipe_bits_18_sigma ? $signed(_result_nz_T_116) : $signed(_result_nz_T_119); // @[Trigonometric.scala 71:21]
  wire  result_ns_19 = $signed(result_nz_19) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_19; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_19_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_19_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_19_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_19_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_193 = 32'sh0 - $signed(result_nz_19); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_194 = $signed(result_nz_19) < 32'sh0 ? $signed(_result_improved_T_193) : $signed(
    result_nz_19); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_198 = 32'sh0 - $signed(result_nextBestPipe_bits_18_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_199 = $signed(result_nextBestPipe_bits_18_z) < 32'sh0 ? $signed(_result_improved_T_198)
     : $signed(result_nextBestPipe_bits_18_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_19 = $signed(_result_improved_T_194) < $signed(_result_improved_T_199); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_19; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_19_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_19_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_19_z; // @[Reg.scala 16:16]
  wire [11:0] _result_nx_T_160 = result_nextPipe_bits_19_y[31:20]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_338 = {{20{_result_nx_T_160[11]}},_result_nx_T_160}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_163 = $signed(result_nextPipe_bits_19_x) - $signed(_GEN_338); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_167 = $signed(result_nextPipe_bits_19_x) + $signed(_GEN_338); // @[Trigonometric.scala 67:94]
  wire [11:0] _result_ny_T_160 = result_nextPipe_bits_19_x[31:20]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_340 = {{20{_result_ny_T_160[11]}},_result_ny_T_160}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_163 = $signed(result_nextPipe_bits_19_y) + $signed(_GEN_340); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_167 = $signed(result_nextPipe_bits_19_y) - $signed(_GEN_340); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_122 = $signed(result_nextPipe_bits_19_z) - 32'sh3ff; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_125 = $signed(result_nextPipe_bits_19_z) + 32'sh3ff; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_20 = result_nextPipe_bits_19_sigma ? $signed(_result_nz_T_122) : $signed(_result_nz_T_125); // @[Trigonometric.scala 71:21]
  wire  result_ns_20 = $signed(result_nz_20) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_20; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_20_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_20_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_20_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_20_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_203 = 32'sh0 - $signed(result_nz_20); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_204 = $signed(result_nz_20) < 32'sh0 ? $signed(_result_improved_T_203) : $signed(
    result_nz_20); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_208 = 32'sh0 - $signed(result_nextBestPipe_bits_19_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_209 = $signed(result_nextBestPipe_bits_19_z) < 32'sh0 ? $signed(_result_improved_T_208)
     : $signed(result_nextBestPipe_bits_19_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_20 = $signed(_result_improved_T_204) < $signed(_result_improved_T_209); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_20; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_20_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_20_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_20_z; // @[Reg.scala 16:16]
  wire [10:0] _result_nx_T_168 = result_nextPipe_bits_20_y[31:21]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_342 = {{21{_result_nx_T_168[10]}},_result_nx_T_168}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_171 = $signed(result_nextPipe_bits_20_x) - $signed(_GEN_342); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_175 = $signed(result_nextPipe_bits_20_x) + $signed(_GEN_342); // @[Trigonometric.scala 67:94]
  wire [10:0] _result_ny_T_168 = result_nextPipe_bits_20_x[31:21]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_344 = {{21{_result_ny_T_168[10]}},_result_ny_T_168}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_171 = $signed(result_nextPipe_bits_20_y) + $signed(_GEN_344); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_175 = $signed(result_nextPipe_bits_20_y) - $signed(_GEN_344); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_128 = $signed(result_nextPipe_bits_20_z) - 32'sh1ff; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_131 = $signed(result_nextPipe_bits_20_z) + 32'sh1ff; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_21 = result_nextPipe_bits_20_sigma ? $signed(_result_nz_T_128) : $signed(_result_nz_T_131); // @[Trigonometric.scala 71:21]
  wire  result_ns_21 = $signed(result_nz_21) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_21; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_21_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_21_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_21_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_21_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_213 = 32'sh0 - $signed(result_nz_21); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_214 = $signed(result_nz_21) < 32'sh0 ? $signed(_result_improved_T_213) : $signed(
    result_nz_21); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_218 = 32'sh0 - $signed(result_nextBestPipe_bits_20_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_219 = $signed(result_nextBestPipe_bits_20_z) < 32'sh0 ? $signed(_result_improved_T_218)
     : $signed(result_nextBestPipe_bits_20_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_21 = $signed(_result_improved_T_214) < $signed(_result_improved_T_219); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_21; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_21_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_21_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_21_z; // @[Reg.scala 16:16]
  wire [9:0] _result_nx_T_176 = result_nextPipe_bits_21_y[31:22]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_346 = {{22{_result_nx_T_176[9]}},_result_nx_T_176}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_179 = $signed(result_nextPipe_bits_21_x) - $signed(_GEN_346); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_183 = $signed(result_nextPipe_bits_21_x) + $signed(_GEN_346); // @[Trigonometric.scala 67:94]
  wire [9:0] _result_ny_T_176 = result_nextPipe_bits_21_x[31:22]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_348 = {{22{_result_ny_T_176[9]}},_result_ny_T_176}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_179 = $signed(result_nextPipe_bits_21_y) + $signed(_GEN_348); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_183 = $signed(result_nextPipe_bits_21_y) - $signed(_GEN_348); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_134 = $signed(result_nextPipe_bits_21_z) - 32'shff; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_137 = $signed(result_nextPipe_bits_21_z) + 32'shff; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_22 = result_nextPipe_bits_21_sigma ? $signed(_result_nz_T_134) : $signed(_result_nz_T_137); // @[Trigonometric.scala 71:21]
  wire  result_ns_22 = $signed(result_nz_22) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_22; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_22_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_22_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_22_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_22_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_223 = 32'sh0 - $signed(result_nz_22); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_224 = $signed(result_nz_22) < 32'sh0 ? $signed(_result_improved_T_223) : $signed(
    result_nz_22); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_228 = 32'sh0 - $signed(result_nextBestPipe_bits_21_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_229 = $signed(result_nextBestPipe_bits_21_z) < 32'sh0 ? $signed(_result_improved_T_228)
     : $signed(result_nextBestPipe_bits_21_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_22 = $signed(_result_improved_T_224) < $signed(_result_improved_T_229); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_22; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_22_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_22_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_22_z; // @[Reg.scala 16:16]
  wire [8:0] _result_nx_T_184 = result_nextPipe_bits_22_y[31:23]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_350 = {{23{_result_nx_T_184[8]}},_result_nx_T_184}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_187 = $signed(result_nextPipe_bits_22_x) - $signed(_GEN_350); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_191 = $signed(result_nextPipe_bits_22_x) + $signed(_GEN_350); // @[Trigonometric.scala 67:94]
  wire [8:0] _result_ny_T_184 = result_nextPipe_bits_22_x[31:23]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_352 = {{23{_result_ny_T_184[8]}},_result_ny_T_184}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_187 = $signed(result_nextPipe_bits_22_y) + $signed(_GEN_352); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_191 = $signed(result_nextPipe_bits_22_y) - $signed(_GEN_352); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_140 = $signed(result_nextPipe_bits_22_z) - 32'sh7f; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_143 = $signed(result_nextPipe_bits_22_z) + 32'sh7f; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_23 = result_nextPipe_bits_22_sigma ? $signed(_result_nz_T_140) : $signed(_result_nz_T_143); // @[Trigonometric.scala 71:21]
  wire  result_ns_23 = $signed(result_nz_23) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_23; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_23_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_23_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_23_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_23_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_233 = 32'sh0 - $signed(result_nz_23); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_234 = $signed(result_nz_23) < 32'sh0 ? $signed(_result_improved_T_233) : $signed(
    result_nz_23); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_238 = 32'sh0 - $signed(result_nextBestPipe_bits_22_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_239 = $signed(result_nextBestPipe_bits_22_z) < 32'sh0 ? $signed(_result_improved_T_238)
     : $signed(result_nextBestPipe_bits_22_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_23 = $signed(_result_improved_T_234) < $signed(_result_improved_T_239); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_23; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_23_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_23_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_23_z; // @[Reg.scala 16:16]
  wire [7:0] _result_nx_T_192 = result_nextPipe_bits_23_y[31:24]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_354 = {{24{_result_nx_T_192[7]}},_result_nx_T_192}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_195 = $signed(result_nextPipe_bits_23_x) - $signed(_GEN_354); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_199 = $signed(result_nextPipe_bits_23_x) + $signed(_GEN_354); // @[Trigonometric.scala 67:94]
  wire [7:0] _result_ny_T_192 = result_nextPipe_bits_23_x[31:24]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_356 = {{24{_result_ny_T_192[7]}},_result_ny_T_192}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_195 = $signed(result_nextPipe_bits_23_y) + $signed(_GEN_356); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_199 = $signed(result_nextPipe_bits_23_y) - $signed(_GEN_356); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_146 = $signed(result_nextPipe_bits_23_z) - 32'sh3f; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_149 = $signed(result_nextPipe_bits_23_z) + 32'sh3f; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_24 = result_nextPipe_bits_23_sigma ? $signed(_result_nz_T_146) : $signed(_result_nz_T_149); // @[Trigonometric.scala 71:21]
  wire  result_ns_24 = $signed(result_nz_24) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_24; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_24_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_24_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_24_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_24_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_243 = 32'sh0 - $signed(result_nz_24); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_244 = $signed(result_nz_24) < 32'sh0 ? $signed(_result_improved_T_243) : $signed(
    result_nz_24); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_248 = 32'sh0 - $signed(result_nextBestPipe_bits_23_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_249 = $signed(result_nextBestPipe_bits_23_z) < 32'sh0 ? $signed(_result_improved_T_248)
     : $signed(result_nextBestPipe_bits_23_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_24 = $signed(_result_improved_T_244) < $signed(_result_improved_T_249); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_24; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_24_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_24_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_24_z; // @[Reg.scala 16:16]
  wire [6:0] _result_nx_T_200 = result_nextPipe_bits_24_y[31:25]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_358 = {{25{_result_nx_T_200[6]}},_result_nx_T_200}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_203 = $signed(result_nextPipe_bits_24_x) - $signed(_GEN_358); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_207 = $signed(result_nextPipe_bits_24_x) + $signed(_GEN_358); // @[Trigonometric.scala 67:94]
  wire [6:0] _result_ny_T_200 = result_nextPipe_bits_24_x[31:25]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_360 = {{25{_result_ny_T_200[6]}},_result_ny_T_200}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_203 = $signed(result_nextPipe_bits_24_y) + $signed(_GEN_360); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_207 = $signed(result_nextPipe_bits_24_y) - $signed(_GEN_360); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_152 = $signed(result_nextPipe_bits_24_z) - 32'sh1f; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_155 = $signed(result_nextPipe_bits_24_z) + 32'sh1f; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_25 = result_nextPipe_bits_24_sigma ? $signed(_result_nz_T_152) : $signed(_result_nz_T_155); // @[Trigonometric.scala 71:21]
  wire  result_ns_25 = $signed(result_nz_25) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_25; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_25_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_25_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_25_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_25_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_253 = 32'sh0 - $signed(result_nz_25); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_254 = $signed(result_nz_25) < 32'sh0 ? $signed(_result_improved_T_253) : $signed(
    result_nz_25); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_258 = 32'sh0 - $signed(result_nextBestPipe_bits_24_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_259 = $signed(result_nextBestPipe_bits_24_z) < 32'sh0 ? $signed(_result_improved_T_258)
     : $signed(result_nextBestPipe_bits_24_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_25 = $signed(_result_improved_T_254) < $signed(_result_improved_T_259); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_25; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_25_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_25_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_25_z; // @[Reg.scala 16:16]
  wire [5:0] _result_nx_T_208 = result_nextPipe_bits_25_y[31:26]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_362 = {{26{_result_nx_T_208[5]}},_result_nx_T_208}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_211 = $signed(result_nextPipe_bits_25_x) - $signed(_GEN_362); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_215 = $signed(result_nextPipe_bits_25_x) + $signed(_GEN_362); // @[Trigonometric.scala 67:94]
  wire [5:0] _result_ny_T_208 = result_nextPipe_bits_25_x[31:26]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_364 = {{26{_result_ny_T_208[5]}},_result_ny_T_208}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_211 = $signed(result_nextPipe_bits_25_y) + $signed(_GEN_364); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_215 = $signed(result_nextPipe_bits_25_y) - $signed(_GEN_364); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_158 = $signed(result_nextPipe_bits_25_z) - 32'shf; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_161 = $signed(result_nextPipe_bits_25_z) + 32'shf; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_26 = result_nextPipe_bits_25_sigma ? $signed(_result_nz_T_158) : $signed(_result_nz_T_161); // @[Trigonometric.scala 71:21]
  wire  result_ns_26 = $signed(result_nz_26) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_26; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_26_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_26_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_26_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_26_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_263 = 32'sh0 - $signed(result_nz_26); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_264 = $signed(result_nz_26) < 32'sh0 ? $signed(_result_improved_T_263) : $signed(
    result_nz_26); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_268 = 32'sh0 - $signed(result_nextBestPipe_bits_25_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_269 = $signed(result_nextBestPipe_bits_25_z) < 32'sh0 ? $signed(_result_improved_T_268)
     : $signed(result_nextBestPipe_bits_25_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_26 = $signed(_result_improved_T_264) < $signed(_result_improved_T_269); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_26; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_26_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_26_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_26_z; // @[Reg.scala 16:16]
  wire [4:0] _result_nx_T_216 = result_nextPipe_bits_26_y[31:27]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_366 = {{27{_result_nx_T_216[4]}},_result_nx_T_216}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_219 = $signed(result_nextPipe_bits_26_x) - $signed(_GEN_366); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_223 = $signed(result_nextPipe_bits_26_x) + $signed(_GEN_366); // @[Trigonometric.scala 67:94]
  wire [4:0] _result_ny_T_216 = result_nextPipe_bits_26_x[31:27]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_368 = {{27{_result_ny_T_216[4]}},_result_ny_T_216}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_219 = $signed(result_nextPipe_bits_26_y) + $signed(_GEN_368); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_223 = $signed(result_nextPipe_bits_26_y) - $signed(_GEN_368); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_164 = $signed(result_nextPipe_bits_26_z) - 32'sh8; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_167 = $signed(result_nextPipe_bits_26_z) + 32'sh8; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_27 = result_nextPipe_bits_26_sigma ? $signed(_result_nz_T_164) : $signed(_result_nz_T_167); // @[Trigonometric.scala 71:21]
  wire  result_ns_27 = $signed(result_nz_27) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_27; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_27_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_27_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_27_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_27_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_273 = 32'sh0 - $signed(result_nz_27); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_274 = $signed(result_nz_27) < 32'sh0 ? $signed(_result_improved_T_273) : $signed(
    result_nz_27); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_278 = 32'sh0 - $signed(result_nextBestPipe_bits_26_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_279 = $signed(result_nextBestPipe_bits_26_z) < 32'sh0 ? $signed(_result_improved_T_278)
     : $signed(result_nextBestPipe_bits_26_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_27 = $signed(_result_improved_T_274) < $signed(_result_improved_T_279); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_27; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_27_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_27_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_27_z; // @[Reg.scala 16:16]
  wire [3:0] _result_nx_T_224 = result_nextPipe_bits_27_y[31:28]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_370 = {{28{_result_nx_T_224[3]}},_result_nx_T_224}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_227 = $signed(result_nextPipe_bits_27_x) - $signed(_GEN_370); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_231 = $signed(result_nextPipe_bits_27_x) + $signed(_GEN_370); // @[Trigonometric.scala 67:94]
  wire [3:0] _result_ny_T_224 = result_nextPipe_bits_27_x[31:28]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_372 = {{28{_result_ny_T_224[3]}},_result_ny_T_224}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_227 = $signed(result_nextPipe_bits_27_y) + $signed(_GEN_372); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_231 = $signed(result_nextPipe_bits_27_y) - $signed(_GEN_372); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_170 = $signed(result_nextPipe_bits_27_z) - 32'sh4; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_173 = $signed(result_nextPipe_bits_27_z) + 32'sh4; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_28 = result_nextPipe_bits_27_sigma ? $signed(_result_nz_T_170) : $signed(_result_nz_T_173); // @[Trigonometric.scala 71:21]
  wire  result_ns_28 = $signed(result_nz_28) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_28; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_28_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_28_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_28_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_28_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_283 = 32'sh0 - $signed(result_nz_28); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_284 = $signed(result_nz_28) < 32'sh0 ? $signed(_result_improved_T_283) : $signed(
    result_nz_28); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_288 = 32'sh0 - $signed(result_nextBestPipe_bits_27_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_289 = $signed(result_nextBestPipe_bits_27_z) < 32'sh0 ? $signed(_result_improved_T_288)
     : $signed(result_nextBestPipe_bits_27_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_28 = $signed(_result_improved_T_284) < $signed(_result_improved_T_289); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_28; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_28_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_28_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_28_z; // @[Reg.scala 16:16]
  wire [2:0] _result_nx_T_232 = result_nextPipe_bits_28_y[31:29]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_374 = {{29{_result_nx_T_232[2]}},_result_nx_T_232}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_235 = $signed(result_nextPipe_bits_28_x) - $signed(_GEN_374); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_239 = $signed(result_nextPipe_bits_28_x) + $signed(_GEN_374); // @[Trigonometric.scala 67:94]
  wire [2:0] _result_ny_T_232 = result_nextPipe_bits_28_x[31:29]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_376 = {{29{_result_ny_T_232[2]}},_result_ny_T_232}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_235 = $signed(result_nextPipe_bits_28_y) + $signed(_GEN_376); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_239 = $signed(result_nextPipe_bits_28_y) - $signed(_GEN_376); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_176 = $signed(result_nextPipe_bits_28_z) - 32'sh2; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_179 = $signed(result_nextPipe_bits_28_z) + 32'sh2; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_29 = result_nextPipe_bits_28_sigma ? $signed(_result_nz_T_176) : $signed(_result_nz_T_179); // @[Trigonometric.scala 71:21]
  wire  result_ns_29 = $signed(result_nz_29) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg  result_nextPipe_valid_29; // @[Valid.scala 127:22]
  reg [31:0] result_nextPipe_bits_29_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_29_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_29_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_29_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_293 = 32'sh0 - $signed(result_nz_29); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_294 = $signed(result_nz_29) < 32'sh0 ? $signed(_result_improved_T_293) : $signed(
    result_nz_29); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_298 = 32'sh0 - $signed(result_nextBestPipe_bits_28_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_299 = $signed(result_nextBestPipe_bits_28_z) < 32'sh0 ? $signed(_result_improved_T_298)
     : $signed(result_nextBestPipe_bits_28_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_29 = $signed(_result_improved_T_294) < $signed(_result_improved_T_299); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_29; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_29_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_29_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_29_z; // @[Reg.scala 16:16]
  wire [1:0] _result_nx_T_240 = result_nextPipe_bits_29_y[31:30]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_378 = {{30{_result_nx_T_240[1]}},_result_nx_T_240}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_243 = $signed(result_nextPipe_bits_29_x) - $signed(_GEN_378); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_247 = $signed(result_nextPipe_bits_29_x) + $signed(_GEN_378); // @[Trigonometric.scala 67:94]
  wire [1:0] _result_ny_T_240 = result_nextPipe_bits_29_x[31:30]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_380 = {{30{_result_ny_T_240[1]}},_result_ny_T_240}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_243 = $signed(result_nextPipe_bits_29_y) + $signed(_GEN_380); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_247 = $signed(result_nextPipe_bits_29_y) - $signed(_GEN_380); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_182 = $signed(result_nextPipe_bits_29_z) - 32'sh1; // @[Trigonometric.scala 71:51]
  wire [31:0] _result_nz_T_185 = $signed(result_nextPipe_bits_29_z) + 32'sh1; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_30 = result_nextPipe_bits_29_sigma ? $signed(_result_nz_T_182) : $signed(_result_nz_T_185); // @[Trigonometric.scala 71:21]
  wire  result_ns_30 = $signed(result_nz_30) > 32'sh0; // @[Trigonometric.scala 72:21]
  reg [31:0] result_nextPipe_bits_30_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_30_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextPipe_bits_30_z; // @[Reg.scala 16:16]
  reg  result_nextPipe_bits_30_sigma; // @[Reg.scala 16:16]
  wire [31:0] _result_improved_T_303 = 32'sh0 - $signed(result_nz_30); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_304 = $signed(result_nz_30) < 32'sh0 ? $signed(_result_improved_T_303) : $signed(
    result_nz_30); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_308 = 32'sh0 - $signed(result_nextBestPipe_bits_29_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_309 = $signed(result_nextBestPipe_bits_29_z) < 32'sh0 ? $signed(_result_improved_T_308)
     : $signed(result_nextBestPipe_bits_29_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_30 = $signed(_result_improved_T_304) < $signed(_result_improved_T_309); // @[Trigonometric.scala 79:19]
  reg  result_nextBestPipe_valid_30; // @[Valid.scala 127:22]
  reg [31:0] result_nextBestPipe_bits_30_x; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_30_y; // @[Reg.scala 16:16]
  reg [31:0] result_nextBestPipe_bits_30_z; // @[Reg.scala 16:16]
  wire  _result_nx_T_248 = result_nextPipe_bits_30_y[31]; // @[Trigonometric.scala 67:69]
  wire [31:0] _GEN_382 = {32{_result_nx_T_248}}; // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_251 = $signed(result_nextPipe_bits_30_x) - $signed(_GEN_382); // @[Trigonometric.scala 67:54]
  wire [31:0] _result_nx_T_255 = $signed(result_nextPipe_bits_30_x) + $signed(_GEN_382); // @[Trigonometric.scala 67:94]
  wire  _result_ny_T_248 = result_nextPipe_bits_30_x[31]; // @[Trigonometric.scala 68:69]
  wire [31:0] _GEN_384 = {32{_result_ny_T_248}}; // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_251 = $signed(result_nextPipe_bits_30_y) + $signed(_GEN_384); // @[Trigonometric.scala 68:54]
  wire [31:0] _result_ny_T_255 = $signed(result_nextPipe_bits_30_y) - $signed(_GEN_384); // @[Trigonometric.scala 68:94]
  wire [31:0] _result_nz_T_188 = $signed(result_nextPipe_bits_30_z) - 32'sh0; // @[Trigonometric.scala 71:51]
  wire [32:0] _result_nz_T_189 = {{1{result_nextPipe_bits_30_z[31]}},result_nextPipe_bits_30_z}; // @[Trigonometric.scala 71:72]
  wire [31:0] _result_nz_T_191 = _result_nz_T_189[31:0]; // @[Trigonometric.scala 71:72]
  wire [31:0] result_nz_31 = result_nextPipe_bits_30_sigma ? $signed(_result_nz_T_188) : $signed(_result_nz_T_191); // @[Trigonometric.scala 71:21]
  wire [31:0] _result_improved_T_313 = 32'sh0 - $signed(result_nz_31); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_314 = $signed(result_nz_31) < 32'sh0 ? $signed(_result_improved_T_313) : $signed(
    result_nz_31); // @[Trigonometric.scala 79:15]
  wire [31:0] _result_improved_T_318 = 32'sh0 - $signed(result_nextBestPipe_bits_30_z); // @[Trigonometric.scala 79:37]
  wire [31:0] _result_improved_T_319 = $signed(result_nextBestPipe_bits_30_z) < 32'sh0 ? $signed(_result_improved_T_318)
     : $signed(result_nextBestPipe_bits_30_z); // @[Trigonometric.scala 79:37]
  wire  result_improved_31 = $signed(_result_improved_T_314) < $signed(_result_improved_T_319); // @[Trigonometric.scala 79:19]
  reg  resultPipe_valid; // @[Valid.scala 127:22]
  reg [31:0] resultPipe_bits_x; // @[Reg.scala 16:16]
  reg [31:0] resultPipe_bits_y; // @[Reg.scala 16:16]
  assign io_result_valid = resultPipe_valid; // @[Valid.scala 122:21 123:17]
  assign io_result_bits_sine = resultPipe_bits_y; // @[Valid.scala 122:21 124:16]
  assign io_result_bits_cosine = resultPipe_bits_x; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      result_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_v <= io_theta_valid; // @[Valid.scala 127:22]
    end
    if (io_theta_valid) begin // @[Reg.scala 17:18]
      result_b_z <= io_theta_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_v_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_v_1 <= io_theta_valid; // @[Valid.scala 127:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid <= result_v; // @[Valid.scala 127:22]
    end
    if (result_v) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_x <= result_nx; // @[Reg.scala 17:22]
    end
    if (result_v) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_z <= result_nz; // @[Reg.scala 17:22]
    end
    if (result_v) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_sigma <= result_ns; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid <= result_v_1; // @[Valid.scala 127:22]
    end
    if (result_v_1) begin // @[Reg.scala 17:18]
      if (result_improved) begin // @[Trigonometric.scala 84:14]
        result_nextBestPipe_bits_x <= result_nx;
      end else begin
        result_nextBestPipe_bits_x <= 32'sh26dd3b6a;
      end
    end
    if (result_v_1) begin // @[Reg.scala 17:18]
      if (result_improved) begin // @[Trigonometric.scala 84:14]
        result_nextBestPipe_bits_y <= 32'sh26dd3b6a;
      end else begin
        result_nextBestPipe_bits_y <= 32'sh0;
      end
    end
    if (result_v_1) begin // @[Reg.scala 17:18]
      if (result_improved) begin // @[Trigonometric.scala 84:14]
        result_nextBestPipe_bits_z <= result_nz;
      end else begin
        result_nextBestPipe_bits_z <= 32'sh40000000;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_1 <= result_nextPipe_valid; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_1_x <= _result_nx_T_11;
      end else begin
        result_nextPipe_bits_1_x <= _result_nx_T_15;
      end
    end
    if (result_nextPipe_valid) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_1_y <= _result_ny_T_11;
      end else begin
        result_nextPipe_bits_1_y <= _result_ny_T_15;
      end
    end
    if (result_nextPipe_valid) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_1_z <= _result_nz_T_8;
      end else begin
        result_nextPipe_bits_1_z <= _result_nz_T_11;
      end
    end
    if (result_nextPipe_valid) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_1_sigma <= result_ns_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_1 <= result_nextBestPipe_valid; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid) begin // @[Reg.scala 17:18]
      if (result_improved_1) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_1_x <= _result_nx_T_11;
        end else begin
          result_nextBestPipe_bits_1_x <= _result_nx_T_15;
        end
      end else begin
        result_nextBestPipe_bits_1_x <= result_nextBestPipe_bits_x;
      end
    end
    if (result_nextBestPipe_valid) begin // @[Reg.scala 17:18]
      if (result_improved_1) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_1_y <= _result_ny_T_11;
        end else begin
          result_nextBestPipe_bits_1_y <= _result_ny_T_15;
        end
      end else begin
        result_nextBestPipe_bits_1_y <= result_nextBestPipe_bits_y;
      end
    end
    if (result_nextBestPipe_valid) begin // @[Reg.scala 17:18]
      if (result_improved_1) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_1_z <= _result_nz_T_8;
        end else begin
          result_nextBestPipe_bits_1_z <= _result_nz_T_11;
        end
      end else begin
        result_nextBestPipe_bits_1_z <= result_nextBestPipe_bits_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_2 <= result_nextPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_1) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_1_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_2_x <= _result_nx_T_19;
      end else begin
        result_nextPipe_bits_2_x <= _result_nx_T_23;
      end
    end
    if (result_nextPipe_valid_1) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_1_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_2_y <= _result_ny_T_19;
      end else begin
        result_nextPipe_bits_2_y <= _result_ny_T_23;
      end
    end
    if (result_nextPipe_valid_1) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_1_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_2_z <= _result_nz_T_14;
      end else begin
        result_nextPipe_bits_2_z <= _result_nz_T_17;
      end
    end
    if (result_nextPipe_valid_1) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_2_sigma <= result_ns_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_2 <= result_nextBestPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_1) begin // @[Reg.scala 17:18]
      if (result_improved_2) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_1_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_2_x <= _result_nx_T_19;
        end else begin
          result_nextBestPipe_bits_2_x <= _result_nx_T_23;
        end
      end else begin
        result_nextBestPipe_bits_2_x <= result_nextBestPipe_bits_1_x;
      end
    end
    if (result_nextBestPipe_valid_1) begin // @[Reg.scala 17:18]
      if (result_improved_2) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_1_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_2_y <= _result_ny_T_19;
        end else begin
          result_nextBestPipe_bits_2_y <= _result_ny_T_23;
        end
      end else begin
        result_nextBestPipe_bits_2_y <= result_nextBestPipe_bits_1_y;
      end
    end
    if (result_nextBestPipe_valid_1) begin // @[Reg.scala 17:18]
      if (result_improved_2) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_1_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_2_z <= _result_nz_T_14;
        end else begin
          result_nextBestPipe_bits_2_z <= _result_nz_T_17;
        end
      end else begin
        result_nextBestPipe_bits_2_z <= result_nextBestPipe_bits_1_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_3 <= result_nextPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_2) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_2_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_3_x <= _result_nx_T_27;
      end else begin
        result_nextPipe_bits_3_x <= _result_nx_T_31;
      end
    end
    if (result_nextPipe_valid_2) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_2_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_3_y <= _result_ny_T_27;
      end else begin
        result_nextPipe_bits_3_y <= _result_ny_T_31;
      end
    end
    if (result_nextPipe_valid_2) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_2_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_3_z <= _result_nz_T_20;
      end else begin
        result_nextPipe_bits_3_z <= _result_nz_T_23;
      end
    end
    if (result_nextPipe_valid_2) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_3_sigma <= result_ns_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_3 <= result_nextBestPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_2) begin // @[Reg.scala 17:18]
      if (result_improved_3) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_2_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_3_x <= _result_nx_T_27;
        end else begin
          result_nextBestPipe_bits_3_x <= _result_nx_T_31;
        end
      end else begin
        result_nextBestPipe_bits_3_x <= result_nextBestPipe_bits_2_x;
      end
    end
    if (result_nextBestPipe_valid_2) begin // @[Reg.scala 17:18]
      if (result_improved_3) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_2_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_3_y <= _result_ny_T_27;
        end else begin
          result_nextBestPipe_bits_3_y <= _result_ny_T_31;
        end
      end else begin
        result_nextBestPipe_bits_3_y <= result_nextBestPipe_bits_2_y;
      end
    end
    if (result_nextBestPipe_valid_2) begin // @[Reg.scala 17:18]
      if (result_improved_3) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_2_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_3_z <= _result_nz_T_20;
        end else begin
          result_nextBestPipe_bits_3_z <= _result_nz_T_23;
        end
      end else begin
        result_nextBestPipe_bits_3_z <= result_nextBestPipe_bits_2_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_4 <= result_nextPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_3) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_3_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_4_x <= _result_nx_T_35;
      end else begin
        result_nextPipe_bits_4_x <= _result_nx_T_39;
      end
    end
    if (result_nextPipe_valid_3) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_3_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_4_y <= _result_ny_T_35;
      end else begin
        result_nextPipe_bits_4_y <= _result_ny_T_39;
      end
    end
    if (result_nextPipe_valid_3) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_3_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_4_z <= _result_nz_T_26;
      end else begin
        result_nextPipe_bits_4_z <= _result_nz_T_29;
      end
    end
    if (result_nextPipe_valid_3) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_4_sigma <= result_ns_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_4 <= result_nextBestPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_3) begin // @[Reg.scala 17:18]
      if (result_improved_4) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_3_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_4_x <= _result_nx_T_35;
        end else begin
          result_nextBestPipe_bits_4_x <= _result_nx_T_39;
        end
      end else begin
        result_nextBestPipe_bits_4_x <= result_nextBestPipe_bits_3_x;
      end
    end
    if (result_nextBestPipe_valid_3) begin // @[Reg.scala 17:18]
      if (result_improved_4) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_3_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_4_y <= _result_ny_T_35;
        end else begin
          result_nextBestPipe_bits_4_y <= _result_ny_T_39;
        end
      end else begin
        result_nextBestPipe_bits_4_y <= result_nextBestPipe_bits_3_y;
      end
    end
    if (result_nextBestPipe_valid_3) begin // @[Reg.scala 17:18]
      if (result_improved_4) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_3_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_4_z <= _result_nz_T_26;
        end else begin
          result_nextBestPipe_bits_4_z <= _result_nz_T_29;
        end
      end else begin
        result_nextBestPipe_bits_4_z <= result_nextBestPipe_bits_3_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_5 <= result_nextPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_4) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_4_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_5_x <= _result_nx_T_43;
      end else begin
        result_nextPipe_bits_5_x <= _result_nx_T_47;
      end
    end
    if (result_nextPipe_valid_4) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_4_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_5_y <= _result_ny_T_43;
      end else begin
        result_nextPipe_bits_5_y <= _result_ny_T_47;
      end
    end
    if (result_nextPipe_valid_4) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_4_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_5_z <= _result_nz_T_32;
      end else begin
        result_nextPipe_bits_5_z <= _result_nz_T_35;
      end
    end
    if (result_nextPipe_valid_4) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_5_sigma <= result_ns_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_5 <= result_nextBestPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_4) begin // @[Reg.scala 17:18]
      if (result_improved_5) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_4_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_5_x <= _result_nx_T_43;
        end else begin
          result_nextBestPipe_bits_5_x <= _result_nx_T_47;
        end
      end else begin
        result_nextBestPipe_bits_5_x <= result_nextBestPipe_bits_4_x;
      end
    end
    if (result_nextBestPipe_valid_4) begin // @[Reg.scala 17:18]
      if (result_improved_5) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_4_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_5_y <= _result_ny_T_43;
        end else begin
          result_nextBestPipe_bits_5_y <= _result_ny_T_47;
        end
      end else begin
        result_nextBestPipe_bits_5_y <= result_nextBestPipe_bits_4_y;
      end
    end
    if (result_nextBestPipe_valid_4) begin // @[Reg.scala 17:18]
      if (result_improved_5) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_4_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_5_z <= _result_nz_T_32;
        end else begin
          result_nextBestPipe_bits_5_z <= _result_nz_T_35;
        end
      end else begin
        result_nextBestPipe_bits_5_z <= result_nextBestPipe_bits_4_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_6 <= result_nextPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_5) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_5_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_6_x <= _result_nx_T_51;
      end else begin
        result_nextPipe_bits_6_x <= _result_nx_T_55;
      end
    end
    if (result_nextPipe_valid_5) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_5_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_6_y <= _result_ny_T_51;
      end else begin
        result_nextPipe_bits_6_y <= _result_ny_T_55;
      end
    end
    if (result_nextPipe_valid_5) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_5_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_6_z <= _result_nz_T_38;
      end else begin
        result_nextPipe_bits_6_z <= _result_nz_T_41;
      end
    end
    if (result_nextPipe_valid_5) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_6_sigma <= result_ns_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_6 <= result_nextBestPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_5) begin // @[Reg.scala 17:18]
      if (result_improved_6) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_5_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_6_x <= _result_nx_T_51;
        end else begin
          result_nextBestPipe_bits_6_x <= _result_nx_T_55;
        end
      end else begin
        result_nextBestPipe_bits_6_x <= result_nextBestPipe_bits_5_x;
      end
    end
    if (result_nextBestPipe_valid_5) begin // @[Reg.scala 17:18]
      if (result_improved_6) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_5_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_6_y <= _result_ny_T_51;
        end else begin
          result_nextBestPipe_bits_6_y <= _result_ny_T_55;
        end
      end else begin
        result_nextBestPipe_bits_6_y <= result_nextBestPipe_bits_5_y;
      end
    end
    if (result_nextBestPipe_valid_5) begin // @[Reg.scala 17:18]
      if (result_improved_6) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_5_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_6_z <= _result_nz_T_38;
        end else begin
          result_nextBestPipe_bits_6_z <= _result_nz_T_41;
        end
      end else begin
        result_nextBestPipe_bits_6_z <= result_nextBestPipe_bits_5_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_7 <= result_nextPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_6) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_6_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_7_x <= _result_nx_T_59;
      end else begin
        result_nextPipe_bits_7_x <= _result_nx_T_63;
      end
    end
    if (result_nextPipe_valid_6) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_6_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_7_y <= _result_ny_T_59;
      end else begin
        result_nextPipe_bits_7_y <= _result_ny_T_63;
      end
    end
    if (result_nextPipe_valid_6) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_6_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_7_z <= _result_nz_T_44;
      end else begin
        result_nextPipe_bits_7_z <= _result_nz_T_47;
      end
    end
    if (result_nextPipe_valid_6) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_7_sigma <= result_ns_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_7 <= result_nextBestPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_6) begin // @[Reg.scala 17:18]
      if (result_improved_7) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_6_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_7_x <= _result_nx_T_59;
        end else begin
          result_nextBestPipe_bits_7_x <= _result_nx_T_63;
        end
      end else begin
        result_nextBestPipe_bits_7_x <= result_nextBestPipe_bits_6_x;
      end
    end
    if (result_nextBestPipe_valid_6) begin // @[Reg.scala 17:18]
      if (result_improved_7) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_6_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_7_y <= _result_ny_T_59;
        end else begin
          result_nextBestPipe_bits_7_y <= _result_ny_T_63;
        end
      end else begin
        result_nextBestPipe_bits_7_y <= result_nextBestPipe_bits_6_y;
      end
    end
    if (result_nextBestPipe_valid_6) begin // @[Reg.scala 17:18]
      if (result_improved_7) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_6_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_7_z <= _result_nz_T_44;
        end else begin
          result_nextBestPipe_bits_7_z <= _result_nz_T_47;
        end
      end else begin
        result_nextBestPipe_bits_7_z <= result_nextBestPipe_bits_6_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_8 <= result_nextPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_7) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_7_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_8_x <= _result_nx_T_67;
      end else begin
        result_nextPipe_bits_8_x <= _result_nx_T_71;
      end
    end
    if (result_nextPipe_valid_7) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_7_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_8_y <= _result_ny_T_67;
      end else begin
        result_nextPipe_bits_8_y <= _result_ny_T_71;
      end
    end
    if (result_nextPipe_valid_7) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_7_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_8_z <= _result_nz_T_50;
      end else begin
        result_nextPipe_bits_8_z <= _result_nz_T_53;
      end
    end
    if (result_nextPipe_valid_7) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_8_sigma <= result_ns_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_8 <= result_nextBestPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_7) begin // @[Reg.scala 17:18]
      if (result_improved_8) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_7_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_8_x <= _result_nx_T_67;
        end else begin
          result_nextBestPipe_bits_8_x <= _result_nx_T_71;
        end
      end else begin
        result_nextBestPipe_bits_8_x <= result_nextBestPipe_bits_7_x;
      end
    end
    if (result_nextBestPipe_valid_7) begin // @[Reg.scala 17:18]
      if (result_improved_8) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_7_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_8_y <= _result_ny_T_67;
        end else begin
          result_nextBestPipe_bits_8_y <= _result_ny_T_71;
        end
      end else begin
        result_nextBestPipe_bits_8_y <= result_nextBestPipe_bits_7_y;
      end
    end
    if (result_nextBestPipe_valid_7) begin // @[Reg.scala 17:18]
      if (result_improved_8) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_7_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_8_z <= _result_nz_T_50;
        end else begin
          result_nextBestPipe_bits_8_z <= _result_nz_T_53;
        end
      end else begin
        result_nextBestPipe_bits_8_z <= result_nextBestPipe_bits_7_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_9 <= result_nextPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_8) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_8_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_9_x <= _result_nx_T_75;
      end else begin
        result_nextPipe_bits_9_x <= _result_nx_T_79;
      end
    end
    if (result_nextPipe_valid_8) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_8_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_9_y <= _result_ny_T_75;
      end else begin
        result_nextPipe_bits_9_y <= _result_ny_T_79;
      end
    end
    if (result_nextPipe_valid_8) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_8_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_9_z <= _result_nz_T_56;
      end else begin
        result_nextPipe_bits_9_z <= _result_nz_T_59;
      end
    end
    if (result_nextPipe_valid_8) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_9_sigma <= result_ns_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_9 <= result_nextBestPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_8) begin // @[Reg.scala 17:18]
      if (result_improved_9) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_8_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_9_x <= _result_nx_T_75;
        end else begin
          result_nextBestPipe_bits_9_x <= _result_nx_T_79;
        end
      end else begin
        result_nextBestPipe_bits_9_x <= result_nextBestPipe_bits_8_x;
      end
    end
    if (result_nextBestPipe_valid_8) begin // @[Reg.scala 17:18]
      if (result_improved_9) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_8_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_9_y <= _result_ny_T_75;
        end else begin
          result_nextBestPipe_bits_9_y <= _result_ny_T_79;
        end
      end else begin
        result_nextBestPipe_bits_9_y <= result_nextBestPipe_bits_8_y;
      end
    end
    if (result_nextBestPipe_valid_8) begin // @[Reg.scala 17:18]
      if (result_improved_9) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_8_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_9_z <= _result_nz_T_56;
        end else begin
          result_nextBestPipe_bits_9_z <= _result_nz_T_59;
        end
      end else begin
        result_nextBestPipe_bits_9_z <= result_nextBestPipe_bits_8_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_10 <= result_nextPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_9) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_9_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_10_x <= _result_nx_T_83;
      end else begin
        result_nextPipe_bits_10_x <= _result_nx_T_87;
      end
    end
    if (result_nextPipe_valid_9) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_9_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_10_y <= _result_ny_T_83;
      end else begin
        result_nextPipe_bits_10_y <= _result_ny_T_87;
      end
    end
    if (result_nextPipe_valid_9) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_9_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_10_z <= _result_nz_T_62;
      end else begin
        result_nextPipe_bits_10_z <= _result_nz_T_65;
      end
    end
    if (result_nextPipe_valid_9) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_10_sigma <= result_ns_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_10 <= result_nextBestPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_9) begin // @[Reg.scala 17:18]
      if (result_improved_10) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_9_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_10_x <= _result_nx_T_83;
        end else begin
          result_nextBestPipe_bits_10_x <= _result_nx_T_87;
        end
      end else begin
        result_nextBestPipe_bits_10_x <= result_nextBestPipe_bits_9_x;
      end
    end
    if (result_nextBestPipe_valid_9) begin // @[Reg.scala 17:18]
      if (result_improved_10) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_9_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_10_y <= _result_ny_T_83;
        end else begin
          result_nextBestPipe_bits_10_y <= _result_ny_T_87;
        end
      end else begin
        result_nextBestPipe_bits_10_y <= result_nextBestPipe_bits_9_y;
      end
    end
    if (result_nextBestPipe_valid_9) begin // @[Reg.scala 17:18]
      if (result_improved_10) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_9_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_10_z <= _result_nz_T_62;
        end else begin
          result_nextBestPipe_bits_10_z <= _result_nz_T_65;
        end
      end else begin
        result_nextBestPipe_bits_10_z <= result_nextBestPipe_bits_9_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_11 <= result_nextPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_10) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_10_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_11_x <= _result_nx_T_91;
      end else begin
        result_nextPipe_bits_11_x <= _result_nx_T_95;
      end
    end
    if (result_nextPipe_valid_10) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_10_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_11_y <= _result_ny_T_91;
      end else begin
        result_nextPipe_bits_11_y <= _result_ny_T_95;
      end
    end
    if (result_nextPipe_valid_10) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_10_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_11_z <= _result_nz_T_68;
      end else begin
        result_nextPipe_bits_11_z <= _result_nz_T_71;
      end
    end
    if (result_nextPipe_valid_10) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_11_sigma <= result_ns_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_11 <= result_nextBestPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_10) begin // @[Reg.scala 17:18]
      if (result_improved_11) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_10_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_11_x <= _result_nx_T_91;
        end else begin
          result_nextBestPipe_bits_11_x <= _result_nx_T_95;
        end
      end else begin
        result_nextBestPipe_bits_11_x <= result_nextBestPipe_bits_10_x;
      end
    end
    if (result_nextBestPipe_valid_10) begin // @[Reg.scala 17:18]
      if (result_improved_11) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_10_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_11_y <= _result_ny_T_91;
        end else begin
          result_nextBestPipe_bits_11_y <= _result_ny_T_95;
        end
      end else begin
        result_nextBestPipe_bits_11_y <= result_nextBestPipe_bits_10_y;
      end
    end
    if (result_nextBestPipe_valid_10) begin // @[Reg.scala 17:18]
      if (result_improved_11) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_10_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_11_z <= _result_nz_T_68;
        end else begin
          result_nextBestPipe_bits_11_z <= _result_nz_T_71;
        end
      end else begin
        result_nextBestPipe_bits_11_z <= result_nextBestPipe_bits_10_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_12 <= result_nextPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_11) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_11_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_12_x <= _result_nx_T_99;
      end else begin
        result_nextPipe_bits_12_x <= _result_nx_T_103;
      end
    end
    if (result_nextPipe_valid_11) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_11_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_12_y <= _result_ny_T_99;
      end else begin
        result_nextPipe_bits_12_y <= _result_ny_T_103;
      end
    end
    if (result_nextPipe_valid_11) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_11_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_12_z <= _result_nz_T_74;
      end else begin
        result_nextPipe_bits_12_z <= _result_nz_T_77;
      end
    end
    if (result_nextPipe_valid_11) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_12_sigma <= result_ns_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_12 <= result_nextBestPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_11) begin // @[Reg.scala 17:18]
      if (result_improved_12) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_11_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_12_x <= _result_nx_T_99;
        end else begin
          result_nextBestPipe_bits_12_x <= _result_nx_T_103;
        end
      end else begin
        result_nextBestPipe_bits_12_x <= result_nextBestPipe_bits_11_x;
      end
    end
    if (result_nextBestPipe_valid_11) begin // @[Reg.scala 17:18]
      if (result_improved_12) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_11_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_12_y <= _result_ny_T_99;
        end else begin
          result_nextBestPipe_bits_12_y <= _result_ny_T_103;
        end
      end else begin
        result_nextBestPipe_bits_12_y <= result_nextBestPipe_bits_11_y;
      end
    end
    if (result_nextBestPipe_valid_11) begin // @[Reg.scala 17:18]
      if (result_improved_12) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_11_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_12_z <= _result_nz_T_74;
        end else begin
          result_nextBestPipe_bits_12_z <= _result_nz_T_77;
        end
      end else begin
        result_nextBestPipe_bits_12_z <= result_nextBestPipe_bits_11_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_13 <= result_nextPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_12) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_12_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_13_x <= _result_nx_T_107;
      end else begin
        result_nextPipe_bits_13_x <= _result_nx_T_111;
      end
    end
    if (result_nextPipe_valid_12) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_12_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_13_y <= _result_ny_T_107;
      end else begin
        result_nextPipe_bits_13_y <= _result_ny_T_111;
      end
    end
    if (result_nextPipe_valid_12) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_12_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_13_z <= _result_nz_T_80;
      end else begin
        result_nextPipe_bits_13_z <= _result_nz_T_83;
      end
    end
    if (result_nextPipe_valid_12) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_13_sigma <= result_ns_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_13 <= result_nextBestPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_12) begin // @[Reg.scala 17:18]
      if (result_improved_13) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_12_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_13_x <= _result_nx_T_107;
        end else begin
          result_nextBestPipe_bits_13_x <= _result_nx_T_111;
        end
      end else begin
        result_nextBestPipe_bits_13_x <= result_nextBestPipe_bits_12_x;
      end
    end
    if (result_nextBestPipe_valid_12) begin // @[Reg.scala 17:18]
      if (result_improved_13) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_12_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_13_y <= _result_ny_T_107;
        end else begin
          result_nextBestPipe_bits_13_y <= _result_ny_T_111;
        end
      end else begin
        result_nextBestPipe_bits_13_y <= result_nextBestPipe_bits_12_y;
      end
    end
    if (result_nextBestPipe_valid_12) begin // @[Reg.scala 17:18]
      if (result_improved_13) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_12_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_13_z <= _result_nz_T_80;
        end else begin
          result_nextBestPipe_bits_13_z <= _result_nz_T_83;
        end
      end else begin
        result_nextBestPipe_bits_13_z <= result_nextBestPipe_bits_12_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_14 <= result_nextPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_13) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_13_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_14_x <= _result_nx_T_115;
      end else begin
        result_nextPipe_bits_14_x <= _result_nx_T_119;
      end
    end
    if (result_nextPipe_valid_13) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_13_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_14_y <= _result_ny_T_115;
      end else begin
        result_nextPipe_bits_14_y <= _result_ny_T_119;
      end
    end
    if (result_nextPipe_valid_13) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_13_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_14_z <= _result_nz_T_86;
      end else begin
        result_nextPipe_bits_14_z <= _result_nz_T_89;
      end
    end
    if (result_nextPipe_valid_13) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_14_sigma <= result_ns_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_14 <= result_nextBestPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_13) begin // @[Reg.scala 17:18]
      if (result_improved_14) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_13_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_14_x <= _result_nx_T_115;
        end else begin
          result_nextBestPipe_bits_14_x <= _result_nx_T_119;
        end
      end else begin
        result_nextBestPipe_bits_14_x <= result_nextBestPipe_bits_13_x;
      end
    end
    if (result_nextBestPipe_valid_13) begin // @[Reg.scala 17:18]
      if (result_improved_14) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_13_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_14_y <= _result_ny_T_115;
        end else begin
          result_nextBestPipe_bits_14_y <= _result_ny_T_119;
        end
      end else begin
        result_nextBestPipe_bits_14_y <= result_nextBestPipe_bits_13_y;
      end
    end
    if (result_nextBestPipe_valid_13) begin // @[Reg.scala 17:18]
      if (result_improved_14) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_13_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_14_z <= _result_nz_T_86;
        end else begin
          result_nextBestPipe_bits_14_z <= _result_nz_T_89;
        end
      end else begin
        result_nextBestPipe_bits_14_z <= result_nextBestPipe_bits_13_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_15 <= result_nextPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_14) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_14_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_15_x <= _result_nx_T_123;
      end else begin
        result_nextPipe_bits_15_x <= _result_nx_T_127;
      end
    end
    if (result_nextPipe_valid_14) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_14_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_15_y <= _result_ny_T_123;
      end else begin
        result_nextPipe_bits_15_y <= _result_ny_T_127;
      end
    end
    if (result_nextPipe_valid_14) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_14_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_15_z <= _result_nz_T_92;
      end else begin
        result_nextPipe_bits_15_z <= _result_nz_T_95;
      end
    end
    if (result_nextPipe_valid_14) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_15_sigma <= result_ns_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_15 <= result_nextBestPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_14) begin // @[Reg.scala 17:18]
      if (result_improved_15) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_14_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_15_x <= _result_nx_T_123;
        end else begin
          result_nextBestPipe_bits_15_x <= _result_nx_T_127;
        end
      end else begin
        result_nextBestPipe_bits_15_x <= result_nextBestPipe_bits_14_x;
      end
    end
    if (result_nextBestPipe_valid_14) begin // @[Reg.scala 17:18]
      if (result_improved_15) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_14_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_15_y <= _result_ny_T_123;
        end else begin
          result_nextBestPipe_bits_15_y <= _result_ny_T_127;
        end
      end else begin
        result_nextBestPipe_bits_15_y <= result_nextBestPipe_bits_14_y;
      end
    end
    if (result_nextBestPipe_valid_14) begin // @[Reg.scala 17:18]
      if (result_improved_15) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_14_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_15_z <= _result_nz_T_92;
        end else begin
          result_nextBestPipe_bits_15_z <= _result_nz_T_95;
        end
      end else begin
        result_nextBestPipe_bits_15_z <= result_nextBestPipe_bits_14_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_16 <= result_nextPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_15) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_15_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_16_x <= _result_nx_T_131;
      end else begin
        result_nextPipe_bits_16_x <= _result_nx_T_135;
      end
    end
    if (result_nextPipe_valid_15) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_15_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_16_y <= _result_ny_T_131;
      end else begin
        result_nextPipe_bits_16_y <= _result_ny_T_135;
      end
    end
    if (result_nextPipe_valid_15) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_15_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_16_z <= _result_nz_T_98;
      end else begin
        result_nextPipe_bits_16_z <= _result_nz_T_101;
      end
    end
    if (result_nextPipe_valid_15) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_16_sigma <= result_ns_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_16 <= result_nextBestPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_15) begin // @[Reg.scala 17:18]
      if (result_improved_16) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_15_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_16_x <= _result_nx_T_131;
        end else begin
          result_nextBestPipe_bits_16_x <= _result_nx_T_135;
        end
      end else begin
        result_nextBestPipe_bits_16_x <= result_nextBestPipe_bits_15_x;
      end
    end
    if (result_nextBestPipe_valid_15) begin // @[Reg.scala 17:18]
      if (result_improved_16) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_15_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_16_y <= _result_ny_T_131;
        end else begin
          result_nextBestPipe_bits_16_y <= _result_ny_T_135;
        end
      end else begin
        result_nextBestPipe_bits_16_y <= result_nextBestPipe_bits_15_y;
      end
    end
    if (result_nextBestPipe_valid_15) begin // @[Reg.scala 17:18]
      if (result_improved_16) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_15_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_16_z <= _result_nz_T_98;
        end else begin
          result_nextBestPipe_bits_16_z <= _result_nz_T_101;
        end
      end else begin
        result_nextBestPipe_bits_16_z <= result_nextBestPipe_bits_15_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_17 <= result_nextPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_16) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_16_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_17_x <= _result_nx_T_139;
      end else begin
        result_nextPipe_bits_17_x <= _result_nx_T_143;
      end
    end
    if (result_nextPipe_valid_16) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_16_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_17_y <= _result_ny_T_139;
      end else begin
        result_nextPipe_bits_17_y <= _result_ny_T_143;
      end
    end
    if (result_nextPipe_valid_16) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_16_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_17_z <= _result_nz_T_104;
      end else begin
        result_nextPipe_bits_17_z <= _result_nz_T_107;
      end
    end
    if (result_nextPipe_valid_16) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_17_sigma <= result_ns_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_17 <= result_nextBestPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_16) begin // @[Reg.scala 17:18]
      if (result_improved_17) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_16_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_17_x <= _result_nx_T_139;
        end else begin
          result_nextBestPipe_bits_17_x <= _result_nx_T_143;
        end
      end else begin
        result_nextBestPipe_bits_17_x <= result_nextBestPipe_bits_16_x;
      end
    end
    if (result_nextBestPipe_valid_16) begin // @[Reg.scala 17:18]
      if (result_improved_17) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_16_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_17_y <= _result_ny_T_139;
        end else begin
          result_nextBestPipe_bits_17_y <= _result_ny_T_143;
        end
      end else begin
        result_nextBestPipe_bits_17_y <= result_nextBestPipe_bits_16_y;
      end
    end
    if (result_nextBestPipe_valid_16) begin // @[Reg.scala 17:18]
      if (result_improved_17) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_16_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_17_z <= _result_nz_T_104;
        end else begin
          result_nextBestPipe_bits_17_z <= _result_nz_T_107;
        end
      end else begin
        result_nextBestPipe_bits_17_z <= result_nextBestPipe_bits_16_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_18 <= result_nextPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_17) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_17_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_18_x <= _result_nx_T_147;
      end else begin
        result_nextPipe_bits_18_x <= _result_nx_T_151;
      end
    end
    if (result_nextPipe_valid_17) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_17_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_18_y <= _result_ny_T_147;
      end else begin
        result_nextPipe_bits_18_y <= _result_ny_T_151;
      end
    end
    if (result_nextPipe_valid_17) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_17_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_18_z <= _result_nz_T_110;
      end else begin
        result_nextPipe_bits_18_z <= _result_nz_T_113;
      end
    end
    if (result_nextPipe_valid_17) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_18_sigma <= result_ns_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_18 <= result_nextBestPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_17) begin // @[Reg.scala 17:18]
      if (result_improved_18) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_17_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_18_x <= _result_nx_T_147;
        end else begin
          result_nextBestPipe_bits_18_x <= _result_nx_T_151;
        end
      end else begin
        result_nextBestPipe_bits_18_x <= result_nextBestPipe_bits_17_x;
      end
    end
    if (result_nextBestPipe_valid_17) begin // @[Reg.scala 17:18]
      if (result_improved_18) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_17_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_18_y <= _result_ny_T_147;
        end else begin
          result_nextBestPipe_bits_18_y <= _result_ny_T_151;
        end
      end else begin
        result_nextBestPipe_bits_18_y <= result_nextBestPipe_bits_17_y;
      end
    end
    if (result_nextBestPipe_valid_17) begin // @[Reg.scala 17:18]
      if (result_improved_18) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_17_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_18_z <= _result_nz_T_110;
        end else begin
          result_nextBestPipe_bits_18_z <= _result_nz_T_113;
        end
      end else begin
        result_nextBestPipe_bits_18_z <= result_nextBestPipe_bits_17_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_19 <= result_nextPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_18) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_18_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_19_x <= _result_nx_T_155;
      end else begin
        result_nextPipe_bits_19_x <= _result_nx_T_159;
      end
    end
    if (result_nextPipe_valid_18) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_18_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_19_y <= _result_ny_T_155;
      end else begin
        result_nextPipe_bits_19_y <= _result_ny_T_159;
      end
    end
    if (result_nextPipe_valid_18) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_18_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_19_z <= _result_nz_T_116;
      end else begin
        result_nextPipe_bits_19_z <= _result_nz_T_119;
      end
    end
    if (result_nextPipe_valid_18) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_19_sigma <= result_ns_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_19 <= result_nextBestPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_18) begin // @[Reg.scala 17:18]
      if (result_improved_19) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_18_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_19_x <= _result_nx_T_155;
        end else begin
          result_nextBestPipe_bits_19_x <= _result_nx_T_159;
        end
      end else begin
        result_nextBestPipe_bits_19_x <= result_nextBestPipe_bits_18_x;
      end
    end
    if (result_nextBestPipe_valid_18) begin // @[Reg.scala 17:18]
      if (result_improved_19) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_18_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_19_y <= _result_ny_T_155;
        end else begin
          result_nextBestPipe_bits_19_y <= _result_ny_T_159;
        end
      end else begin
        result_nextBestPipe_bits_19_y <= result_nextBestPipe_bits_18_y;
      end
    end
    if (result_nextBestPipe_valid_18) begin // @[Reg.scala 17:18]
      if (result_improved_19) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_18_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_19_z <= _result_nz_T_116;
        end else begin
          result_nextBestPipe_bits_19_z <= _result_nz_T_119;
        end
      end else begin
        result_nextBestPipe_bits_19_z <= result_nextBestPipe_bits_18_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_20 <= result_nextPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_19) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_19_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_20_x <= _result_nx_T_163;
      end else begin
        result_nextPipe_bits_20_x <= _result_nx_T_167;
      end
    end
    if (result_nextPipe_valid_19) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_19_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_20_y <= _result_ny_T_163;
      end else begin
        result_nextPipe_bits_20_y <= _result_ny_T_167;
      end
    end
    if (result_nextPipe_valid_19) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_19_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_20_z <= _result_nz_T_122;
      end else begin
        result_nextPipe_bits_20_z <= _result_nz_T_125;
      end
    end
    if (result_nextPipe_valid_19) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_20_sigma <= result_ns_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_20 <= result_nextBestPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_19) begin // @[Reg.scala 17:18]
      if (result_improved_20) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_19_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_20_x <= _result_nx_T_163;
        end else begin
          result_nextBestPipe_bits_20_x <= _result_nx_T_167;
        end
      end else begin
        result_nextBestPipe_bits_20_x <= result_nextBestPipe_bits_19_x;
      end
    end
    if (result_nextBestPipe_valid_19) begin // @[Reg.scala 17:18]
      if (result_improved_20) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_19_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_20_y <= _result_ny_T_163;
        end else begin
          result_nextBestPipe_bits_20_y <= _result_ny_T_167;
        end
      end else begin
        result_nextBestPipe_bits_20_y <= result_nextBestPipe_bits_19_y;
      end
    end
    if (result_nextBestPipe_valid_19) begin // @[Reg.scala 17:18]
      if (result_improved_20) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_19_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_20_z <= _result_nz_T_122;
        end else begin
          result_nextBestPipe_bits_20_z <= _result_nz_T_125;
        end
      end else begin
        result_nextBestPipe_bits_20_z <= result_nextBestPipe_bits_19_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_21 <= result_nextPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_20) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_20_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_21_x <= _result_nx_T_171;
      end else begin
        result_nextPipe_bits_21_x <= _result_nx_T_175;
      end
    end
    if (result_nextPipe_valid_20) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_20_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_21_y <= _result_ny_T_171;
      end else begin
        result_nextPipe_bits_21_y <= _result_ny_T_175;
      end
    end
    if (result_nextPipe_valid_20) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_20_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_21_z <= _result_nz_T_128;
      end else begin
        result_nextPipe_bits_21_z <= _result_nz_T_131;
      end
    end
    if (result_nextPipe_valid_20) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_21_sigma <= result_ns_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_21 <= result_nextBestPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_20) begin // @[Reg.scala 17:18]
      if (result_improved_21) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_20_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_21_x <= _result_nx_T_171;
        end else begin
          result_nextBestPipe_bits_21_x <= _result_nx_T_175;
        end
      end else begin
        result_nextBestPipe_bits_21_x <= result_nextBestPipe_bits_20_x;
      end
    end
    if (result_nextBestPipe_valid_20) begin // @[Reg.scala 17:18]
      if (result_improved_21) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_20_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_21_y <= _result_ny_T_171;
        end else begin
          result_nextBestPipe_bits_21_y <= _result_ny_T_175;
        end
      end else begin
        result_nextBestPipe_bits_21_y <= result_nextBestPipe_bits_20_y;
      end
    end
    if (result_nextBestPipe_valid_20) begin // @[Reg.scala 17:18]
      if (result_improved_21) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_20_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_21_z <= _result_nz_T_128;
        end else begin
          result_nextBestPipe_bits_21_z <= _result_nz_T_131;
        end
      end else begin
        result_nextBestPipe_bits_21_z <= result_nextBestPipe_bits_20_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_22 <= result_nextPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_21) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_21_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_22_x <= _result_nx_T_179;
      end else begin
        result_nextPipe_bits_22_x <= _result_nx_T_183;
      end
    end
    if (result_nextPipe_valid_21) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_21_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_22_y <= _result_ny_T_179;
      end else begin
        result_nextPipe_bits_22_y <= _result_ny_T_183;
      end
    end
    if (result_nextPipe_valid_21) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_21_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_22_z <= _result_nz_T_134;
      end else begin
        result_nextPipe_bits_22_z <= _result_nz_T_137;
      end
    end
    if (result_nextPipe_valid_21) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_22_sigma <= result_ns_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_22 <= result_nextBestPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_21) begin // @[Reg.scala 17:18]
      if (result_improved_22) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_21_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_22_x <= _result_nx_T_179;
        end else begin
          result_nextBestPipe_bits_22_x <= _result_nx_T_183;
        end
      end else begin
        result_nextBestPipe_bits_22_x <= result_nextBestPipe_bits_21_x;
      end
    end
    if (result_nextBestPipe_valid_21) begin // @[Reg.scala 17:18]
      if (result_improved_22) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_21_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_22_y <= _result_ny_T_179;
        end else begin
          result_nextBestPipe_bits_22_y <= _result_ny_T_183;
        end
      end else begin
        result_nextBestPipe_bits_22_y <= result_nextBestPipe_bits_21_y;
      end
    end
    if (result_nextBestPipe_valid_21) begin // @[Reg.scala 17:18]
      if (result_improved_22) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_21_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_22_z <= _result_nz_T_134;
        end else begin
          result_nextBestPipe_bits_22_z <= _result_nz_T_137;
        end
      end else begin
        result_nextBestPipe_bits_22_z <= result_nextBestPipe_bits_21_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_23 <= result_nextPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_22) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_22_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_23_x <= _result_nx_T_187;
      end else begin
        result_nextPipe_bits_23_x <= _result_nx_T_191;
      end
    end
    if (result_nextPipe_valid_22) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_22_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_23_y <= _result_ny_T_187;
      end else begin
        result_nextPipe_bits_23_y <= _result_ny_T_191;
      end
    end
    if (result_nextPipe_valid_22) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_22_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_23_z <= _result_nz_T_140;
      end else begin
        result_nextPipe_bits_23_z <= _result_nz_T_143;
      end
    end
    if (result_nextPipe_valid_22) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_23_sigma <= result_ns_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_23 <= result_nextBestPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_22) begin // @[Reg.scala 17:18]
      if (result_improved_23) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_22_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_23_x <= _result_nx_T_187;
        end else begin
          result_nextBestPipe_bits_23_x <= _result_nx_T_191;
        end
      end else begin
        result_nextBestPipe_bits_23_x <= result_nextBestPipe_bits_22_x;
      end
    end
    if (result_nextBestPipe_valid_22) begin // @[Reg.scala 17:18]
      if (result_improved_23) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_22_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_23_y <= _result_ny_T_187;
        end else begin
          result_nextBestPipe_bits_23_y <= _result_ny_T_191;
        end
      end else begin
        result_nextBestPipe_bits_23_y <= result_nextBestPipe_bits_22_y;
      end
    end
    if (result_nextBestPipe_valid_22) begin // @[Reg.scala 17:18]
      if (result_improved_23) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_22_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_23_z <= _result_nz_T_140;
        end else begin
          result_nextBestPipe_bits_23_z <= _result_nz_T_143;
        end
      end else begin
        result_nextBestPipe_bits_23_z <= result_nextBestPipe_bits_22_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_24 <= result_nextPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_23) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_23_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_24_x <= _result_nx_T_195;
      end else begin
        result_nextPipe_bits_24_x <= _result_nx_T_199;
      end
    end
    if (result_nextPipe_valid_23) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_23_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_24_y <= _result_ny_T_195;
      end else begin
        result_nextPipe_bits_24_y <= _result_ny_T_199;
      end
    end
    if (result_nextPipe_valid_23) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_23_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_24_z <= _result_nz_T_146;
      end else begin
        result_nextPipe_bits_24_z <= _result_nz_T_149;
      end
    end
    if (result_nextPipe_valid_23) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_24_sigma <= result_ns_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_24 <= result_nextBestPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_23) begin // @[Reg.scala 17:18]
      if (result_improved_24) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_23_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_24_x <= _result_nx_T_195;
        end else begin
          result_nextBestPipe_bits_24_x <= _result_nx_T_199;
        end
      end else begin
        result_nextBestPipe_bits_24_x <= result_nextBestPipe_bits_23_x;
      end
    end
    if (result_nextBestPipe_valid_23) begin // @[Reg.scala 17:18]
      if (result_improved_24) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_23_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_24_y <= _result_ny_T_195;
        end else begin
          result_nextBestPipe_bits_24_y <= _result_ny_T_199;
        end
      end else begin
        result_nextBestPipe_bits_24_y <= result_nextBestPipe_bits_23_y;
      end
    end
    if (result_nextBestPipe_valid_23) begin // @[Reg.scala 17:18]
      if (result_improved_24) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_23_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_24_z <= _result_nz_T_146;
        end else begin
          result_nextBestPipe_bits_24_z <= _result_nz_T_149;
        end
      end else begin
        result_nextBestPipe_bits_24_z <= result_nextBestPipe_bits_23_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_25 <= result_nextPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_24) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_24_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_25_x <= _result_nx_T_203;
      end else begin
        result_nextPipe_bits_25_x <= _result_nx_T_207;
      end
    end
    if (result_nextPipe_valid_24) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_24_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_25_y <= _result_ny_T_203;
      end else begin
        result_nextPipe_bits_25_y <= _result_ny_T_207;
      end
    end
    if (result_nextPipe_valid_24) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_24_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_25_z <= _result_nz_T_152;
      end else begin
        result_nextPipe_bits_25_z <= _result_nz_T_155;
      end
    end
    if (result_nextPipe_valid_24) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_25_sigma <= result_ns_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_25 <= result_nextBestPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_24) begin // @[Reg.scala 17:18]
      if (result_improved_25) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_24_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_25_x <= _result_nx_T_203;
        end else begin
          result_nextBestPipe_bits_25_x <= _result_nx_T_207;
        end
      end else begin
        result_nextBestPipe_bits_25_x <= result_nextBestPipe_bits_24_x;
      end
    end
    if (result_nextBestPipe_valid_24) begin // @[Reg.scala 17:18]
      if (result_improved_25) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_24_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_25_y <= _result_ny_T_203;
        end else begin
          result_nextBestPipe_bits_25_y <= _result_ny_T_207;
        end
      end else begin
        result_nextBestPipe_bits_25_y <= result_nextBestPipe_bits_24_y;
      end
    end
    if (result_nextBestPipe_valid_24) begin // @[Reg.scala 17:18]
      if (result_improved_25) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_24_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_25_z <= _result_nz_T_152;
        end else begin
          result_nextBestPipe_bits_25_z <= _result_nz_T_155;
        end
      end else begin
        result_nextBestPipe_bits_25_z <= result_nextBestPipe_bits_24_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_26 <= result_nextPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_25) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_25_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_26_x <= _result_nx_T_211;
      end else begin
        result_nextPipe_bits_26_x <= _result_nx_T_215;
      end
    end
    if (result_nextPipe_valid_25) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_25_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_26_y <= _result_ny_T_211;
      end else begin
        result_nextPipe_bits_26_y <= _result_ny_T_215;
      end
    end
    if (result_nextPipe_valid_25) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_25_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_26_z <= _result_nz_T_158;
      end else begin
        result_nextPipe_bits_26_z <= _result_nz_T_161;
      end
    end
    if (result_nextPipe_valid_25) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_26_sigma <= result_ns_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_26 <= result_nextBestPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_25) begin // @[Reg.scala 17:18]
      if (result_improved_26) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_25_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_26_x <= _result_nx_T_211;
        end else begin
          result_nextBestPipe_bits_26_x <= _result_nx_T_215;
        end
      end else begin
        result_nextBestPipe_bits_26_x <= result_nextBestPipe_bits_25_x;
      end
    end
    if (result_nextBestPipe_valid_25) begin // @[Reg.scala 17:18]
      if (result_improved_26) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_25_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_26_y <= _result_ny_T_211;
        end else begin
          result_nextBestPipe_bits_26_y <= _result_ny_T_215;
        end
      end else begin
        result_nextBestPipe_bits_26_y <= result_nextBestPipe_bits_25_y;
      end
    end
    if (result_nextBestPipe_valid_25) begin // @[Reg.scala 17:18]
      if (result_improved_26) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_25_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_26_z <= _result_nz_T_158;
        end else begin
          result_nextBestPipe_bits_26_z <= _result_nz_T_161;
        end
      end else begin
        result_nextBestPipe_bits_26_z <= result_nextBestPipe_bits_25_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_27 <= result_nextPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_26) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_26_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_27_x <= _result_nx_T_219;
      end else begin
        result_nextPipe_bits_27_x <= _result_nx_T_223;
      end
    end
    if (result_nextPipe_valid_26) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_26_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_27_y <= _result_ny_T_219;
      end else begin
        result_nextPipe_bits_27_y <= _result_ny_T_223;
      end
    end
    if (result_nextPipe_valid_26) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_26_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_27_z <= _result_nz_T_164;
      end else begin
        result_nextPipe_bits_27_z <= _result_nz_T_167;
      end
    end
    if (result_nextPipe_valid_26) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_27_sigma <= result_ns_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_27 <= result_nextBestPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_26) begin // @[Reg.scala 17:18]
      if (result_improved_27) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_26_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_27_x <= _result_nx_T_219;
        end else begin
          result_nextBestPipe_bits_27_x <= _result_nx_T_223;
        end
      end else begin
        result_nextBestPipe_bits_27_x <= result_nextBestPipe_bits_26_x;
      end
    end
    if (result_nextBestPipe_valid_26) begin // @[Reg.scala 17:18]
      if (result_improved_27) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_26_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_27_y <= _result_ny_T_219;
        end else begin
          result_nextBestPipe_bits_27_y <= _result_ny_T_223;
        end
      end else begin
        result_nextBestPipe_bits_27_y <= result_nextBestPipe_bits_26_y;
      end
    end
    if (result_nextBestPipe_valid_26) begin // @[Reg.scala 17:18]
      if (result_improved_27) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_26_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_27_z <= _result_nz_T_164;
        end else begin
          result_nextBestPipe_bits_27_z <= _result_nz_T_167;
        end
      end else begin
        result_nextBestPipe_bits_27_z <= result_nextBestPipe_bits_26_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_28 <= result_nextPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_27) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_27_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_28_x <= _result_nx_T_227;
      end else begin
        result_nextPipe_bits_28_x <= _result_nx_T_231;
      end
    end
    if (result_nextPipe_valid_27) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_27_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_28_y <= _result_ny_T_227;
      end else begin
        result_nextPipe_bits_28_y <= _result_ny_T_231;
      end
    end
    if (result_nextPipe_valid_27) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_27_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_28_z <= _result_nz_T_170;
      end else begin
        result_nextPipe_bits_28_z <= _result_nz_T_173;
      end
    end
    if (result_nextPipe_valid_27) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_28_sigma <= result_ns_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_28 <= result_nextBestPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_27) begin // @[Reg.scala 17:18]
      if (result_improved_28) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_27_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_28_x <= _result_nx_T_227;
        end else begin
          result_nextBestPipe_bits_28_x <= _result_nx_T_231;
        end
      end else begin
        result_nextBestPipe_bits_28_x <= result_nextBestPipe_bits_27_x;
      end
    end
    if (result_nextBestPipe_valid_27) begin // @[Reg.scala 17:18]
      if (result_improved_28) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_27_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_28_y <= _result_ny_T_227;
        end else begin
          result_nextBestPipe_bits_28_y <= _result_ny_T_231;
        end
      end else begin
        result_nextBestPipe_bits_28_y <= result_nextBestPipe_bits_27_y;
      end
    end
    if (result_nextBestPipe_valid_27) begin // @[Reg.scala 17:18]
      if (result_improved_28) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_27_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_28_z <= _result_nz_T_170;
        end else begin
          result_nextBestPipe_bits_28_z <= _result_nz_T_173;
        end
      end else begin
        result_nextBestPipe_bits_28_z <= result_nextBestPipe_bits_27_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextPipe_valid_29 <= result_nextPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (result_nextPipe_valid_28) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_28_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_29_x <= _result_nx_T_235;
      end else begin
        result_nextPipe_bits_29_x <= _result_nx_T_239;
      end
    end
    if (result_nextPipe_valid_28) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_28_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_29_y <= _result_ny_T_235;
      end else begin
        result_nextPipe_bits_29_y <= _result_ny_T_239;
      end
    end
    if (result_nextPipe_valid_28) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_28_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_29_z <= _result_nz_T_176;
      end else begin
        result_nextPipe_bits_29_z <= _result_nz_T_179;
      end
    end
    if (result_nextPipe_valid_28) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_29_sigma <= result_ns_29; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_29 <= result_nextBestPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_28) begin // @[Reg.scala 17:18]
      if (result_improved_29) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_28_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_29_x <= _result_nx_T_235;
        end else begin
          result_nextBestPipe_bits_29_x <= _result_nx_T_239;
        end
      end else begin
        result_nextBestPipe_bits_29_x <= result_nextBestPipe_bits_28_x;
      end
    end
    if (result_nextBestPipe_valid_28) begin // @[Reg.scala 17:18]
      if (result_improved_29) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_28_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_29_y <= _result_ny_T_235;
        end else begin
          result_nextBestPipe_bits_29_y <= _result_ny_T_239;
        end
      end else begin
        result_nextBestPipe_bits_29_y <= result_nextBestPipe_bits_28_y;
      end
    end
    if (result_nextBestPipe_valid_28) begin // @[Reg.scala 17:18]
      if (result_improved_29) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_28_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_29_z <= _result_nz_T_176;
        end else begin
          result_nextBestPipe_bits_29_z <= _result_nz_T_179;
        end
      end else begin
        result_nextBestPipe_bits_29_z <= result_nextBestPipe_bits_28_z;
      end
    end
    if (result_nextPipe_valid_29) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_29_sigma) begin // @[Trigonometric.scala 67:24]
        result_nextPipe_bits_30_x <= _result_nx_T_243;
      end else begin
        result_nextPipe_bits_30_x <= _result_nx_T_247;
      end
    end
    if (result_nextPipe_valid_29) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_29_sigma) begin // @[Trigonometric.scala 68:24]
        result_nextPipe_bits_30_y <= _result_ny_T_243;
      end else begin
        result_nextPipe_bits_30_y <= _result_ny_T_247;
      end
    end
    if (result_nextPipe_valid_29) begin // @[Reg.scala 17:18]
      if (result_nextPipe_bits_29_sigma) begin // @[Trigonometric.scala 71:21]
        result_nextPipe_bits_30_z <= _result_nz_T_182;
      end else begin
        result_nextPipe_bits_30_z <= _result_nz_T_185;
      end
    end
    if (result_nextPipe_valid_29) begin // @[Reg.scala 17:18]
      result_nextPipe_bits_30_sigma <= result_ns_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_nextBestPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_nextBestPipe_valid_30 <= result_nextBestPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_29) begin // @[Reg.scala 17:18]
      if (result_improved_30) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_29_sigma) begin // @[Trigonometric.scala 67:24]
          result_nextBestPipe_bits_30_x <= _result_nx_T_243;
        end else begin
          result_nextBestPipe_bits_30_x <= _result_nx_T_247;
        end
      end else begin
        result_nextBestPipe_bits_30_x <= result_nextBestPipe_bits_29_x;
      end
    end
    if (result_nextBestPipe_valid_29) begin // @[Reg.scala 17:18]
      if (result_improved_30) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_29_sigma) begin // @[Trigonometric.scala 68:24]
          result_nextBestPipe_bits_30_y <= _result_ny_T_243;
        end else begin
          result_nextBestPipe_bits_30_y <= _result_ny_T_247;
        end
      end else begin
        result_nextBestPipe_bits_30_y <= result_nextBestPipe_bits_29_y;
      end
    end
    if (result_nextBestPipe_valid_29) begin // @[Reg.scala 17:18]
      if (result_improved_30) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_29_sigma) begin // @[Trigonometric.scala 71:21]
          result_nextBestPipe_bits_30_z <= _result_nz_T_182;
        end else begin
          result_nextBestPipe_bits_30_z <= _result_nz_T_185;
        end
      end else begin
        result_nextBestPipe_bits_30_z <= result_nextBestPipe_bits_29_z;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      resultPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      resultPipe_valid <= result_nextBestPipe_valid_30; // @[Valid.scala 127:22]
    end
    if (result_nextBestPipe_valid_30) begin // @[Reg.scala 17:18]
      if (result_improved_31) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_30_sigma) begin // @[Trigonometric.scala 67:24]
          resultPipe_bits_x <= _result_nx_T_251;
        end else begin
          resultPipe_bits_x <= _result_nx_T_255;
        end
      end else begin
        resultPipe_bits_x <= result_nextBestPipe_bits_30_x;
      end
    end
    if (result_nextBestPipe_valid_30) begin // @[Reg.scala 17:18]
      if (result_improved_31) begin // @[Trigonometric.scala 84:14]
        if (result_nextPipe_bits_30_sigma) begin // @[Trigonometric.scala 68:24]
          resultPipe_bits_y <= _result_ny_T_251;
        end else begin
          resultPipe_bits_y <= _result_ny_T_255;
        end
      end else begin
        resultPipe_bits_y <= result_nextBestPipe_bits_30_y;
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  result_v = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  result_b_z = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  result_v_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  result_nextPipe_valid = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  result_nextPipe_bits_x = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  result_nextPipe_bits_z = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  result_nextPipe_bits_sigma = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  result_nextBestPipe_valid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  result_nextBestPipe_bits_x = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  result_nextBestPipe_bits_y = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  result_nextBestPipe_bits_z = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  result_nextPipe_valid_1 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  result_nextPipe_bits_1_x = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  result_nextPipe_bits_1_y = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  result_nextPipe_bits_1_z = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  result_nextPipe_bits_1_sigma = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  result_nextBestPipe_valid_1 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  result_nextBestPipe_bits_1_x = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  result_nextBestPipe_bits_1_y = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  result_nextBestPipe_bits_1_z = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  result_nextPipe_valid_2 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  result_nextPipe_bits_2_x = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  result_nextPipe_bits_2_y = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  result_nextPipe_bits_2_z = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  result_nextPipe_bits_2_sigma = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  result_nextBestPipe_valid_2 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  result_nextBestPipe_bits_2_x = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  result_nextBestPipe_bits_2_y = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  result_nextBestPipe_bits_2_z = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  result_nextPipe_valid_3 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  result_nextPipe_bits_3_x = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  result_nextPipe_bits_3_y = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  result_nextPipe_bits_3_z = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  result_nextPipe_bits_3_sigma = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  result_nextBestPipe_valid_3 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  result_nextBestPipe_bits_3_x = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  result_nextBestPipe_bits_3_y = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  result_nextBestPipe_bits_3_z = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  result_nextPipe_valid_4 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  result_nextPipe_bits_4_x = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  result_nextPipe_bits_4_y = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  result_nextPipe_bits_4_z = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  result_nextPipe_bits_4_sigma = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  result_nextBestPipe_valid_4 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  result_nextBestPipe_bits_4_x = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  result_nextBestPipe_bits_4_y = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  result_nextBestPipe_bits_4_z = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  result_nextPipe_valid_5 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  result_nextPipe_bits_5_x = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  result_nextPipe_bits_5_y = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  result_nextPipe_bits_5_z = _RAND_50[31:0];
  _RAND_51 = {1{`RANDOM}};
  result_nextPipe_bits_5_sigma = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  result_nextBestPipe_valid_5 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  result_nextBestPipe_bits_5_x = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  result_nextBestPipe_bits_5_y = _RAND_54[31:0];
  _RAND_55 = {1{`RANDOM}};
  result_nextBestPipe_bits_5_z = _RAND_55[31:0];
  _RAND_56 = {1{`RANDOM}};
  result_nextPipe_valid_6 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  result_nextPipe_bits_6_x = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  result_nextPipe_bits_6_y = _RAND_58[31:0];
  _RAND_59 = {1{`RANDOM}};
  result_nextPipe_bits_6_z = _RAND_59[31:0];
  _RAND_60 = {1{`RANDOM}};
  result_nextPipe_bits_6_sigma = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  result_nextBestPipe_valid_6 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  result_nextBestPipe_bits_6_x = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  result_nextBestPipe_bits_6_y = _RAND_63[31:0];
  _RAND_64 = {1{`RANDOM}};
  result_nextBestPipe_bits_6_z = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  result_nextPipe_valid_7 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  result_nextPipe_bits_7_x = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  result_nextPipe_bits_7_y = _RAND_67[31:0];
  _RAND_68 = {1{`RANDOM}};
  result_nextPipe_bits_7_z = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  result_nextPipe_bits_7_sigma = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  result_nextBestPipe_valid_7 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  result_nextBestPipe_bits_7_x = _RAND_71[31:0];
  _RAND_72 = {1{`RANDOM}};
  result_nextBestPipe_bits_7_y = _RAND_72[31:0];
  _RAND_73 = {1{`RANDOM}};
  result_nextBestPipe_bits_7_z = _RAND_73[31:0];
  _RAND_74 = {1{`RANDOM}};
  result_nextPipe_valid_8 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  result_nextPipe_bits_8_x = _RAND_75[31:0];
  _RAND_76 = {1{`RANDOM}};
  result_nextPipe_bits_8_y = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  result_nextPipe_bits_8_z = _RAND_77[31:0];
  _RAND_78 = {1{`RANDOM}};
  result_nextPipe_bits_8_sigma = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  result_nextBestPipe_valid_8 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  result_nextBestPipe_bits_8_x = _RAND_80[31:0];
  _RAND_81 = {1{`RANDOM}};
  result_nextBestPipe_bits_8_y = _RAND_81[31:0];
  _RAND_82 = {1{`RANDOM}};
  result_nextBestPipe_bits_8_z = _RAND_82[31:0];
  _RAND_83 = {1{`RANDOM}};
  result_nextPipe_valid_9 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  result_nextPipe_bits_9_x = _RAND_84[31:0];
  _RAND_85 = {1{`RANDOM}};
  result_nextPipe_bits_9_y = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  result_nextPipe_bits_9_z = _RAND_86[31:0];
  _RAND_87 = {1{`RANDOM}};
  result_nextPipe_bits_9_sigma = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  result_nextBestPipe_valid_9 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  result_nextBestPipe_bits_9_x = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  result_nextBestPipe_bits_9_y = _RAND_90[31:0];
  _RAND_91 = {1{`RANDOM}};
  result_nextBestPipe_bits_9_z = _RAND_91[31:0];
  _RAND_92 = {1{`RANDOM}};
  result_nextPipe_valid_10 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  result_nextPipe_bits_10_x = _RAND_93[31:0];
  _RAND_94 = {1{`RANDOM}};
  result_nextPipe_bits_10_y = _RAND_94[31:0];
  _RAND_95 = {1{`RANDOM}};
  result_nextPipe_bits_10_z = _RAND_95[31:0];
  _RAND_96 = {1{`RANDOM}};
  result_nextPipe_bits_10_sigma = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  result_nextBestPipe_valid_10 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  result_nextBestPipe_bits_10_x = _RAND_98[31:0];
  _RAND_99 = {1{`RANDOM}};
  result_nextBestPipe_bits_10_y = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  result_nextBestPipe_bits_10_z = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  result_nextPipe_valid_11 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  result_nextPipe_bits_11_x = _RAND_102[31:0];
  _RAND_103 = {1{`RANDOM}};
  result_nextPipe_bits_11_y = _RAND_103[31:0];
  _RAND_104 = {1{`RANDOM}};
  result_nextPipe_bits_11_z = _RAND_104[31:0];
  _RAND_105 = {1{`RANDOM}};
  result_nextPipe_bits_11_sigma = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  result_nextBestPipe_valid_11 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  result_nextBestPipe_bits_11_x = _RAND_107[31:0];
  _RAND_108 = {1{`RANDOM}};
  result_nextBestPipe_bits_11_y = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  result_nextBestPipe_bits_11_z = _RAND_109[31:0];
  _RAND_110 = {1{`RANDOM}};
  result_nextPipe_valid_12 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  result_nextPipe_bits_12_x = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  result_nextPipe_bits_12_y = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  result_nextPipe_bits_12_z = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  result_nextPipe_bits_12_sigma = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  result_nextBestPipe_valid_12 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  result_nextBestPipe_bits_12_x = _RAND_116[31:0];
  _RAND_117 = {1{`RANDOM}};
  result_nextBestPipe_bits_12_y = _RAND_117[31:0];
  _RAND_118 = {1{`RANDOM}};
  result_nextBestPipe_bits_12_z = _RAND_118[31:0];
  _RAND_119 = {1{`RANDOM}};
  result_nextPipe_valid_13 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  result_nextPipe_bits_13_x = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  result_nextPipe_bits_13_y = _RAND_121[31:0];
  _RAND_122 = {1{`RANDOM}};
  result_nextPipe_bits_13_z = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  result_nextPipe_bits_13_sigma = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  result_nextBestPipe_valid_13 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  result_nextBestPipe_bits_13_x = _RAND_125[31:0];
  _RAND_126 = {1{`RANDOM}};
  result_nextBestPipe_bits_13_y = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  result_nextBestPipe_bits_13_z = _RAND_127[31:0];
  _RAND_128 = {1{`RANDOM}};
  result_nextPipe_valid_14 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  result_nextPipe_bits_14_x = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  result_nextPipe_bits_14_y = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  result_nextPipe_bits_14_z = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  result_nextPipe_bits_14_sigma = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  result_nextBestPipe_valid_14 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  result_nextBestPipe_bits_14_x = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  result_nextBestPipe_bits_14_y = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  result_nextBestPipe_bits_14_z = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  result_nextPipe_valid_15 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  result_nextPipe_bits_15_x = _RAND_138[31:0];
  _RAND_139 = {1{`RANDOM}};
  result_nextPipe_bits_15_y = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  result_nextPipe_bits_15_z = _RAND_140[31:0];
  _RAND_141 = {1{`RANDOM}};
  result_nextPipe_bits_15_sigma = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  result_nextBestPipe_valid_15 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  result_nextBestPipe_bits_15_x = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  result_nextBestPipe_bits_15_y = _RAND_144[31:0];
  _RAND_145 = {1{`RANDOM}};
  result_nextBestPipe_bits_15_z = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  result_nextPipe_valid_16 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  result_nextPipe_bits_16_x = _RAND_147[31:0];
  _RAND_148 = {1{`RANDOM}};
  result_nextPipe_bits_16_y = _RAND_148[31:0];
  _RAND_149 = {1{`RANDOM}};
  result_nextPipe_bits_16_z = _RAND_149[31:0];
  _RAND_150 = {1{`RANDOM}};
  result_nextPipe_bits_16_sigma = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  result_nextBestPipe_valid_16 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  result_nextBestPipe_bits_16_x = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  result_nextBestPipe_bits_16_y = _RAND_153[31:0];
  _RAND_154 = {1{`RANDOM}};
  result_nextBestPipe_bits_16_z = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  result_nextPipe_valid_17 = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  result_nextPipe_bits_17_x = _RAND_156[31:0];
  _RAND_157 = {1{`RANDOM}};
  result_nextPipe_bits_17_y = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  result_nextPipe_bits_17_z = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  result_nextPipe_bits_17_sigma = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  result_nextBestPipe_valid_17 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  result_nextBestPipe_bits_17_x = _RAND_161[31:0];
  _RAND_162 = {1{`RANDOM}};
  result_nextBestPipe_bits_17_y = _RAND_162[31:0];
  _RAND_163 = {1{`RANDOM}};
  result_nextBestPipe_bits_17_z = _RAND_163[31:0];
  _RAND_164 = {1{`RANDOM}};
  result_nextPipe_valid_18 = _RAND_164[0:0];
  _RAND_165 = {1{`RANDOM}};
  result_nextPipe_bits_18_x = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  result_nextPipe_bits_18_y = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  result_nextPipe_bits_18_z = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  result_nextPipe_bits_18_sigma = _RAND_168[0:0];
  _RAND_169 = {1{`RANDOM}};
  result_nextBestPipe_valid_18 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  result_nextBestPipe_bits_18_x = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  result_nextBestPipe_bits_18_y = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  result_nextBestPipe_bits_18_z = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  result_nextPipe_valid_19 = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  result_nextPipe_bits_19_x = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  result_nextPipe_bits_19_y = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  result_nextPipe_bits_19_z = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  result_nextPipe_bits_19_sigma = _RAND_177[0:0];
  _RAND_178 = {1{`RANDOM}};
  result_nextBestPipe_valid_19 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  result_nextBestPipe_bits_19_x = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  result_nextBestPipe_bits_19_y = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  result_nextBestPipe_bits_19_z = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  result_nextPipe_valid_20 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  result_nextPipe_bits_20_x = _RAND_183[31:0];
  _RAND_184 = {1{`RANDOM}};
  result_nextPipe_bits_20_y = _RAND_184[31:0];
  _RAND_185 = {1{`RANDOM}};
  result_nextPipe_bits_20_z = _RAND_185[31:0];
  _RAND_186 = {1{`RANDOM}};
  result_nextPipe_bits_20_sigma = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  result_nextBestPipe_valid_20 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  result_nextBestPipe_bits_20_x = _RAND_188[31:0];
  _RAND_189 = {1{`RANDOM}};
  result_nextBestPipe_bits_20_y = _RAND_189[31:0];
  _RAND_190 = {1{`RANDOM}};
  result_nextBestPipe_bits_20_z = _RAND_190[31:0];
  _RAND_191 = {1{`RANDOM}};
  result_nextPipe_valid_21 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  result_nextPipe_bits_21_x = _RAND_192[31:0];
  _RAND_193 = {1{`RANDOM}};
  result_nextPipe_bits_21_y = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  result_nextPipe_bits_21_z = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  result_nextPipe_bits_21_sigma = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  result_nextBestPipe_valid_21 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  result_nextBestPipe_bits_21_x = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  result_nextBestPipe_bits_21_y = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  result_nextBestPipe_bits_21_z = _RAND_199[31:0];
  _RAND_200 = {1{`RANDOM}};
  result_nextPipe_valid_22 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  result_nextPipe_bits_22_x = _RAND_201[31:0];
  _RAND_202 = {1{`RANDOM}};
  result_nextPipe_bits_22_y = _RAND_202[31:0];
  _RAND_203 = {1{`RANDOM}};
  result_nextPipe_bits_22_z = _RAND_203[31:0];
  _RAND_204 = {1{`RANDOM}};
  result_nextPipe_bits_22_sigma = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  result_nextBestPipe_valid_22 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  result_nextBestPipe_bits_22_x = _RAND_206[31:0];
  _RAND_207 = {1{`RANDOM}};
  result_nextBestPipe_bits_22_y = _RAND_207[31:0];
  _RAND_208 = {1{`RANDOM}};
  result_nextBestPipe_bits_22_z = _RAND_208[31:0];
  _RAND_209 = {1{`RANDOM}};
  result_nextPipe_valid_23 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  result_nextPipe_bits_23_x = _RAND_210[31:0];
  _RAND_211 = {1{`RANDOM}};
  result_nextPipe_bits_23_y = _RAND_211[31:0];
  _RAND_212 = {1{`RANDOM}};
  result_nextPipe_bits_23_z = _RAND_212[31:0];
  _RAND_213 = {1{`RANDOM}};
  result_nextPipe_bits_23_sigma = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  result_nextBestPipe_valid_23 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  result_nextBestPipe_bits_23_x = _RAND_215[31:0];
  _RAND_216 = {1{`RANDOM}};
  result_nextBestPipe_bits_23_y = _RAND_216[31:0];
  _RAND_217 = {1{`RANDOM}};
  result_nextBestPipe_bits_23_z = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  result_nextPipe_valid_24 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  result_nextPipe_bits_24_x = _RAND_219[31:0];
  _RAND_220 = {1{`RANDOM}};
  result_nextPipe_bits_24_y = _RAND_220[31:0];
  _RAND_221 = {1{`RANDOM}};
  result_nextPipe_bits_24_z = _RAND_221[31:0];
  _RAND_222 = {1{`RANDOM}};
  result_nextPipe_bits_24_sigma = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  result_nextBestPipe_valid_24 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  result_nextBestPipe_bits_24_x = _RAND_224[31:0];
  _RAND_225 = {1{`RANDOM}};
  result_nextBestPipe_bits_24_y = _RAND_225[31:0];
  _RAND_226 = {1{`RANDOM}};
  result_nextBestPipe_bits_24_z = _RAND_226[31:0];
  _RAND_227 = {1{`RANDOM}};
  result_nextPipe_valid_25 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  result_nextPipe_bits_25_x = _RAND_228[31:0];
  _RAND_229 = {1{`RANDOM}};
  result_nextPipe_bits_25_y = _RAND_229[31:0];
  _RAND_230 = {1{`RANDOM}};
  result_nextPipe_bits_25_z = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  result_nextPipe_bits_25_sigma = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  result_nextBestPipe_valid_25 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  result_nextBestPipe_bits_25_x = _RAND_233[31:0];
  _RAND_234 = {1{`RANDOM}};
  result_nextBestPipe_bits_25_y = _RAND_234[31:0];
  _RAND_235 = {1{`RANDOM}};
  result_nextBestPipe_bits_25_z = _RAND_235[31:0];
  _RAND_236 = {1{`RANDOM}};
  result_nextPipe_valid_26 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  result_nextPipe_bits_26_x = _RAND_237[31:0];
  _RAND_238 = {1{`RANDOM}};
  result_nextPipe_bits_26_y = _RAND_238[31:0];
  _RAND_239 = {1{`RANDOM}};
  result_nextPipe_bits_26_z = _RAND_239[31:0];
  _RAND_240 = {1{`RANDOM}};
  result_nextPipe_bits_26_sigma = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  result_nextBestPipe_valid_26 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  result_nextBestPipe_bits_26_x = _RAND_242[31:0];
  _RAND_243 = {1{`RANDOM}};
  result_nextBestPipe_bits_26_y = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  result_nextBestPipe_bits_26_z = _RAND_244[31:0];
  _RAND_245 = {1{`RANDOM}};
  result_nextPipe_valid_27 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  result_nextPipe_bits_27_x = _RAND_246[31:0];
  _RAND_247 = {1{`RANDOM}};
  result_nextPipe_bits_27_y = _RAND_247[31:0];
  _RAND_248 = {1{`RANDOM}};
  result_nextPipe_bits_27_z = _RAND_248[31:0];
  _RAND_249 = {1{`RANDOM}};
  result_nextPipe_bits_27_sigma = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  result_nextBestPipe_valid_27 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  result_nextBestPipe_bits_27_x = _RAND_251[31:0];
  _RAND_252 = {1{`RANDOM}};
  result_nextBestPipe_bits_27_y = _RAND_252[31:0];
  _RAND_253 = {1{`RANDOM}};
  result_nextBestPipe_bits_27_z = _RAND_253[31:0];
  _RAND_254 = {1{`RANDOM}};
  result_nextPipe_valid_28 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  result_nextPipe_bits_28_x = _RAND_255[31:0];
  _RAND_256 = {1{`RANDOM}};
  result_nextPipe_bits_28_y = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  result_nextPipe_bits_28_z = _RAND_257[31:0];
  _RAND_258 = {1{`RANDOM}};
  result_nextPipe_bits_28_sigma = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  result_nextBestPipe_valid_28 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  result_nextBestPipe_bits_28_x = _RAND_260[31:0];
  _RAND_261 = {1{`RANDOM}};
  result_nextBestPipe_bits_28_y = _RAND_261[31:0];
  _RAND_262 = {1{`RANDOM}};
  result_nextBestPipe_bits_28_z = _RAND_262[31:0];
  _RAND_263 = {1{`RANDOM}};
  result_nextPipe_valid_29 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  result_nextPipe_bits_29_x = _RAND_264[31:0];
  _RAND_265 = {1{`RANDOM}};
  result_nextPipe_bits_29_y = _RAND_265[31:0];
  _RAND_266 = {1{`RANDOM}};
  result_nextPipe_bits_29_z = _RAND_266[31:0];
  _RAND_267 = {1{`RANDOM}};
  result_nextPipe_bits_29_sigma = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  result_nextBestPipe_valid_29 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  result_nextBestPipe_bits_29_x = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  result_nextBestPipe_bits_29_y = _RAND_270[31:0];
  _RAND_271 = {1{`RANDOM}};
  result_nextBestPipe_bits_29_z = _RAND_271[31:0];
  _RAND_272 = {1{`RANDOM}};
  result_nextPipe_bits_30_x = _RAND_272[31:0];
  _RAND_273 = {1{`RANDOM}};
  result_nextPipe_bits_30_y = _RAND_273[31:0];
  _RAND_274 = {1{`RANDOM}};
  result_nextPipe_bits_30_z = _RAND_274[31:0];
  _RAND_275 = {1{`RANDOM}};
  result_nextPipe_bits_30_sigma = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  result_nextBestPipe_valid_30 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  result_nextBestPipe_bits_30_x = _RAND_277[31:0];
  _RAND_278 = {1{`RANDOM}};
  result_nextBestPipe_bits_30_y = _RAND_278[31:0];
  _RAND_279 = {1{`RANDOM}};
  result_nextBestPipe_bits_30_z = _RAND_279[31:0];
  _RAND_280 = {1{`RANDOM}};
  resultPipe_valid = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  resultPipe_bits_x = _RAND_281[31:0];
  _RAND_282 = {1{`RANDOM}};
  resultPipe_bits_y = _RAND_282[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SquareRootLog(
  input         clock,
  input         reset,
  input         io_uniform_valid,
  input  [31:0] io_uniform_bits,
  output        io_result_valid,
  output [51:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
`endif // RANDOMIZE_REG_INIT
  reg [51:0] arg; // @[SquareRootLog.scala 49:16]
  wire [34:0] _GEN_10 = {$signed(io_uniform_bits), 3'h0}; // @[SquareRootLog.scala 49:16 50:{26,32}]
  reg  result_v; // @[Valid.scala 127:22]
  wire [103:0] _result_mul_T = 52'sh441b23a29c7 * $signed(arg); // @[SquareRootLog.scala 42:24]
  wire [71:0] _GEN_11 = _result_mul_T[103:32]; // @[SquareRootLog.scala 41:21 42:11]
  wire [51:0] result_mul = _GEN_11[51:0]; // @[SquareRootLog.scala 41:21 42:11]
  wire [51:0] result_next = $signed(result_mul) - 52'sh129b3b5f1bef; // @[SquareRootLog.scala 44:19]
  reg  result_v_1; // @[Valid.scala 127:22]
  reg [51:0] result_b_1; // @[Reg.scala 16:16]
  reg [51:0] result_REG; // @[SquareRootLog.scala 45:51]
  wire [103:0] _result_mul_T_1 = $signed(result_b_1) * $signed(result_REG); // @[SquareRootLog.scala 42:24]
  wire [71:0] _GEN_13 = _result_mul_T_1[103:32]; // @[SquareRootLog.scala 41:21 42:11]
  wire [51:0] result_mul_1 = _GEN_13[51:0]; // @[SquareRootLog.scala 41:21 42:11]
  wire [51:0] result_next_1 = $signed(result_mul_1) + 52'sh21b2370ed3d8; // @[SquareRootLog.scala 44:19]
  reg  result_v_2; // @[Valid.scala 127:22]
  reg [51:0] result_b_2; // @[Reg.scala 16:16]
  reg [51:0] result_REG_1; // @[SquareRootLog.scala 45:51]
  wire [103:0] _result_mul_T_2 = $signed(result_b_2) * $signed(result_REG_1); // @[SquareRootLog.scala 42:24]
  wire [71:0] _GEN_15 = _result_mul_T_2[103:32]; // @[SquareRootLog.scala 41:21 42:11]
  wire [51:0] result_mul_2 = _GEN_15[51:0]; // @[SquareRootLog.scala 41:21 42:11]
  wire [51:0] result_next_2 = $signed(result_mul_2) - 52'sh20b8922291fb; // @[SquareRootLog.scala 44:19]
  reg  result_v_3; // @[Valid.scala 127:22]
  reg [51:0] result_b_3; // @[Reg.scala 16:16]
  reg [51:0] result_REG_2; // @[SquareRootLog.scala 45:51]
  wire [103:0] _result_mul_T_3 = $signed(result_b_3) * $signed(result_REG_2); // @[SquareRootLog.scala 42:24]
  wire [71:0] _GEN_17 = _result_mul_T_3[103:32]; // @[SquareRootLog.scala 41:21 42:11]
  wire [51:0] result_mul_3 = _GEN_17[51:0]; // @[SquareRootLog.scala 41:21 42:11]
  wire [51:0] result_next_3 = $signed(result_mul_3) + 52'sh126c2a5e353f; // @[SquareRootLog.scala 44:19]
  reg  result_v_4; // @[Valid.scala 127:22]
  reg [51:0] result_b_4; // @[Reg.scala 16:16]
  reg [51:0] result_REG_3; // @[SquareRootLog.scala 45:51]
  wire [103:0] _result_mul_T_4 = $signed(result_b_4) * $signed(result_REG_3); // @[SquareRootLog.scala 42:24]
  wire [71:0] _GEN_19 = _result_mul_T_4[103:32]; // @[SquareRootLog.scala 41:21 42:11]
  wire [51:0] result_mul_4 = _GEN_19[51:0]; // @[SquareRootLog.scala 41:21 42:11]
  wire [51:0] result_next_4 = $signed(result_mul_4) - 52'sh614d1ba5e35; // @[SquareRootLog.scala 44:19]
  reg  result_v_5; // @[Valid.scala 127:22]
  reg [51:0] result_b_5; // @[Reg.scala 16:16]
  reg [51:0] result_REG_4; // @[SquareRootLog.scala 45:51]
  wire [103:0] _result_mul_T_5 = $signed(result_b_5) * $signed(result_REG_4); // @[SquareRootLog.scala 42:24]
  wire [71:0] _GEN_21 = _result_mul_T_5[103:32]; // @[SquareRootLog.scala 41:21 42:11]
  wire [51:0] result_mul_5 = _GEN_21[51:0]; // @[SquareRootLog.scala 41:21 42:11]
  wire [51:0] result_next_5 = $signed(result_mul_5) + 52'sh12459f59cd0; // @[SquareRootLog.scala 44:19]
  reg  result_v_6; // @[Valid.scala 127:22]
  reg [51:0] result_b_6; // @[Reg.scala 16:16]
  reg [51:0] result_REG_5; // @[SquareRootLog.scala 45:51]
  wire [103:0] _result_mul_T_6 = $signed(result_b_6) * $signed(result_REG_5); // @[SquareRootLog.scala 42:24]
  wire [71:0] _GEN_23 = _result_mul_T_6[103:32]; // @[SquareRootLog.scala 41:21 42:11]
  wire [51:0] result_mul_6 = _GEN_23[51:0]; // @[SquareRootLog.scala 41:21 42:11]
  wire [51:0] result_next_6 = $signed(result_mul_6) - 52'sh1f22f5d85f; // @[SquareRootLog.scala 44:19]
  reg  result_v_7; // @[Valid.scala 127:22]
  reg [51:0] result_b_7; // @[Reg.scala 16:16]
  reg [51:0] result_REG_6; // @[SquareRootLog.scala 45:51]
  wire [103:0] _result_mul_T_7 = $signed(result_b_7) * $signed(result_REG_6); // @[SquareRootLog.scala 42:24]
  wire [71:0] _GEN_25 = _result_mul_T_7[103:32]; // @[SquareRootLog.scala 41:21 42:11]
  wire [51:0] result_mul_7 = _GEN_25[51:0]; // @[SquareRootLog.scala 41:21 42:11]
  wire [51:0] result_next_7 = $signed(result_mul_7) + 52'sh37316176f; // @[SquareRootLog.scala 44:19]
  reg  resultPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] resultPipe_bits; // @[Reg.scala 16:16]
  assign io_result_valid = resultPipe_valid; // @[Valid.scala 122:21 123:17]
  assign io_result_bits = resultPipe_bits; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    if (io_uniform_valid) begin // @[SquareRootLog.scala 50:26]
      arg <= {{17{_GEN_10[34]}},_GEN_10}; // @[SquareRootLog.scala 50:32]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_v <= io_uniform_valid; // @[Valid.scala 127:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      result_v_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_v_1 <= result_v; // @[Valid.scala 127:22]
    end
    if (result_v) begin // @[Reg.scala 17:18]
      result_b_1 <= result_next; // @[Reg.scala 17:22]
    end
    result_REG <= arg; // @[SquareRootLog.scala 45:51]
    if (reset) begin // @[Valid.scala 127:22]
      result_v_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_v_2 <= result_v_1; // @[Valid.scala 127:22]
    end
    if (result_v_1) begin // @[Reg.scala 17:18]
      result_b_2 <= result_next_1; // @[Reg.scala 17:22]
    end
    result_REG_1 <= result_REG; // @[SquareRootLog.scala 45:51]
    if (reset) begin // @[Valid.scala 127:22]
      result_v_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_v_3 <= result_v_2; // @[Valid.scala 127:22]
    end
    if (result_v_2) begin // @[Reg.scala 17:18]
      result_b_3 <= result_next_2; // @[Reg.scala 17:22]
    end
    result_REG_2 <= result_REG_1; // @[SquareRootLog.scala 45:51]
    if (reset) begin // @[Valid.scala 127:22]
      result_v_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_v_4 <= result_v_3; // @[Valid.scala 127:22]
    end
    if (result_v_3) begin // @[Reg.scala 17:18]
      result_b_4 <= result_next_3; // @[Reg.scala 17:22]
    end
    result_REG_3 <= result_REG_2; // @[SquareRootLog.scala 45:51]
    if (reset) begin // @[Valid.scala 127:22]
      result_v_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_v_5 <= result_v_4; // @[Valid.scala 127:22]
    end
    if (result_v_4) begin // @[Reg.scala 17:18]
      result_b_5 <= result_next_4; // @[Reg.scala 17:22]
    end
    result_REG_4 <= result_REG_3; // @[SquareRootLog.scala 45:51]
    if (reset) begin // @[Valid.scala 127:22]
      result_v_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_v_6 <= result_v_5; // @[Valid.scala 127:22]
    end
    if (result_v_5) begin // @[Reg.scala 17:18]
      result_b_6 <= result_next_5; // @[Reg.scala 17:22]
    end
    result_REG_5 <= result_REG_4; // @[SquareRootLog.scala 45:51]
    if (reset) begin // @[Valid.scala 127:22]
      result_v_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      result_v_7 <= result_v_6; // @[Valid.scala 127:22]
    end
    if (result_v_6) begin // @[Reg.scala 17:18]
      result_b_7 <= result_next_6; // @[Reg.scala 17:22]
    end
    result_REG_6 <= result_REG_5; // @[SquareRootLog.scala 45:51]
    if (reset) begin // @[Valid.scala 127:22]
      resultPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      resultPipe_valid <= result_v_7; // @[Valid.scala 127:22]
    end
    if (result_v_7) begin // @[Reg.scala 17:18]
      resultPipe_bits <= result_next_7; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  arg = _RAND_0[51:0];
  _RAND_1 = {1{`RANDOM}};
  result_v = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  result_v_1 = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  result_b_1 = _RAND_3[51:0];
  _RAND_4 = {2{`RANDOM}};
  result_REG = _RAND_4[51:0];
  _RAND_5 = {1{`RANDOM}};
  result_v_2 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  result_b_2 = _RAND_6[51:0];
  _RAND_7 = {2{`RANDOM}};
  result_REG_1 = _RAND_7[51:0];
  _RAND_8 = {1{`RANDOM}};
  result_v_3 = _RAND_8[0:0];
  _RAND_9 = {2{`RANDOM}};
  result_b_3 = _RAND_9[51:0];
  _RAND_10 = {2{`RANDOM}};
  result_REG_2 = _RAND_10[51:0];
  _RAND_11 = {1{`RANDOM}};
  result_v_4 = _RAND_11[0:0];
  _RAND_12 = {2{`RANDOM}};
  result_b_4 = _RAND_12[51:0];
  _RAND_13 = {2{`RANDOM}};
  result_REG_3 = _RAND_13[51:0];
  _RAND_14 = {1{`RANDOM}};
  result_v_5 = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  result_b_5 = _RAND_15[51:0];
  _RAND_16 = {2{`RANDOM}};
  result_REG_4 = _RAND_16[51:0];
  _RAND_17 = {1{`RANDOM}};
  result_v_6 = _RAND_17[0:0];
  _RAND_18 = {2{`RANDOM}};
  result_b_6 = _RAND_18[51:0];
  _RAND_19 = {2{`RANDOM}};
  result_REG_5 = _RAND_19[51:0];
  _RAND_20 = {1{`RANDOM}};
  result_v_7 = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  result_b_7 = _RAND_21[51:0];
  _RAND_22 = {2{`RANDOM}};
  result_REG_6 = _RAND_22[51:0];
  _RAND_23 = {1{`RANDOM}};
  resultPipe_valid = _RAND_23[0:0];
  _RAND_24 = {2{`RANDOM}};
  resultPipe_bits = _RAND_24[51:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoxMuller(
  input         clock,
  input         reset,
  output        io_g1_valid,
  output [51:0] io_g1_bits,
  output        io_g2_valid,
  output [51:0] io_g2_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [95:0] _RAND_77;
`endif // RANDOMIZE_REG_INIT
  wire  rng1_clock; // @[BoxMuller.scala 51:20]
  wire  rng1_reset; // @[BoxMuller.scala 51:20]
  wire  rng1_io_rand_valid; // @[BoxMuller.scala 51:20]
  wire [31:0] rng1_io_rand_bits; // @[BoxMuller.scala 51:20]
  wire  rng2_clock; // @[BoxMuller.scala 52:20]
  wire  rng2_reset; // @[BoxMuller.scala 52:20]
  wire  rng2_io_rand_valid; // @[BoxMuller.scala 52:20]
  wire [31:0] rng2_io_rand_bits; // @[BoxMuller.scala 52:20]
  wire  trigonometric_clock; // @[BoxMuller.scala 55:29]
  wire  trigonometric_reset; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_theta_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_theta_bits; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_result_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_sine; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_cosine; // @[BoxMuller.scala 55:29]
  wire  sqrt_log_clock; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_reset; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_uniform_valid; // @[BoxMuller.scala 84:24]
  wire [31:0] sqrt_log_io_uniform_bits; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_result_valid; // @[BoxMuller.scala 84:24]
  wire [51:0] sqrt_log_io_result_bits; // @[BoxMuller.scala 84:24]
  wire [30:0] _theta_T_3 = {2'h0,rng1_io_rand_bits[28:0]}; // @[BoxMuller.scala 62:18]
  wire [62:0] _theta_T_4 = $signed(_theta_T_3) * 32'sh6487ed51; // @[BoxMuller.scala 62:26]
  reg  quadrantPipe_valid; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_1; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_1; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_2; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_2; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_3; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_3; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_4; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_4; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_5; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_5; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_6; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_6; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_7; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_7; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_8; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_8; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_9; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_9; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_10; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_10; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_11; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_11; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_12; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_12; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_13; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_13; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_14; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_14; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_15; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_15; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_16; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_16; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_17; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_17; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_18; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_18; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_19; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_19; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_20; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_20; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_21; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_21; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_22; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_22; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_23; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_23; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_24; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_24; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_25; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_25; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_26; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_26; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_27; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_27; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_28; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_28; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_29; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_29; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_30; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_30; // @[Reg.scala 16:16]
  reg [1:0] quadrantPipe_bits_31; // @[Reg.scala 16:16]
  reg  trigonometric_io_theta_v; // @[Valid.scala 127:22]
  reg [31:0] trigonometric_io_theta_b; // @[Reg.scala 16:16]
  wire [33:0] _GEN_40 = _theta_T_4[62:29]; // @[BoxMuller.scala 59:19 61:9]
  wire [31:0] theta = _GEN_40[31:0]; // @[BoxMuller.scala 59:19 61:9]
  wire  _cosine_T = quadrantPipe_bits_31 == 2'h0; // @[BoxMuller.scala 70:21]
  wire  _cosine_T_2 = quadrantPipe_bits_31 == 2'h0 | quadrantPipe_bits_31 == 2'h3; // @[BoxMuller.scala 70:29]
  wire [31:0] _cosine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_cosine); // @[BoxMuller.scala 72:7]
  reg  cosinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] cosinePipe_bits; // @[Reg.scala 16:16]
  wire  _sine_T_2 = _cosine_T | quadrantPipe_bits_31 == 2'h2; // @[BoxMuller.scala 78:29]
  wire [31:0] _sine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_sine); // @[BoxMuller.scala 80:7]
  reg  sinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] sinePipe_bits; // @[Reg.scala 16:16]
  reg  signPipe_bits; // @[Reg.scala 16:16]
  wire [28:0] _sqrt_log_io_uniform_T_1 = rng2_io_rand_bits[28:0]; // @[BoxMuller.scala 87:89]
  reg  sqrt_log_io_uniform_v; // @[Valid.scala 127:22]
  reg [28:0] sqrt_log_io_uniform_b; // @[Reg.scala 16:16]
  wire [51:0] _sign_adjusted_T_3 = 52'sh0 - $signed(sqrt_log_io_result_bits); // @[BoxMuller.scala 93:7]
  reg  sign_adjustedPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] sign_adjustedPipe_bits; // @[Reg.scala 16:16]
  wire  _io_g1_T = sign_adjustedPipe_valid & cosinePipe_valid; // @[BoxMuller.scala 99:25]
  wire [83:0] _io_g1_T_1 = $signed(cosinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 100:17]
  reg  io_g1_v; // @[Valid.scala 127:22]
  reg [83:0] io_g1_b; // @[Reg.scala 16:16]
  wire  _io_g2_T = sign_adjustedPipe_valid & sinePipe_valid; // @[BoxMuller.scala 103:25]
  wire [83:0] _io_g2_T_1 = $signed(sinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 104:15]
  reg  io_g2_v; // @[Valid.scala 127:22]
  reg [83:0] io_g2_b; // @[Reg.scala 16:16]
  wire [53:0] _GEN_42 = io_g1_b[83:30]; // @[BoxMuller.scala 98:9]
  wire [53:0] _GEN_44 = io_g2_b[83:30]; // @[BoxMuller.scala 102:9]
  wire [32:0] _GEN_46 = {$signed(trigonometric_io_theta_b), 1'h0}; // @[BoxMuller.scala 65:26]
  TauswortheUniform rng1 ( // @[BoxMuller.scala 51:20]
    .clock(rng1_clock),
    .reset(rng1_reset),
    .io_rand_valid(rng1_io_rand_valid),
    .io_rand_bits(rng1_io_rand_bits)
  );
  TauswortheUniform_1 rng2 ( // @[BoxMuller.scala 52:20]
    .clock(rng2_clock),
    .reset(rng2_reset),
    .io_rand_valid(rng2_io_rand_valid),
    .io_rand_bits(rng2_io_rand_bits)
  );
  Trigonometric trigonometric ( // @[BoxMuller.scala 55:29]
    .clock(trigonometric_clock),
    .reset(trigonometric_reset),
    .io_theta_valid(trigonometric_io_theta_valid),
    .io_theta_bits(trigonometric_io_theta_bits),
    .io_result_valid(trigonometric_io_result_valid),
    .io_result_bits_sine(trigonometric_io_result_bits_sine),
    .io_result_bits_cosine(trigonometric_io_result_bits_cosine)
  );
  SquareRootLog sqrt_log ( // @[BoxMuller.scala 84:24]
    .clock(sqrt_log_clock),
    .reset(sqrt_log_reset),
    .io_uniform_valid(sqrt_log_io_uniform_valid),
    .io_uniform_bits(sqrt_log_io_uniform_bits),
    .io_result_valid(sqrt_log_io_result_valid),
    .io_result_bits(sqrt_log_io_result_bits)
  );
  assign io_g1_valid = io_g1_v; // @[Valid.scala 122:21 123:17]
  assign io_g1_bits = _GEN_42[51:0]; // @[BoxMuller.scala 98:9]
  assign io_g2_valid = io_g2_v; // @[Valid.scala 122:21 123:17]
  assign io_g2_bits = _GEN_44[51:0]; // @[BoxMuller.scala 102:9]
  assign rng1_clock = clock;
  assign rng1_reset = reset;
  assign rng2_clock = clock;
  assign rng2_reset = reset;
  assign trigonometric_clock = clock;
  assign trigonometric_reset = reset;
  assign trigonometric_io_theta_valid = trigonometric_io_theta_v; // @[Valid.scala 122:21 123:17]
  assign trigonometric_io_theta_bits = _GEN_46[31:0]; // @[BoxMuller.scala 65:26]
  assign sqrt_log_clock = clock;
  assign sqrt_log_reset = reset;
  assign sqrt_log_io_uniform_valid = sqrt_log_io_uniform_v; // @[Valid.scala 122:21 123:17]
  assign sqrt_log_io_uniform_bits = {{3{sqrt_log_io_uniform_b[28]}},sqrt_log_io_uniform_b}; // @[BoxMuller.scala 87:23]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits <= rng1_io_rand_bits[31:30]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_1 <= quadrantPipe_valid; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_1 <= quadrantPipe_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_2 <= quadrantPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_1) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_2 <= quadrantPipe_bits_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_3 <= quadrantPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_2) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_3 <= quadrantPipe_bits_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_4 <= quadrantPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_3) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_4 <= quadrantPipe_bits_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_5 <= quadrantPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_4) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_5 <= quadrantPipe_bits_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_6 <= quadrantPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_5) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_6 <= quadrantPipe_bits_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_7 <= quadrantPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_6) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_7 <= quadrantPipe_bits_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_8 <= quadrantPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_7) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_8 <= quadrantPipe_bits_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_9 <= quadrantPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_8) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_9 <= quadrantPipe_bits_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_10 <= quadrantPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_9) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_10 <= quadrantPipe_bits_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_11 <= quadrantPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_10) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_11 <= quadrantPipe_bits_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_12 <= quadrantPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_11) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_12 <= quadrantPipe_bits_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_13 <= quadrantPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_12) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_13 <= quadrantPipe_bits_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_14 <= quadrantPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_13) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_14 <= quadrantPipe_bits_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_15 <= quadrantPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_14) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_15 <= quadrantPipe_bits_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_16 <= quadrantPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_15) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_16 <= quadrantPipe_bits_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_17 <= quadrantPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_16) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_17 <= quadrantPipe_bits_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_18 <= quadrantPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_17) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_18 <= quadrantPipe_bits_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_19 <= quadrantPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_18) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_19 <= quadrantPipe_bits_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_20 <= quadrantPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_19) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_20 <= quadrantPipe_bits_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_21 <= quadrantPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_20) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_21 <= quadrantPipe_bits_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_22 <= quadrantPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_21) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_22 <= quadrantPipe_bits_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_23 <= quadrantPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_22) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_23 <= quadrantPipe_bits_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_24 <= quadrantPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_23) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_24 <= quadrantPipe_bits_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_25 <= quadrantPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_24) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_25 <= quadrantPipe_bits_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_26 <= quadrantPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_25) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_26 <= quadrantPipe_bits_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_27 <= quadrantPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_26) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_27 <= quadrantPipe_bits_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_28 <= quadrantPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_27) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_28 <= quadrantPipe_bits_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_29 <= quadrantPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_28) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_29 <= quadrantPipe_bits_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_30 <= quadrantPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_29) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_30 <= quadrantPipe_bits_29; // @[Reg.scala 17:22]
    end
    if (quadrantPipe_valid_30) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_31 <= quadrantPipe_bits_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      trigonometric_io_theta_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      trigonometric_io_theta_v <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      trigonometric_io_theta_b <= theta; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      cosinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      cosinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_cosine_T_2) begin // @[BoxMuller.scala 69:8]
        cosinePipe_bits <= trigonometric_io_result_bits_cosine;
      end else begin
        cosinePipe_bits <= _cosine_T_5;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      sinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_sine_T_2) begin // @[BoxMuller.scala 77:8]
        sinePipe_bits <= trigonometric_io_result_bits_sine;
      end else begin
        sinePipe_bits <= _sine_T_5;
      end
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      signPipe_bits <= rng2_io_rand_bits[31]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sqrt_log_io_uniform_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sqrt_log_io_uniform_v <= rng2_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      sqrt_log_io_uniform_b <= _sqrt_log_io_uniform_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sign_adjustedPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sign_adjustedPipe_valid <= sqrt_log_io_result_valid; // @[Valid.scala 127:22]
    end
    if (sqrt_log_io_result_valid) begin // @[Reg.scala 17:18]
      if (signPipe_bits) begin // @[BoxMuller.scala 91:8]
        sign_adjustedPipe_bits <= _sign_adjusted_T_3;
      end else begin
        sign_adjustedPipe_bits <= sqrt_log_io_result_bits;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g1_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g1_v <= _io_g1_T; // @[Valid.scala 127:22]
    end
    if (_io_g1_T) begin // @[Reg.scala 17:18]
      io_g1_b <= _io_g1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g2_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g2_v <= _io_g2_T; // @[Valid.scala 127:22]
    end
    if (_io_g2_T) begin // @[Reg.scala 17:18]
      io_g2_b <= _io_g2_T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quadrantPipe_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  quadrantPipe_bits = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  quadrantPipe_valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  quadrantPipe_bits_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  quadrantPipe_valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  quadrantPipe_bits_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  quadrantPipe_valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quadrantPipe_bits_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  quadrantPipe_valid_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  quadrantPipe_bits_4 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  quadrantPipe_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  quadrantPipe_bits_5 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  quadrantPipe_valid_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  quadrantPipe_bits_6 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  quadrantPipe_valid_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  quadrantPipe_bits_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  quadrantPipe_valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  quadrantPipe_bits_8 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  quadrantPipe_valid_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  quadrantPipe_bits_9 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  quadrantPipe_valid_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  quadrantPipe_bits_10 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  quadrantPipe_valid_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  quadrantPipe_bits_11 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  quadrantPipe_valid_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  quadrantPipe_bits_12 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  quadrantPipe_valid_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  quadrantPipe_bits_13 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  quadrantPipe_valid_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  quadrantPipe_bits_14 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  quadrantPipe_valid_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  quadrantPipe_bits_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  quadrantPipe_valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  quadrantPipe_bits_16 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  quadrantPipe_valid_17 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  quadrantPipe_bits_17 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  quadrantPipe_valid_18 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  quadrantPipe_bits_18 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  quadrantPipe_valid_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  quadrantPipe_bits_19 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  quadrantPipe_valid_20 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  quadrantPipe_bits_20 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  quadrantPipe_valid_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  quadrantPipe_bits_21 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  quadrantPipe_valid_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  quadrantPipe_bits_22 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  quadrantPipe_valid_23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  quadrantPipe_bits_23 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  quadrantPipe_valid_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  quadrantPipe_bits_24 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  quadrantPipe_valid_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  quadrantPipe_bits_25 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  quadrantPipe_valid_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  quadrantPipe_bits_26 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  quadrantPipe_valid_27 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  quadrantPipe_bits_27 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  quadrantPipe_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  quadrantPipe_bits_28 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  quadrantPipe_valid_29 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  quadrantPipe_bits_29 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  quadrantPipe_valid_30 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  quadrantPipe_bits_30 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  quadrantPipe_bits_31 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  trigonometric_io_theta_v = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  trigonometric_io_theta_b = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cosinePipe_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cosinePipe_bits = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sinePipe_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sinePipe_bits = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  signPipe_bits = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sqrt_log_io_uniform_v = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sqrt_log_io_uniform_b = _RAND_71[28:0];
  _RAND_72 = {1{`RANDOM}};
  sign_adjustedPipe_valid = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  sign_adjustedPipe_bits = _RAND_73[51:0];
  _RAND_74 = {1{`RANDOM}};
  io_g1_v = _RAND_74[0:0];
  _RAND_75 = {3{`RANDOM}};
  io_g1_b = _RAND_75[83:0];
  _RAND_76 = {1{`RANDOM}};
  io_g2_v = _RAND_76[0:0];
  _RAND_77 = {3{`RANDOM}};
  io_g2_b = _RAND_77[83:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MonteCarlo(
  input         clock,
  input         reset,
  output        io_request_0_ready,
  input         io_request_0_valid,
  input  [31:0] io_request_0_bits_time_steps,
  input  [31:0] io_request_0_bits_start_value,
  input  [31:0] io_request_0_bits_coefficient1,
  input  [31:0] io_request_0_bits_coefficient2,
  output        io_request_1_ready,
  input         io_request_1_valid,
  input  [31:0] io_request_1_bits_time_steps,
  input  [31:0] io_request_1_bits_start_value,
  input  [31:0] io_request_1_bits_coefficient1,
  input  [31:0] io_request_1_bits_coefficient2,
  input         io_response_0_ready,
  output        io_response_0_valid,
  output [31:0] io_response_0_bits,
  input         io_response_1_ready,
  output        io_response_1_valid,
  output [31:0] io_response_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rng_clock; // @[MonteCarlo.scala 42:19]
  wire  rng_reset; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g1_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g1_bits; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g2_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g2_bits; // @[MonteCarlo.scala 42:19]
  wire  initialized = rng_io_g1_valid & rng_io_g2_valid; // @[MonteCarlo.scala 47:37]
  reg [2:0] state; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_2 = $signed(io_request_0_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_3 = io_request_0_ready & io_request_0_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1; // @[Reg.scala 16:16]
  reg [31:0] c2; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_1 = io_request_0_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step; // @[Reg.scala 16:16]
  reg [31:0] price; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T = $signed(price) * $signed(c1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T = $signed(rng_io_g1_bits) * $signed(c2); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T = $signed(price) * $signed(partial_res2); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_2 = $signed(partial_res3) + $signed(partial_res1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_3 = counter == last_step ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_4 = counter == last_step ? counter : _counter_T_1; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_7 = io_response_0_ready & io_response_0_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_5 = _T_7 ? 3'h1 : state; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_6 = 3'h5 == state ? _GEN_5 : state; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_7 = 3'h4 == state ? $signed(_price_T_2) : $signed(price); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_3 : _GEN_6; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_9 = 3'h4 == state ? _GEN_4 : counter; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_64 = {$signed(partial_res3), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_10 = 3'h3 == state ? $signed(_partial_res3_T) : $signed({{12{_GEN_64[51]}},_GEN_64}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_11 = 3'h3 == state ? 3'h4 : _GEN_8; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_65 = {$signed(partial_res1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_14 = 3'h2 == state ? $signed(_partial_res1_T) : $signed({{12{_GEN_65[51]}},_GEN_65}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_66 = {$signed(partial_res2), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_15 = 3'h2 == state ? $signed(_partial_res2_T) : $signed({{20{_GEN_66[63]}},_GEN_66}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_17 = 3'h2 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_10); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_23 = 3'h1 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_14); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_24 = 3'h1 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_15); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_25 = 3'h1 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_17); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_29 = 3'h0 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_23); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_30 = 3'h0 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_24); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_31 = 3'h0 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_25); // @[MonteCarlo.scala 66:19 60:27]
  reg [2:0] state_1; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_6 = $signed(io_request_1_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_7 = io_request_1_ready & io_request_1_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1_1; // @[Reg.scala 16:16]
  reg [31:0] c2_1; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_4 = io_request_1_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step_1; // @[Reg.scala 16:16]
  reg [31:0] price_1; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1_1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2_1; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3_1; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter_1; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T_1 = $signed(price_1) * $signed(c1_1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T_1 = $signed(rng_io_g2_bits) * $signed(c2_1); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T_1 = $signed(price_1) * $signed(partial_res2_1); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_5 = $signed(partial_res3_1) + $signed(partial_res1_1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_35 = counter_1 == last_step_1 ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_36 = counter_1 == last_step_1 ? counter_1 : _counter_T_3; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_15 = io_response_1_ready & io_response_1_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_37 = _T_15 ? 3'h1 : state_1; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_38 = 3'h5 == state_1 ? _GEN_37 : state_1; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_39 = 3'h4 == state_1 ? $signed(_price_T_5) : $signed(price_1); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_40 = 3'h4 == state_1 ? _GEN_35 : _GEN_38; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_41 = 3'h4 == state_1 ? _GEN_36 : counter_1; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_74 = {$signed(partial_res3_1), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_42 = 3'h3 == state_1 ? $signed(_partial_res3_T_1) : $signed({{12{_GEN_74[51]}},_GEN_74}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_43 = 3'h3 == state_1 ? 3'h4 : _GEN_40; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_75 = {$signed(partial_res1_1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_46 = 3'h2 == state_1 ? $signed(_partial_res1_T_1) : $signed({{12{_GEN_75[51]}},_GEN_75}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_76 = {$signed(partial_res2_1), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_47 = 3'h2 == state_1 ? $signed(_partial_res2_T_1) : $signed({{20{_GEN_76[63]}},_GEN_76}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_49 = 3'h2 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_42); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_55 = 3'h1 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_46); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_56 = 3'h1 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_47); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_57 = 3'h1 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_49); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_61 = 3'h0 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_55); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_62 = 3'h0 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_56); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_63 = 3'h0 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_57); // @[MonteCarlo.scala 66:19 60:27]
  wire [43:0] _GEN_84 = _GEN_29[63:20];
  wire [51:0] _GEN_86 = _GEN_30[83:32];
  wire [43:0] _GEN_88 = _GEN_31[63:20];
  wire [43:0] _GEN_90 = _GEN_61[63:20];
  wire [51:0] _GEN_92 = _GEN_62[83:32];
  wire [43:0] _GEN_94 = _GEN_63[63:20];
  BoxMuller rng ( // @[MonteCarlo.scala 42:19]
    .clock(rng_clock),
    .reset(rng_reset),
    .io_g1_valid(rng_io_g1_valid),
    .io_g1_bits(rng_io_g1_bits),
    .io_g2_valid(rng_io_g2_valid),
    .io_g2_bits(rng_io_g2_bits)
  );
  assign io_request_0_ready = state == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_request_1_ready = state_1 == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_response_0_valid = state == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_0_bits = price; // @[MonteCarlo.scala 65:16]
  assign io_response_1_valid = state_1 == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_1_bits = price_1; // @[MonteCarlo.scala 65:16]
  assign rng_clock = clock;
  assign rng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state <= 3'h1;
      end else begin
        state <= 3'h0;
      end
    end else if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_3) begin // @[MonteCarlo.scala 71:23]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[MonteCarlo.scala 66:19]
      state <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state <= _GEN_11;
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c1 <= _c1_T_2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c2 <= io_request_0_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      last_step <= _last_step_T_1; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        price <= io_request_0_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          price <= _GEN_7;
        end
      end
    end
    partial_res1 <= _GEN_84[31:0];
    partial_res2 <= _GEN_86[31:0];
    partial_res3 <= _GEN_88[31:0];
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        counter <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          counter <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state_1 <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state_1 <= 3'h1;
      end else begin
        state_1 <= 3'h0;
      end
    end else if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_7) begin // @[MonteCarlo.scala 71:23]
        state_1 <= 3'h2;
      end else begin
        state_1 <= 3'h1;
      end
    end else if (3'h2 == state_1) begin // @[MonteCarlo.scala 66:19]
      state_1 <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state_1 <= _GEN_43;
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c1_1 <= _c1_T_6; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c2_1 <= io_request_1_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      last_step_1 <= _last_step_T_4; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        price_1 <= io_request_1_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          price_1 <= _GEN_39;
        end
      end
    end
    partial_res1_1 <= _GEN_90[31:0];
    partial_res2_1 <= _GEN_92[31:0];
    partial_res3_1 <= _GEN_94[31:0];
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        counter_1 <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          counter_1 <= _GEN_41;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  c1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_step = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  price = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  partial_res1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  partial_res2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  partial_res3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  c1_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_step_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  price_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  partial_res1_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  partial_res2_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  partial_res3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  counter_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_2(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h233a5c2d : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h77d0940 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h263e2e8f : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_3(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h3204a9db : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h1553734a : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h102d7c12 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoxMuller_1(
  input         clock,
  input         reset,
  output        io_g1_valid,
  output [51:0] io_g1_bits,
  output        io_g2_valid,
  output [51:0] io_g2_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [95:0] _RAND_77;
`endif // RANDOMIZE_REG_INIT
  wire  rng1_clock; // @[BoxMuller.scala 51:20]
  wire  rng1_reset; // @[BoxMuller.scala 51:20]
  wire  rng1_io_rand_valid; // @[BoxMuller.scala 51:20]
  wire [31:0] rng1_io_rand_bits; // @[BoxMuller.scala 51:20]
  wire  rng2_clock; // @[BoxMuller.scala 52:20]
  wire  rng2_reset; // @[BoxMuller.scala 52:20]
  wire  rng2_io_rand_valid; // @[BoxMuller.scala 52:20]
  wire [31:0] rng2_io_rand_bits; // @[BoxMuller.scala 52:20]
  wire  trigonometric_clock; // @[BoxMuller.scala 55:29]
  wire  trigonometric_reset; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_theta_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_theta_bits; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_result_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_sine; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_cosine; // @[BoxMuller.scala 55:29]
  wire  sqrt_log_clock; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_reset; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_uniform_valid; // @[BoxMuller.scala 84:24]
  wire [31:0] sqrt_log_io_uniform_bits; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_result_valid; // @[BoxMuller.scala 84:24]
  wire [51:0] sqrt_log_io_result_bits; // @[BoxMuller.scala 84:24]
  wire [30:0] _theta_T_3 = {2'h0,rng1_io_rand_bits[28:0]}; // @[BoxMuller.scala 62:18]
  wire [62:0] _theta_T_4 = $signed(_theta_T_3) * 32'sh6487ed51; // @[BoxMuller.scala 62:26]
  reg  quadrantPipe_valid; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_1; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_1; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_2; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_2; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_3; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_3; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_4; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_4; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_5; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_5; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_6; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_6; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_7; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_7; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_8; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_8; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_9; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_9; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_10; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_10; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_11; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_11; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_12; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_12; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_13; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_13; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_14; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_14; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_15; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_15; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_16; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_16; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_17; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_17; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_18; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_18; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_19; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_19; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_20; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_20; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_21; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_21; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_22; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_22; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_23; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_23; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_24; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_24; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_25; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_25; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_26; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_26; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_27; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_27; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_28; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_28; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_29; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_29; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_30; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_30; // @[Reg.scala 16:16]
  reg [1:0] quadrantPipe_bits_31; // @[Reg.scala 16:16]
  reg  trigonometric_io_theta_v; // @[Valid.scala 127:22]
  reg [31:0] trigonometric_io_theta_b; // @[Reg.scala 16:16]
  wire [33:0] _GEN_40 = _theta_T_4[62:29]; // @[BoxMuller.scala 59:19 61:9]
  wire [31:0] theta = _GEN_40[31:0]; // @[BoxMuller.scala 59:19 61:9]
  wire  _cosine_T = quadrantPipe_bits_31 == 2'h0; // @[BoxMuller.scala 70:21]
  wire  _cosine_T_2 = quadrantPipe_bits_31 == 2'h0 | quadrantPipe_bits_31 == 2'h3; // @[BoxMuller.scala 70:29]
  wire [31:0] _cosine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_cosine); // @[BoxMuller.scala 72:7]
  reg  cosinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] cosinePipe_bits; // @[Reg.scala 16:16]
  wire  _sine_T_2 = _cosine_T | quadrantPipe_bits_31 == 2'h2; // @[BoxMuller.scala 78:29]
  wire [31:0] _sine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_sine); // @[BoxMuller.scala 80:7]
  reg  sinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] sinePipe_bits; // @[Reg.scala 16:16]
  reg  signPipe_bits; // @[Reg.scala 16:16]
  wire [28:0] _sqrt_log_io_uniform_T_1 = rng2_io_rand_bits[28:0]; // @[BoxMuller.scala 87:89]
  reg  sqrt_log_io_uniform_v; // @[Valid.scala 127:22]
  reg [28:0] sqrt_log_io_uniform_b; // @[Reg.scala 16:16]
  wire [51:0] _sign_adjusted_T_3 = 52'sh0 - $signed(sqrt_log_io_result_bits); // @[BoxMuller.scala 93:7]
  reg  sign_adjustedPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] sign_adjustedPipe_bits; // @[Reg.scala 16:16]
  wire  _io_g1_T = sign_adjustedPipe_valid & cosinePipe_valid; // @[BoxMuller.scala 99:25]
  wire [83:0] _io_g1_T_1 = $signed(cosinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 100:17]
  reg  io_g1_v; // @[Valid.scala 127:22]
  reg [83:0] io_g1_b; // @[Reg.scala 16:16]
  wire  _io_g2_T = sign_adjustedPipe_valid & sinePipe_valid; // @[BoxMuller.scala 103:25]
  wire [83:0] _io_g2_T_1 = $signed(sinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 104:15]
  reg  io_g2_v; // @[Valid.scala 127:22]
  reg [83:0] io_g2_b; // @[Reg.scala 16:16]
  wire [53:0] _GEN_42 = io_g1_b[83:30]; // @[BoxMuller.scala 98:9]
  wire [53:0] _GEN_44 = io_g2_b[83:30]; // @[BoxMuller.scala 102:9]
  wire [32:0] _GEN_46 = {$signed(trigonometric_io_theta_b), 1'h0}; // @[BoxMuller.scala 65:26]
  TauswortheUniform_2 rng1 ( // @[BoxMuller.scala 51:20]
    .clock(rng1_clock),
    .reset(rng1_reset),
    .io_rand_valid(rng1_io_rand_valid),
    .io_rand_bits(rng1_io_rand_bits)
  );
  TauswortheUniform_3 rng2 ( // @[BoxMuller.scala 52:20]
    .clock(rng2_clock),
    .reset(rng2_reset),
    .io_rand_valid(rng2_io_rand_valid),
    .io_rand_bits(rng2_io_rand_bits)
  );
  Trigonometric trigonometric ( // @[BoxMuller.scala 55:29]
    .clock(trigonometric_clock),
    .reset(trigonometric_reset),
    .io_theta_valid(trigonometric_io_theta_valid),
    .io_theta_bits(trigonometric_io_theta_bits),
    .io_result_valid(trigonometric_io_result_valid),
    .io_result_bits_sine(trigonometric_io_result_bits_sine),
    .io_result_bits_cosine(trigonometric_io_result_bits_cosine)
  );
  SquareRootLog sqrt_log ( // @[BoxMuller.scala 84:24]
    .clock(sqrt_log_clock),
    .reset(sqrt_log_reset),
    .io_uniform_valid(sqrt_log_io_uniform_valid),
    .io_uniform_bits(sqrt_log_io_uniform_bits),
    .io_result_valid(sqrt_log_io_result_valid),
    .io_result_bits(sqrt_log_io_result_bits)
  );
  assign io_g1_valid = io_g1_v; // @[Valid.scala 122:21 123:17]
  assign io_g1_bits = _GEN_42[51:0]; // @[BoxMuller.scala 98:9]
  assign io_g2_valid = io_g2_v; // @[Valid.scala 122:21 123:17]
  assign io_g2_bits = _GEN_44[51:0]; // @[BoxMuller.scala 102:9]
  assign rng1_clock = clock;
  assign rng1_reset = reset;
  assign rng2_clock = clock;
  assign rng2_reset = reset;
  assign trigonometric_clock = clock;
  assign trigonometric_reset = reset;
  assign trigonometric_io_theta_valid = trigonometric_io_theta_v; // @[Valid.scala 122:21 123:17]
  assign trigonometric_io_theta_bits = _GEN_46[31:0]; // @[BoxMuller.scala 65:26]
  assign sqrt_log_clock = clock;
  assign sqrt_log_reset = reset;
  assign sqrt_log_io_uniform_valid = sqrt_log_io_uniform_v; // @[Valid.scala 122:21 123:17]
  assign sqrt_log_io_uniform_bits = {{3{sqrt_log_io_uniform_b[28]}},sqrt_log_io_uniform_b}; // @[BoxMuller.scala 87:23]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits <= rng1_io_rand_bits[31:30]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_1 <= quadrantPipe_valid; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_1 <= quadrantPipe_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_2 <= quadrantPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_1) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_2 <= quadrantPipe_bits_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_3 <= quadrantPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_2) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_3 <= quadrantPipe_bits_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_4 <= quadrantPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_3) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_4 <= quadrantPipe_bits_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_5 <= quadrantPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_4) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_5 <= quadrantPipe_bits_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_6 <= quadrantPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_5) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_6 <= quadrantPipe_bits_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_7 <= quadrantPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_6) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_7 <= quadrantPipe_bits_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_8 <= quadrantPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_7) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_8 <= quadrantPipe_bits_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_9 <= quadrantPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_8) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_9 <= quadrantPipe_bits_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_10 <= quadrantPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_9) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_10 <= quadrantPipe_bits_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_11 <= quadrantPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_10) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_11 <= quadrantPipe_bits_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_12 <= quadrantPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_11) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_12 <= quadrantPipe_bits_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_13 <= quadrantPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_12) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_13 <= quadrantPipe_bits_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_14 <= quadrantPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_13) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_14 <= quadrantPipe_bits_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_15 <= quadrantPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_14) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_15 <= quadrantPipe_bits_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_16 <= quadrantPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_15) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_16 <= quadrantPipe_bits_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_17 <= quadrantPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_16) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_17 <= quadrantPipe_bits_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_18 <= quadrantPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_17) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_18 <= quadrantPipe_bits_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_19 <= quadrantPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_18) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_19 <= quadrantPipe_bits_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_20 <= quadrantPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_19) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_20 <= quadrantPipe_bits_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_21 <= quadrantPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_20) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_21 <= quadrantPipe_bits_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_22 <= quadrantPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_21) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_22 <= quadrantPipe_bits_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_23 <= quadrantPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_22) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_23 <= quadrantPipe_bits_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_24 <= quadrantPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_23) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_24 <= quadrantPipe_bits_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_25 <= quadrantPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_24) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_25 <= quadrantPipe_bits_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_26 <= quadrantPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_25) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_26 <= quadrantPipe_bits_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_27 <= quadrantPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_26) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_27 <= quadrantPipe_bits_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_28 <= quadrantPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_27) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_28 <= quadrantPipe_bits_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_29 <= quadrantPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_28) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_29 <= quadrantPipe_bits_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_30 <= quadrantPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_29) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_30 <= quadrantPipe_bits_29; // @[Reg.scala 17:22]
    end
    if (quadrantPipe_valid_30) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_31 <= quadrantPipe_bits_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      trigonometric_io_theta_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      trigonometric_io_theta_v <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      trigonometric_io_theta_b <= theta; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      cosinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      cosinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_cosine_T_2) begin // @[BoxMuller.scala 69:8]
        cosinePipe_bits <= trigonometric_io_result_bits_cosine;
      end else begin
        cosinePipe_bits <= _cosine_T_5;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      sinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_sine_T_2) begin // @[BoxMuller.scala 77:8]
        sinePipe_bits <= trigonometric_io_result_bits_sine;
      end else begin
        sinePipe_bits <= _sine_T_5;
      end
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      signPipe_bits <= rng2_io_rand_bits[31]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sqrt_log_io_uniform_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sqrt_log_io_uniform_v <= rng2_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      sqrt_log_io_uniform_b <= _sqrt_log_io_uniform_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sign_adjustedPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sign_adjustedPipe_valid <= sqrt_log_io_result_valid; // @[Valid.scala 127:22]
    end
    if (sqrt_log_io_result_valid) begin // @[Reg.scala 17:18]
      if (signPipe_bits) begin // @[BoxMuller.scala 91:8]
        sign_adjustedPipe_bits <= _sign_adjusted_T_3;
      end else begin
        sign_adjustedPipe_bits <= sqrt_log_io_result_bits;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g1_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g1_v <= _io_g1_T; // @[Valid.scala 127:22]
    end
    if (_io_g1_T) begin // @[Reg.scala 17:18]
      io_g1_b <= _io_g1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g2_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g2_v <= _io_g2_T; // @[Valid.scala 127:22]
    end
    if (_io_g2_T) begin // @[Reg.scala 17:18]
      io_g2_b <= _io_g2_T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quadrantPipe_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  quadrantPipe_bits = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  quadrantPipe_valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  quadrantPipe_bits_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  quadrantPipe_valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  quadrantPipe_bits_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  quadrantPipe_valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quadrantPipe_bits_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  quadrantPipe_valid_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  quadrantPipe_bits_4 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  quadrantPipe_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  quadrantPipe_bits_5 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  quadrantPipe_valid_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  quadrantPipe_bits_6 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  quadrantPipe_valid_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  quadrantPipe_bits_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  quadrantPipe_valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  quadrantPipe_bits_8 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  quadrantPipe_valid_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  quadrantPipe_bits_9 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  quadrantPipe_valid_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  quadrantPipe_bits_10 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  quadrantPipe_valid_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  quadrantPipe_bits_11 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  quadrantPipe_valid_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  quadrantPipe_bits_12 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  quadrantPipe_valid_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  quadrantPipe_bits_13 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  quadrantPipe_valid_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  quadrantPipe_bits_14 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  quadrantPipe_valid_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  quadrantPipe_bits_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  quadrantPipe_valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  quadrantPipe_bits_16 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  quadrantPipe_valid_17 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  quadrantPipe_bits_17 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  quadrantPipe_valid_18 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  quadrantPipe_bits_18 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  quadrantPipe_valid_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  quadrantPipe_bits_19 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  quadrantPipe_valid_20 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  quadrantPipe_bits_20 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  quadrantPipe_valid_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  quadrantPipe_bits_21 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  quadrantPipe_valid_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  quadrantPipe_bits_22 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  quadrantPipe_valid_23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  quadrantPipe_bits_23 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  quadrantPipe_valid_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  quadrantPipe_bits_24 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  quadrantPipe_valid_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  quadrantPipe_bits_25 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  quadrantPipe_valid_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  quadrantPipe_bits_26 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  quadrantPipe_valid_27 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  quadrantPipe_bits_27 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  quadrantPipe_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  quadrantPipe_bits_28 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  quadrantPipe_valid_29 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  quadrantPipe_bits_29 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  quadrantPipe_valid_30 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  quadrantPipe_bits_30 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  quadrantPipe_bits_31 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  trigonometric_io_theta_v = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  trigonometric_io_theta_b = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cosinePipe_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cosinePipe_bits = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sinePipe_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sinePipe_bits = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  signPipe_bits = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sqrt_log_io_uniform_v = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sqrt_log_io_uniform_b = _RAND_71[28:0];
  _RAND_72 = {1{`RANDOM}};
  sign_adjustedPipe_valid = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  sign_adjustedPipe_bits = _RAND_73[51:0];
  _RAND_74 = {1{`RANDOM}};
  io_g1_v = _RAND_74[0:0];
  _RAND_75 = {3{`RANDOM}};
  io_g1_b = _RAND_75[83:0];
  _RAND_76 = {1{`RANDOM}};
  io_g2_v = _RAND_76[0:0];
  _RAND_77 = {3{`RANDOM}};
  io_g2_b = _RAND_77[83:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MonteCarlo_1(
  input         clock,
  input         reset,
  output        io_request_0_ready,
  input         io_request_0_valid,
  input  [31:0] io_request_0_bits_time_steps,
  input  [31:0] io_request_0_bits_start_value,
  input  [31:0] io_request_0_bits_coefficient1,
  input  [31:0] io_request_0_bits_coefficient2,
  output        io_request_1_ready,
  input         io_request_1_valid,
  input  [31:0] io_request_1_bits_time_steps,
  input  [31:0] io_request_1_bits_start_value,
  input  [31:0] io_request_1_bits_coefficient1,
  input  [31:0] io_request_1_bits_coefficient2,
  input         io_response_0_ready,
  output        io_response_0_valid,
  output [31:0] io_response_0_bits,
  input         io_response_1_ready,
  output        io_response_1_valid,
  output [31:0] io_response_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rng_clock; // @[MonteCarlo.scala 42:19]
  wire  rng_reset; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g1_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g1_bits; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g2_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g2_bits; // @[MonteCarlo.scala 42:19]
  wire  initialized = rng_io_g1_valid & rng_io_g2_valid; // @[MonteCarlo.scala 47:37]
  reg [2:0] state; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_2 = $signed(io_request_0_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_3 = io_request_0_ready & io_request_0_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1; // @[Reg.scala 16:16]
  reg [31:0] c2; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_1 = io_request_0_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step; // @[Reg.scala 16:16]
  reg [31:0] price; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T = $signed(price) * $signed(c1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T = $signed(rng_io_g1_bits) * $signed(c2); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T = $signed(price) * $signed(partial_res2); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_2 = $signed(partial_res3) + $signed(partial_res1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_3 = counter == last_step ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_4 = counter == last_step ? counter : _counter_T_1; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_7 = io_response_0_ready & io_response_0_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_5 = _T_7 ? 3'h1 : state; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_6 = 3'h5 == state ? _GEN_5 : state; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_7 = 3'h4 == state ? $signed(_price_T_2) : $signed(price); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_3 : _GEN_6; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_9 = 3'h4 == state ? _GEN_4 : counter; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_64 = {$signed(partial_res3), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_10 = 3'h3 == state ? $signed(_partial_res3_T) : $signed({{12{_GEN_64[51]}},_GEN_64}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_11 = 3'h3 == state ? 3'h4 : _GEN_8; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_65 = {$signed(partial_res1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_14 = 3'h2 == state ? $signed(_partial_res1_T) : $signed({{12{_GEN_65[51]}},_GEN_65}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_66 = {$signed(partial_res2), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_15 = 3'h2 == state ? $signed(_partial_res2_T) : $signed({{20{_GEN_66[63]}},_GEN_66}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_17 = 3'h2 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_10); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_23 = 3'h1 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_14); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_24 = 3'h1 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_15); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_25 = 3'h1 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_17); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_29 = 3'h0 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_23); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_30 = 3'h0 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_24); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_31 = 3'h0 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_25); // @[MonteCarlo.scala 66:19 60:27]
  reg [2:0] state_1; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_6 = $signed(io_request_1_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_7 = io_request_1_ready & io_request_1_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1_1; // @[Reg.scala 16:16]
  reg [31:0] c2_1; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_4 = io_request_1_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step_1; // @[Reg.scala 16:16]
  reg [31:0] price_1; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1_1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2_1; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3_1; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter_1; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T_1 = $signed(price_1) * $signed(c1_1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T_1 = $signed(rng_io_g2_bits) * $signed(c2_1); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T_1 = $signed(price_1) * $signed(partial_res2_1); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_5 = $signed(partial_res3_1) + $signed(partial_res1_1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_35 = counter_1 == last_step_1 ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_36 = counter_1 == last_step_1 ? counter_1 : _counter_T_3; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_15 = io_response_1_ready & io_response_1_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_37 = _T_15 ? 3'h1 : state_1; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_38 = 3'h5 == state_1 ? _GEN_37 : state_1; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_39 = 3'h4 == state_1 ? $signed(_price_T_5) : $signed(price_1); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_40 = 3'h4 == state_1 ? _GEN_35 : _GEN_38; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_41 = 3'h4 == state_1 ? _GEN_36 : counter_1; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_74 = {$signed(partial_res3_1), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_42 = 3'h3 == state_1 ? $signed(_partial_res3_T_1) : $signed({{12{_GEN_74[51]}},_GEN_74}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_43 = 3'h3 == state_1 ? 3'h4 : _GEN_40; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_75 = {$signed(partial_res1_1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_46 = 3'h2 == state_1 ? $signed(_partial_res1_T_1) : $signed({{12{_GEN_75[51]}},_GEN_75}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_76 = {$signed(partial_res2_1), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_47 = 3'h2 == state_1 ? $signed(_partial_res2_T_1) : $signed({{20{_GEN_76[63]}},_GEN_76}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_49 = 3'h2 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_42); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_55 = 3'h1 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_46); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_56 = 3'h1 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_47); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_57 = 3'h1 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_49); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_61 = 3'h0 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_55); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_62 = 3'h0 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_56); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_63 = 3'h0 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_57); // @[MonteCarlo.scala 66:19 60:27]
  wire [43:0] _GEN_84 = _GEN_29[63:20];
  wire [51:0] _GEN_86 = _GEN_30[83:32];
  wire [43:0] _GEN_88 = _GEN_31[63:20];
  wire [43:0] _GEN_90 = _GEN_61[63:20];
  wire [51:0] _GEN_92 = _GEN_62[83:32];
  wire [43:0] _GEN_94 = _GEN_63[63:20];
  BoxMuller_1 rng ( // @[MonteCarlo.scala 42:19]
    .clock(rng_clock),
    .reset(rng_reset),
    .io_g1_valid(rng_io_g1_valid),
    .io_g1_bits(rng_io_g1_bits),
    .io_g2_valid(rng_io_g2_valid),
    .io_g2_bits(rng_io_g2_bits)
  );
  assign io_request_0_ready = state == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_request_1_ready = state_1 == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_response_0_valid = state == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_0_bits = price; // @[MonteCarlo.scala 65:16]
  assign io_response_1_valid = state_1 == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_1_bits = price_1; // @[MonteCarlo.scala 65:16]
  assign rng_clock = clock;
  assign rng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state <= 3'h1;
      end else begin
        state <= 3'h0;
      end
    end else if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_3) begin // @[MonteCarlo.scala 71:23]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[MonteCarlo.scala 66:19]
      state <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state <= _GEN_11;
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c1 <= _c1_T_2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c2 <= io_request_0_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      last_step <= _last_step_T_1; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        price <= io_request_0_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          price <= _GEN_7;
        end
      end
    end
    partial_res1 <= _GEN_84[31:0];
    partial_res2 <= _GEN_86[31:0];
    partial_res3 <= _GEN_88[31:0];
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        counter <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          counter <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state_1 <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state_1 <= 3'h1;
      end else begin
        state_1 <= 3'h0;
      end
    end else if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_7) begin // @[MonteCarlo.scala 71:23]
        state_1 <= 3'h2;
      end else begin
        state_1 <= 3'h1;
      end
    end else if (3'h2 == state_1) begin // @[MonteCarlo.scala 66:19]
      state_1 <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state_1 <= _GEN_43;
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c1_1 <= _c1_T_6; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c2_1 <= io_request_1_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      last_step_1 <= _last_step_T_4; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        price_1 <= io_request_1_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          price_1 <= _GEN_39;
        end
      end
    end
    partial_res1_1 <= _GEN_90[31:0];
    partial_res2_1 <= _GEN_92[31:0];
    partial_res3_1 <= _GEN_94[31:0];
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        counter_1 <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          counter_1 <= _GEN_41;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  c1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_step = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  price = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  partial_res1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  partial_res2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  partial_res3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  c1_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_step_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  price_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  partial_res1_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  partial_res2_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  partial_res3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  counter_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_4(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h18a6f088 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h273bfa53 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h3f07a4cb : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_5(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h3ee683d6 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h384486c2 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h17a2c41 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoxMuller_2(
  input         clock,
  input         reset,
  output        io_g1_valid,
  output [51:0] io_g1_bits,
  output        io_g2_valid,
  output [51:0] io_g2_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [95:0] _RAND_77;
`endif // RANDOMIZE_REG_INIT
  wire  rng1_clock; // @[BoxMuller.scala 51:20]
  wire  rng1_reset; // @[BoxMuller.scala 51:20]
  wire  rng1_io_rand_valid; // @[BoxMuller.scala 51:20]
  wire [31:0] rng1_io_rand_bits; // @[BoxMuller.scala 51:20]
  wire  rng2_clock; // @[BoxMuller.scala 52:20]
  wire  rng2_reset; // @[BoxMuller.scala 52:20]
  wire  rng2_io_rand_valid; // @[BoxMuller.scala 52:20]
  wire [31:0] rng2_io_rand_bits; // @[BoxMuller.scala 52:20]
  wire  trigonometric_clock; // @[BoxMuller.scala 55:29]
  wire  trigonometric_reset; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_theta_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_theta_bits; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_result_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_sine; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_cosine; // @[BoxMuller.scala 55:29]
  wire  sqrt_log_clock; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_reset; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_uniform_valid; // @[BoxMuller.scala 84:24]
  wire [31:0] sqrt_log_io_uniform_bits; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_result_valid; // @[BoxMuller.scala 84:24]
  wire [51:0] sqrt_log_io_result_bits; // @[BoxMuller.scala 84:24]
  wire [30:0] _theta_T_3 = {2'h0,rng1_io_rand_bits[28:0]}; // @[BoxMuller.scala 62:18]
  wire [62:0] _theta_T_4 = $signed(_theta_T_3) * 32'sh6487ed51; // @[BoxMuller.scala 62:26]
  reg  quadrantPipe_valid; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_1; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_1; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_2; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_2; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_3; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_3; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_4; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_4; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_5; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_5; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_6; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_6; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_7; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_7; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_8; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_8; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_9; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_9; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_10; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_10; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_11; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_11; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_12; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_12; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_13; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_13; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_14; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_14; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_15; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_15; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_16; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_16; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_17; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_17; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_18; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_18; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_19; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_19; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_20; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_20; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_21; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_21; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_22; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_22; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_23; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_23; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_24; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_24; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_25; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_25; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_26; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_26; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_27; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_27; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_28; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_28; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_29; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_29; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_30; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_30; // @[Reg.scala 16:16]
  reg [1:0] quadrantPipe_bits_31; // @[Reg.scala 16:16]
  reg  trigonometric_io_theta_v; // @[Valid.scala 127:22]
  reg [31:0] trigonometric_io_theta_b; // @[Reg.scala 16:16]
  wire [33:0] _GEN_40 = _theta_T_4[62:29]; // @[BoxMuller.scala 59:19 61:9]
  wire [31:0] theta = _GEN_40[31:0]; // @[BoxMuller.scala 59:19 61:9]
  wire  _cosine_T = quadrantPipe_bits_31 == 2'h0; // @[BoxMuller.scala 70:21]
  wire  _cosine_T_2 = quadrantPipe_bits_31 == 2'h0 | quadrantPipe_bits_31 == 2'h3; // @[BoxMuller.scala 70:29]
  wire [31:0] _cosine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_cosine); // @[BoxMuller.scala 72:7]
  reg  cosinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] cosinePipe_bits; // @[Reg.scala 16:16]
  wire  _sine_T_2 = _cosine_T | quadrantPipe_bits_31 == 2'h2; // @[BoxMuller.scala 78:29]
  wire [31:0] _sine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_sine); // @[BoxMuller.scala 80:7]
  reg  sinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] sinePipe_bits; // @[Reg.scala 16:16]
  reg  signPipe_bits; // @[Reg.scala 16:16]
  wire [28:0] _sqrt_log_io_uniform_T_1 = rng2_io_rand_bits[28:0]; // @[BoxMuller.scala 87:89]
  reg  sqrt_log_io_uniform_v; // @[Valid.scala 127:22]
  reg [28:0] sqrt_log_io_uniform_b; // @[Reg.scala 16:16]
  wire [51:0] _sign_adjusted_T_3 = 52'sh0 - $signed(sqrt_log_io_result_bits); // @[BoxMuller.scala 93:7]
  reg  sign_adjustedPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] sign_adjustedPipe_bits; // @[Reg.scala 16:16]
  wire  _io_g1_T = sign_adjustedPipe_valid & cosinePipe_valid; // @[BoxMuller.scala 99:25]
  wire [83:0] _io_g1_T_1 = $signed(cosinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 100:17]
  reg  io_g1_v; // @[Valid.scala 127:22]
  reg [83:0] io_g1_b; // @[Reg.scala 16:16]
  wire  _io_g2_T = sign_adjustedPipe_valid & sinePipe_valid; // @[BoxMuller.scala 103:25]
  wire [83:0] _io_g2_T_1 = $signed(sinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 104:15]
  reg  io_g2_v; // @[Valid.scala 127:22]
  reg [83:0] io_g2_b; // @[Reg.scala 16:16]
  wire [53:0] _GEN_42 = io_g1_b[83:30]; // @[BoxMuller.scala 98:9]
  wire [53:0] _GEN_44 = io_g2_b[83:30]; // @[BoxMuller.scala 102:9]
  wire [32:0] _GEN_46 = {$signed(trigonometric_io_theta_b), 1'h0}; // @[BoxMuller.scala 65:26]
  TauswortheUniform_4 rng1 ( // @[BoxMuller.scala 51:20]
    .clock(rng1_clock),
    .reset(rng1_reset),
    .io_rand_valid(rng1_io_rand_valid),
    .io_rand_bits(rng1_io_rand_bits)
  );
  TauswortheUniform_5 rng2 ( // @[BoxMuller.scala 52:20]
    .clock(rng2_clock),
    .reset(rng2_reset),
    .io_rand_valid(rng2_io_rand_valid),
    .io_rand_bits(rng2_io_rand_bits)
  );
  Trigonometric trigonometric ( // @[BoxMuller.scala 55:29]
    .clock(trigonometric_clock),
    .reset(trigonometric_reset),
    .io_theta_valid(trigonometric_io_theta_valid),
    .io_theta_bits(trigonometric_io_theta_bits),
    .io_result_valid(trigonometric_io_result_valid),
    .io_result_bits_sine(trigonometric_io_result_bits_sine),
    .io_result_bits_cosine(trigonometric_io_result_bits_cosine)
  );
  SquareRootLog sqrt_log ( // @[BoxMuller.scala 84:24]
    .clock(sqrt_log_clock),
    .reset(sqrt_log_reset),
    .io_uniform_valid(sqrt_log_io_uniform_valid),
    .io_uniform_bits(sqrt_log_io_uniform_bits),
    .io_result_valid(sqrt_log_io_result_valid),
    .io_result_bits(sqrt_log_io_result_bits)
  );
  assign io_g1_valid = io_g1_v; // @[Valid.scala 122:21 123:17]
  assign io_g1_bits = _GEN_42[51:0]; // @[BoxMuller.scala 98:9]
  assign io_g2_valid = io_g2_v; // @[Valid.scala 122:21 123:17]
  assign io_g2_bits = _GEN_44[51:0]; // @[BoxMuller.scala 102:9]
  assign rng1_clock = clock;
  assign rng1_reset = reset;
  assign rng2_clock = clock;
  assign rng2_reset = reset;
  assign trigonometric_clock = clock;
  assign trigonometric_reset = reset;
  assign trigonometric_io_theta_valid = trigonometric_io_theta_v; // @[Valid.scala 122:21 123:17]
  assign trigonometric_io_theta_bits = _GEN_46[31:0]; // @[BoxMuller.scala 65:26]
  assign sqrt_log_clock = clock;
  assign sqrt_log_reset = reset;
  assign sqrt_log_io_uniform_valid = sqrt_log_io_uniform_v; // @[Valid.scala 122:21 123:17]
  assign sqrt_log_io_uniform_bits = {{3{sqrt_log_io_uniform_b[28]}},sqrt_log_io_uniform_b}; // @[BoxMuller.scala 87:23]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits <= rng1_io_rand_bits[31:30]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_1 <= quadrantPipe_valid; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_1 <= quadrantPipe_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_2 <= quadrantPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_1) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_2 <= quadrantPipe_bits_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_3 <= quadrantPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_2) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_3 <= quadrantPipe_bits_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_4 <= quadrantPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_3) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_4 <= quadrantPipe_bits_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_5 <= quadrantPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_4) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_5 <= quadrantPipe_bits_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_6 <= quadrantPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_5) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_6 <= quadrantPipe_bits_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_7 <= quadrantPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_6) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_7 <= quadrantPipe_bits_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_8 <= quadrantPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_7) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_8 <= quadrantPipe_bits_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_9 <= quadrantPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_8) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_9 <= quadrantPipe_bits_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_10 <= quadrantPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_9) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_10 <= quadrantPipe_bits_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_11 <= quadrantPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_10) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_11 <= quadrantPipe_bits_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_12 <= quadrantPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_11) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_12 <= quadrantPipe_bits_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_13 <= quadrantPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_12) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_13 <= quadrantPipe_bits_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_14 <= quadrantPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_13) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_14 <= quadrantPipe_bits_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_15 <= quadrantPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_14) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_15 <= quadrantPipe_bits_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_16 <= quadrantPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_15) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_16 <= quadrantPipe_bits_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_17 <= quadrantPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_16) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_17 <= quadrantPipe_bits_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_18 <= quadrantPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_17) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_18 <= quadrantPipe_bits_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_19 <= quadrantPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_18) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_19 <= quadrantPipe_bits_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_20 <= quadrantPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_19) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_20 <= quadrantPipe_bits_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_21 <= quadrantPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_20) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_21 <= quadrantPipe_bits_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_22 <= quadrantPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_21) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_22 <= quadrantPipe_bits_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_23 <= quadrantPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_22) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_23 <= quadrantPipe_bits_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_24 <= quadrantPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_23) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_24 <= quadrantPipe_bits_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_25 <= quadrantPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_24) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_25 <= quadrantPipe_bits_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_26 <= quadrantPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_25) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_26 <= quadrantPipe_bits_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_27 <= quadrantPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_26) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_27 <= quadrantPipe_bits_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_28 <= quadrantPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_27) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_28 <= quadrantPipe_bits_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_29 <= quadrantPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_28) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_29 <= quadrantPipe_bits_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_30 <= quadrantPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_29) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_30 <= quadrantPipe_bits_29; // @[Reg.scala 17:22]
    end
    if (quadrantPipe_valid_30) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_31 <= quadrantPipe_bits_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      trigonometric_io_theta_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      trigonometric_io_theta_v <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      trigonometric_io_theta_b <= theta; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      cosinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      cosinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_cosine_T_2) begin // @[BoxMuller.scala 69:8]
        cosinePipe_bits <= trigonometric_io_result_bits_cosine;
      end else begin
        cosinePipe_bits <= _cosine_T_5;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      sinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_sine_T_2) begin // @[BoxMuller.scala 77:8]
        sinePipe_bits <= trigonometric_io_result_bits_sine;
      end else begin
        sinePipe_bits <= _sine_T_5;
      end
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      signPipe_bits <= rng2_io_rand_bits[31]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sqrt_log_io_uniform_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sqrt_log_io_uniform_v <= rng2_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      sqrt_log_io_uniform_b <= _sqrt_log_io_uniform_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sign_adjustedPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sign_adjustedPipe_valid <= sqrt_log_io_result_valid; // @[Valid.scala 127:22]
    end
    if (sqrt_log_io_result_valid) begin // @[Reg.scala 17:18]
      if (signPipe_bits) begin // @[BoxMuller.scala 91:8]
        sign_adjustedPipe_bits <= _sign_adjusted_T_3;
      end else begin
        sign_adjustedPipe_bits <= sqrt_log_io_result_bits;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g1_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g1_v <= _io_g1_T; // @[Valid.scala 127:22]
    end
    if (_io_g1_T) begin // @[Reg.scala 17:18]
      io_g1_b <= _io_g1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g2_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g2_v <= _io_g2_T; // @[Valid.scala 127:22]
    end
    if (_io_g2_T) begin // @[Reg.scala 17:18]
      io_g2_b <= _io_g2_T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quadrantPipe_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  quadrantPipe_bits = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  quadrantPipe_valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  quadrantPipe_bits_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  quadrantPipe_valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  quadrantPipe_bits_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  quadrantPipe_valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quadrantPipe_bits_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  quadrantPipe_valid_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  quadrantPipe_bits_4 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  quadrantPipe_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  quadrantPipe_bits_5 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  quadrantPipe_valid_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  quadrantPipe_bits_6 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  quadrantPipe_valid_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  quadrantPipe_bits_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  quadrantPipe_valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  quadrantPipe_bits_8 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  quadrantPipe_valid_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  quadrantPipe_bits_9 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  quadrantPipe_valid_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  quadrantPipe_bits_10 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  quadrantPipe_valid_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  quadrantPipe_bits_11 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  quadrantPipe_valid_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  quadrantPipe_bits_12 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  quadrantPipe_valid_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  quadrantPipe_bits_13 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  quadrantPipe_valid_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  quadrantPipe_bits_14 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  quadrantPipe_valid_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  quadrantPipe_bits_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  quadrantPipe_valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  quadrantPipe_bits_16 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  quadrantPipe_valid_17 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  quadrantPipe_bits_17 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  quadrantPipe_valid_18 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  quadrantPipe_bits_18 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  quadrantPipe_valid_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  quadrantPipe_bits_19 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  quadrantPipe_valid_20 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  quadrantPipe_bits_20 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  quadrantPipe_valid_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  quadrantPipe_bits_21 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  quadrantPipe_valid_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  quadrantPipe_bits_22 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  quadrantPipe_valid_23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  quadrantPipe_bits_23 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  quadrantPipe_valid_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  quadrantPipe_bits_24 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  quadrantPipe_valid_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  quadrantPipe_bits_25 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  quadrantPipe_valid_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  quadrantPipe_bits_26 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  quadrantPipe_valid_27 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  quadrantPipe_bits_27 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  quadrantPipe_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  quadrantPipe_bits_28 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  quadrantPipe_valid_29 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  quadrantPipe_bits_29 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  quadrantPipe_valid_30 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  quadrantPipe_bits_30 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  quadrantPipe_bits_31 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  trigonometric_io_theta_v = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  trigonometric_io_theta_b = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cosinePipe_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cosinePipe_bits = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sinePipe_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sinePipe_bits = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  signPipe_bits = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sqrt_log_io_uniform_v = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sqrt_log_io_uniform_b = _RAND_71[28:0];
  _RAND_72 = {1{`RANDOM}};
  sign_adjustedPipe_valid = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  sign_adjustedPipe_bits = _RAND_73[51:0];
  _RAND_74 = {1{`RANDOM}};
  io_g1_v = _RAND_74[0:0];
  _RAND_75 = {3{`RANDOM}};
  io_g1_b = _RAND_75[83:0];
  _RAND_76 = {1{`RANDOM}};
  io_g2_v = _RAND_76[0:0];
  _RAND_77 = {3{`RANDOM}};
  io_g2_b = _RAND_77[83:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MonteCarlo_2(
  input         clock,
  input         reset,
  output        io_request_0_ready,
  input         io_request_0_valid,
  input  [31:0] io_request_0_bits_time_steps,
  input  [31:0] io_request_0_bits_start_value,
  input  [31:0] io_request_0_bits_coefficient1,
  input  [31:0] io_request_0_bits_coefficient2,
  output        io_request_1_ready,
  input         io_request_1_valid,
  input  [31:0] io_request_1_bits_time_steps,
  input  [31:0] io_request_1_bits_start_value,
  input  [31:0] io_request_1_bits_coefficient1,
  input  [31:0] io_request_1_bits_coefficient2,
  input         io_response_0_ready,
  output        io_response_0_valid,
  output [31:0] io_response_0_bits,
  input         io_response_1_ready,
  output        io_response_1_valid,
  output [31:0] io_response_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rng_clock; // @[MonteCarlo.scala 42:19]
  wire  rng_reset; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g1_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g1_bits; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g2_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g2_bits; // @[MonteCarlo.scala 42:19]
  wire  initialized = rng_io_g1_valid & rng_io_g2_valid; // @[MonteCarlo.scala 47:37]
  reg [2:0] state; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_2 = $signed(io_request_0_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_3 = io_request_0_ready & io_request_0_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1; // @[Reg.scala 16:16]
  reg [31:0] c2; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_1 = io_request_0_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step; // @[Reg.scala 16:16]
  reg [31:0] price; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T = $signed(price) * $signed(c1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T = $signed(rng_io_g1_bits) * $signed(c2); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T = $signed(price) * $signed(partial_res2); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_2 = $signed(partial_res3) + $signed(partial_res1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_3 = counter == last_step ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_4 = counter == last_step ? counter : _counter_T_1; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_7 = io_response_0_ready & io_response_0_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_5 = _T_7 ? 3'h1 : state; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_6 = 3'h5 == state ? _GEN_5 : state; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_7 = 3'h4 == state ? $signed(_price_T_2) : $signed(price); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_3 : _GEN_6; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_9 = 3'h4 == state ? _GEN_4 : counter; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_64 = {$signed(partial_res3), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_10 = 3'h3 == state ? $signed(_partial_res3_T) : $signed({{12{_GEN_64[51]}},_GEN_64}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_11 = 3'h3 == state ? 3'h4 : _GEN_8; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_65 = {$signed(partial_res1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_14 = 3'h2 == state ? $signed(_partial_res1_T) : $signed({{12{_GEN_65[51]}},_GEN_65}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_66 = {$signed(partial_res2), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_15 = 3'h2 == state ? $signed(_partial_res2_T) : $signed({{20{_GEN_66[63]}},_GEN_66}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_17 = 3'h2 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_10); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_23 = 3'h1 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_14); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_24 = 3'h1 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_15); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_25 = 3'h1 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_17); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_29 = 3'h0 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_23); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_30 = 3'h0 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_24); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_31 = 3'h0 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_25); // @[MonteCarlo.scala 66:19 60:27]
  reg [2:0] state_1; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_6 = $signed(io_request_1_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_7 = io_request_1_ready & io_request_1_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1_1; // @[Reg.scala 16:16]
  reg [31:0] c2_1; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_4 = io_request_1_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step_1; // @[Reg.scala 16:16]
  reg [31:0] price_1; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1_1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2_1; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3_1; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter_1; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T_1 = $signed(price_1) * $signed(c1_1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T_1 = $signed(rng_io_g2_bits) * $signed(c2_1); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T_1 = $signed(price_1) * $signed(partial_res2_1); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_5 = $signed(partial_res3_1) + $signed(partial_res1_1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_35 = counter_1 == last_step_1 ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_36 = counter_1 == last_step_1 ? counter_1 : _counter_T_3; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_15 = io_response_1_ready & io_response_1_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_37 = _T_15 ? 3'h1 : state_1; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_38 = 3'h5 == state_1 ? _GEN_37 : state_1; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_39 = 3'h4 == state_1 ? $signed(_price_T_5) : $signed(price_1); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_40 = 3'h4 == state_1 ? _GEN_35 : _GEN_38; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_41 = 3'h4 == state_1 ? _GEN_36 : counter_1; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_74 = {$signed(partial_res3_1), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_42 = 3'h3 == state_1 ? $signed(_partial_res3_T_1) : $signed({{12{_GEN_74[51]}},_GEN_74}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_43 = 3'h3 == state_1 ? 3'h4 : _GEN_40; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_75 = {$signed(partial_res1_1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_46 = 3'h2 == state_1 ? $signed(_partial_res1_T_1) : $signed({{12{_GEN_75[51]}},_GEN_75}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_76 = {$signed(partial_res2_1), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_47 = 3'h2 == state_1 ? $signed(_partial_res2_T_1) : $signed({{20{_GEN_76[63]}},_GEN_76}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_49 = 3'h2 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_42); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_55 = 3'h1 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_46); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_56 = 3'h1 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_47); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_57 = 3'h1 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_49); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_61 = 3'h0 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_55); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_62 = 3'h0 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_56); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_63 = 3'h0 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_57); // @[MonteCarlo.scala 66:19 60:27]
  wire [43:0] _GEN_84 = _GEN_29[63:20];
  wire [51:0] _GEN_86 = _GEN_30[83:32];
  wire [43:0] _GEN_88 = _GEN_31[63:20];
  wire [43:0] _GEN_90 = _GEN_61[63:20];
  wire [51:0] _GEN_92 = _GEN_62[83:32];
  wire [43:0] _GEN_94 = _GEN_63[63:20];
  BoxMuller_2 rng ( // @[MonteCarlo.scala 42:19]
    .clock(rng_clock),
    .reset(rng_reset),
    .io_g1_valid(rng_io_g1_valid),
    .io_g1_bits(rng_io_g1_bits),
    .io_g2_valid(rng_io_g2_valid),
    .io_g2_bits(rng_io_g2_bits)
  );
  assign io_request_0_ready = state == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_request_1_ready = state_1 == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_response_0_valid = state == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_0_bits = price; // @[MonteCarlo.scala 65:16]
  assign io_response_1_valid = state_1 == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_1_bits = price_1; // @[MonteCarlo.scala 65:16]
  assign rng_clock = clock;
  assign rng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state <= 3'h1;
      end else begin
        state <= 3'h0;
      end
    end else if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_3) begin // @[MonteCarlo.scala 71:23]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[MonteCarlo.scala 66:19]
      state <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state <= _GEN_11;
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c1 <= _c1_T_2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c2 <= io_request_0_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      last_step <= _last_step_T_1; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        price <= io_request_0_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          price <= _GEN_7;
        end
      end
    end
    partial_res1 <= _GEN_84[31:0];
    partial_res2 <= _GEN_86[31:0];
    partial_res3 <= _GEN_88[31:0];
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        counter <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          counter <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state_1 <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state_1 <= 3'h1;
      end else begin
        state_1 <= 3'h0;
      end
    end else if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_7) begin // @[MonteCarlo.scala 71:23]
        state_1 <= 3'h2;
      end else begin
        state_1 <= 3'h1;
      end
    end else if (3'h2 == state_1) begin // @[MonteCarlo.scala 66:19]
      state_1 <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state_1 <= _GEN_43;
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c1_1 <= _c1_T_6; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c2_1 <= io_request_1_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      last_step_1 <= _last_step_T_4; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        price_1 <= io_request_1_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          price_1 <= _GEN_39;
        end
      end
    end
    partial_res1_1 <= _GEN_90[31:0];
    partial_res2_1 <= _GEN_92[31:0];
    partial_res3_1 <= _GEN_94[31:0];
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        counter_1 <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          counter_1 <= _GEN_41;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  c1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_step = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  price = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  partial_res1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  partial_res2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  partial_res3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  c1_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_step_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  price_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  partial_res1_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  partial_res2_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  partial_res3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  counter_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_6(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h3c3d6d3c : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'hb43343c : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h1198d883 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_7(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h1407249c : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h83fd9d6 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h178cea3d : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoxMuller_3(
  input         clock,
  input         reset,
  output        io_g1_valid,
  output [51:0] io_g1_bits,
  output        io_g2_valid,
  output [51:0] io_g2_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [95:0] _RAND_77;
`endif // RANDOMIZE_REG_INIT
  wire  rng1_clock; // @[BoxMuller.scala 51:20]
  wire  rng1_reset; // @[BoxMuller.scala 51:20]
  wire  rng1_io_rand_valid; // @[BoxMuller.scala 51:20]
  wire [31:0] rng1_io_rand_bits; // @[BoxMuller.scala 51:20]
  wire  rng2_clock; // @[BoxMuller.scala 52:20]
  wire  rng2_reset; // @[BoxMuller.scala 52:20]
  wire  rng2_io_rand_valid; // @[BoxMuller.scala 52:20]
  wire [31:0] rng2_io_rand_bits; // @[BoxMuller.scala 52:20]
  wire  trigonometric_clock; // @[BoxMuller.scala 55:29]
  wire  trigonometric_reset; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_theta_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_theta_bits; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_result_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_sine; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_cosine; // @[BoxMuller.scala 55:29]
  wire  sqrt_log_clock; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_reset; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_uniform_valid; // @[BoxMuller.scala 84:24]
  wire [31:0] sqrt_log_io_uniform_bits; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_result_valid; // @[BoxMuller.scala 84:24]
  wire [51:0] sqrt_log_io_result_bits; // @[BoxMuller.scala 84:24]
  wire [30:0] _theta_T_3 = {2'h0,rng1_io_rand_bits[28:0]}; // @[BoxMuller.scala 62:18]
  wire [62:0] _theta_T_4 = $signed(_theta_T_3) * 32'sh6487ed51; // @[BoxMuller.scala 62:26]
  reg  quadrantPipe_valid; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_1; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_1; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_2; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_2; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_3; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_3; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_4; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_4; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_5; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_5; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_6; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_6; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_7; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_7; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_8; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_8; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_9; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_9; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_10; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_10; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_11; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_11; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_12; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_12; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_13; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_13; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_14; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_14; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_15; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_15; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_16; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_16; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_17; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_17; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_18; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_18; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_19; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_19; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_20; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_20; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_21; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_21; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_22; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_22; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_23; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_23; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_24; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_24; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_25; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_25; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_26; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_26; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_27; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_27; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_28; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_28; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_29; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_29; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_30; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_30; // @[Reg.scala 16:16]
  reg [1:0] quadrantPipe_bits_31; // @[Reg.scala 16:16]
  reg  trigonometric_io_theta_v; // @[Valid.scala 127:22]
  reg [31:0] trigonometric_io_theta_b; // @[Reg.scala 16:16]
  wire [33:0] _GEN_40 = _theta_T_4[62:29]; // @[BoxMuller.scala 59:19 61:9]
  wire [31:0] theta = _GEN_40[31:0]; // @[BoxMuller.scala 59:19 61:9]
  wire  _cosine_T = quadrantPipe_bits_31 == 2'h0; // @[BoxMuller.scala 70:21]
  wire  _cosine_T_2 = quadrantPipe_bits_31 == 2'h0 | quadrantPipe_bits_31 == 2'h3; // @[BoxMuller.scala 70:29]
  wire [31:0] _cosine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_cosine); // @[BoxMuller.scala 72:7]
  reg  cosinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] cosinePipe_bits; // @[Reg.scala 16:16]
  wire  _sine_T_2 = _cosine_T | quadrantPipe_bits_31 == 2'h2; // @[BoxMuller.scala 78:29]
  wire [31:0] _sine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_sine); // @[BoxMuller.scala 80:7]
  reg  sinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] sinePipe_bits; // @[Reg.scala 16:16]
  reg  signPipe_bits; // @[Reg.scala 16:16]
  wire [28:0] _sqrt_log_io_uniform_T_1 = rng2_io_rand_bits[28:0]; // @[BoxMuller.scala 87:89]
  reg  sqrt_log_io_uniform_v; // @[Valid.scala 127:22]
  reg [28:0] sqrt_log_io_uniform_b; // @[Reg.scala 16:16]
  wire [51:0] _sign_adjusted_T_3 = 52'sh0 - $signed(sqrt_log_io_result_bits); // @[BoxMuller.scala 93:7]
  reg  sign_adjustedPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] sign_adjustedPipe_bits; // @[Reg.scala 16:16]
  wire  _io_g1_T = sign_adjustedPipe_valid & cosinePipe_valid; // @[BoxMuller.scala 99:25]
  wire [83:0] _io_g1_T_1 = $signed(cosinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 100:17]
  reg  io_g1_v; // @[Valid.scala 127:22]
  reg [83:0] io_g1_b; // @[Reg.scala 16:16]
  wire  _io_g2_T = sign_adjustedPipe_valid & sinePipe_valid; // @[BoxMuller.scala 103:25]
  wire [83:0] _io_g2_T_1 = $signed(sinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 104:15]
  reg  io_g2_v; // @[Valid.scala 127:22]
  reg [83:0] io_g2_b; // @[Reg.scala 16:16]
  wire [53:0] _GEN_42 = io_g1_b[83:30]; // @[BoxMuller.scala 98:9]
  wire [53:0] _GEN_44 = io_g2_b[83:30]; // @[BoxMuller.scala 102:9]
  wire [32:0] _GEN_46 = {$signed(trigonometric_io_theta_b), 1'h0}; // @[BoxMuller.scala 65:26]
  TauswortheUniform_6 rng1 ( // @[BoxMuller.scala 51:20]
    .clock(rng1_clock),
    .reset(rng1_reset),
    .io_rand_valid(rng1_io_rand_valid),
    .io_rand_bits(rng1_io_rand_bits)
  );
  TauswortheUniform_7 rng2 ( // @[BoxMuller.scala 52:20]
    .clock(rng2_clock),
    .reset(rng2_reset),
    .io_rand_valid(rng2_io_rand_valid),
    .io_rand_bits(rng2_io_rand_bits)
  );
  Trigonometric trigonometric ( // @[BoxMuller.scala 55:29]
    .clock(trigonometric_clock),
    .reset(trigonometric_reset),
    .io_theta_valid(trigonometric_io_theta_valid),
    .io_theta_bits(trigonometric_io_theta_bits),
    .io_result_valid(trigonometric_io_result_valid),
    .io_result_bits_sine(trigonometric_io_result_bits_sine),
    .io_result_bits_cosine(trigonometric_io_result_bits_cosine)
  );
  SquareRootLog sqrt_log ( // @[BoxMuller.scala 84:24]
    .clock(sqrt_log_clock),
    .reset(sqrt_log_reset),
    .io_uniform_valid(sqrt_log_io_uniform_valid),
    .io_uniform_bits(sqrt_log_io_uniform_bits),
    .io_result_valid(sqrt_log_io_result_valid),
    .io_result_bits(sqrt_log_io_result_bits)
  );
  assign io_g1_valid = io_g1_v; // @[Valid.scala 122:21 123:17]
  assign io_g1_bits = _GEN_42[51:0]; // @[BoxMuller.scala 98:9]
  assign io_g2_valid = io_g2_v; // @[Valid.scala 122:21 123:17]
  assign io_g2_bits = _GEN_44[51:0]; // @[BoxMuller.scala 102:9]
  assign rng1_clock = clock;
  assign rng1_reset = reset;
  assign rng2_clock = clock;
  assign rng2_reset = reset;
  assign trigonometric_clock = clock;
  assign trigonometric_reset = reset;
  assign trigonometric_io_theta_valid = trigonometric_io_theta_v; // @[Valid.scala 122:21 123:17]
  assign trigonometric_io_theta_bits = _GEN_46[31:0]; // @[BoxMuller.scala 65:26]
  assign sqrt_log_clock = clock;
  assign sqrt_log_reset = reset;
  assign sqrt_log_io_uniform_valid = sqrt_log_io_uniform_v; // @[Valid.scala 122:21 123:17]
  assign sqrt_log_io_uniform_bits = {{3{sqrt_log_io_uniform_b[28]}},sqrt_log_io_uniform_b}; // @[BoxMuller.scala 87:23]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits <= rng1_io_rand_bits[31:30]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_1 <= quadrantPipe_valid; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_1 <= quadrantPipe_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_2 <= quadrantPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_1) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_2 <= quadrantPipe_bits_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_3 <= quadrantPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_2) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_3 <= quadrantPipe_bits_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_4 <= quadrantPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_3) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_4 <= quadrantPipe_bits_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_5 <= quadrantPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_4) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_5 <= quadrantPipe_bits_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_6 <= quadrantPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_5) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_6 <= quadrantPipe_bits_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_7 <= quadrantPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_6) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_7 <= quadrantPipe_bits_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_8 <= quadrantPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_7) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_8 <= quadrantPipe_bits_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_9 <= quadrantPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_8) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_9 <= quadrantPipe_bits_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_10 <= quadrantPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_9) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_10 <= quadrantPipe_bits_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_11 <= quadrantPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_10) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_11 <= quadrantPipe_bits_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_12 <= quadrantPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_11) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_12 <= quadrantPipe_bits_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_13 <= quadrantPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_12) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_13 <= quadrantPipe_bits_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_14 <= quadrantPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_13) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_14 <= quadrantPipe_bits_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_15 <= quadrantPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_14) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_15 <= quadrantPipe_bits_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_16 <= quadrantPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_15) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_16 <= quadrantPipe_bits_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_17 <= quadrantPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_16) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_17 <= quadrantPipe_bits_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_18 <= quadrantPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_17) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_18 <= quadrantPipe_bits_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_19 <= quadrantPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_18) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_19 <= quadrantPipe_bits_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_20 <= quadrantPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_19) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_20 <= quadrantPipe_bits_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_21 <= quadrantPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_20) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_21 <= quadrantPipe_bits_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_22 <= quadrantPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_21) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_22 <= quadrantPipe_bits_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_23 <= quadrantPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_22) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_23 <= quadrantPipe_bits_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_24 <= quadrantPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_23) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_24 <= quadrantPipe_bits_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_25 <= quadrantPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_24) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_25 <= quadrantPipe_bits_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_26 <= quadrantPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_25) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_26 <= quadrantPipe_bits_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_27 <= quadrantPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_26) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_27 <= quadrantPipe_bits_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_28 <= quadrantPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_27) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_28 <= quadrantPipe_bits_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_29 <= quadrantPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_28) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_29 <= quadrantPipe_bits_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_30 <= quadrantPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_29) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_30 <= quadrantPipe_bits_29; // @[Reg.scala 17:22]
    end
    if (quadrantPipe_valid_30) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_31 <= quadrantPipe_bits_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      trigonometric_io_theta_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      trigonometric_io_theta_v <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      trigonometric_io_theta_b <= theta; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      cosinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      cosinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_cosine_T_2) begin // @[BoxMuller.scala 69:8]
        cosinePipe_bits <= trigonometric_io_result_bits_cosine;
      end else begin
        cosinePipe_bits <= _cosine_T_5;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      sinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_sine_T_2) begin // @[BoxMuller.scala 77:8]
        sinePipe_bits <= trigonometric_io_result_bits_sine;
      end else begin
        sinePipe_bits <= _sine_T_5;
      end
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      signPipe_bits <= rng2_io_rand_bits[31]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sqrt_log_io_uniform_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sqrt_log_io_uniform_v <= rng2_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      sqrt_log_io_uniform_b <= _sqrt_log_io_uniform_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sign_adjustedPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sign_adjustedPipe_valid <= sqrt_log_io_result_valid; // @[Valid.scala 127:22]
    end
    if (sqrt_log_io_result_valid) begin // @[Reg.scala 17:18]
      if (signPipe_bits) begin // @[BoxMuller.scala 91:8]
        sign_adjustedPipe_bits <= _sign_adjusted_T_3;
      end else begin
        sign_adjustedPipe_bits <= sqrt_log_io_result_bits;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g1_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g1_v <= _io_g1_T; // @[Valid.scala 127:22]
    end
    if (_io_g1_T) begin // @[Reg.scala 17:18]
      io_g1_b <= _io_g1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g2_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g2_v <= _io_g2_T; // @[Valid.scala 127:22]
    end
    if (_io_g2_T) begin // @[Reg.scala 17:18]
      io_g2_b <= _io_g2_T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quadrantPipe_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  quadrantPipe_bits = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  quadrantPipe_valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  quadrantPipe_bits_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  quadrantPipe_valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  quadrantPipe_bits_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  quadrantPipe_valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quadrantPipe_bits_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  quadrantPipe_valid_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  quadrantPipe_bits_4 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  quadrantPipe_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  quadrantPipe_bits_5 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  quadrantPipe_valid_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  quadrantPipe_bits_6 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  quadrantPipe_valid_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  quadrantPipe_bits_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  quadrantPipe_valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  quadrantPipe_bits_8 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  quadrantPipe_valid_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  quadrantPipe_bits_9 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  quadrantPipe_valid_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  quadrantPipe_bits_10 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  quadrantPipe_valid_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  quadrantPipe_bits_11 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  quadrantPipe_valid_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  quadrantPipe_bits_12 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  quadrantPipe_valid_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  quadrantPipe_bits_13 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  quadrantPipe_valid_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  quadrantPipe_bits_14 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  quadrantPipe_valid_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  quadrantPipe_bits_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  quadrantPipe_valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  quadrantPipe_bits_16 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  quadrantPipe_valid_17 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  quadrantPipe_bits_17 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  quadrantPipe_valid_18 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  quadrantPipe_bits_18 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  quadrantPipe_valid_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  quadrantPipe_bits_19 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  quadrantPipe_valid_20 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  quadrantPipe_bits_20 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  quadrantPipe_valid_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  quadrantPipe_bits_21 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  quadrantPipe_valid_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  quadrantPipe_bits_22 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  quadrantPipe_valid_23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  quadrantPipe_bits_23 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  quadrantPipe_valid_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  quadrantPipe_bits_24 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  quadrantPipe_valid_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  quadrantPipe_bits_25 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  quadrantPipe_valid_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  quadrantPipe_bits_26 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  quadrantPipe_valid_27 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  quadrantPipe_bits_27 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  quadrantPipe_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  quadrantPipe_bits_28 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  quadrantPipe_valid_29 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  quadrantPipe_bits_29 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  quadrantPipe_valid_30 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  quadrantPipe_bits_30 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  quadrantPipe_bits_31 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  trigonometric_io_theta_v = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  trigonometric_io_theta_b = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cosinePipe_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cosinePipe_bits = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sinePipe_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sinePipe_bits = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  signPipe_bits = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sqrt_log_io_uniform_v = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sqrt_log_io_uniform_b = _RAND_71[28:0];
  _RAND_72 = {1{`RANDOM}};
  sign_adjustedPipe_valid = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  sign_adjustedPipe_bits = _RAND_73[51:0];
  _RAND_74 = {1{`RANDOM}};
  io_g1_v = _RAND_74[0:0];
  _RAND_75 = {3{`RANDOM}};
  io_g1_b = _RAND_75[83:0];
  _RAND_76 = {1{`RANDOM}};
  io_g2_v = _RAND_76[0:0];
  _RAND_77 = {3{`RANDOM}};
  io_g2_b = _RAND_77[83:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MonteCarlo_3(
  input         clock,
  input         reset,
  output        io_request_0_ready,
  input         io_request_0_valid,
  input  [31:0] io_request_0_bits_time_steps,
  input  [31:0] io_request_0_bits_start_value,
  input  [31:0] io_request_0_bits_coefficient1,
  input  [31:0] io_request_0_bits_coefficient2,
  output        io_request_1_ready,
  input         io_request_1_valid,
  input  [31:0] io_request_1_bits_time_steps,
  input  [31:0] io_request_1_bits_start_value,
  input  [31:0] io_request_1_bits_coefficient1,
  input  [31:0] io_request_1_bits_coefficient2,
  input         io_response_0_ready,
  output        io_response_0_valid,
  output [31:0] io_response_0_bits,
  input         io_response_1_ready,
  output        io_response_1_valid,
  output [31:0] io_response_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rng_clock; // @[MonteCarlo.scala 42:19]
  wire  rng_reset; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g1_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g1_bits; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g2_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g2_bits; // @[MonteCarlo.scala 42:19]
  wire  initialized = rng_io_g1_valid & rng_io_g2_valid; // @[MonteCarlo.scala 47:37]
  reg [2:0] state; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_2 = $signed(io_request_0_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_3 = io_request_0_ready & io_request_0_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1; // @[Reg.scala 16:16]
  reg [31:0] c2; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_1 = io_request_0_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step; // @[Reg.scala 16:16]
  reg [31:0] price; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T = $signed(price) * $signed(c1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T = $signed(rng_io_g1_bits) * $signed(c2); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T = $signed(price) * $signed(partial_res2); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_2 = $signed(partial_res3) + $signed(partial_res1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_3 = counter == last_step ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_4 = counter == last_step ? counter : _counter_T_1; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_7 = io_response_0_ready & io_response_0_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_5 = _T_7 ? 3'h1 : state; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_6 = 3'h5 == state ? _GEN_5 : state; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_7 = 3'h4 == state ? $signed(_price_T_2) : $signed(price); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_3 : _GEN_6; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_9 = 3'h4 == state ? _GEN_4 : counter; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_64 = {$signed(partial_res3), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_10 = 3'h3 == state ? $signed(_partial_res3_T) : $signed({{12{_GEN_64[51]}},_GEN_64}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_11 = 3'h3 == state ? 3'h4 : _GEN_8; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_65 = {$signed(partial_res1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_14 = 3'h2 == state ? $signed(_partial_res1_T) : $signed({{12{_GEN_65[51]}},_GEN_65}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_66 = {$signed(partial_res2), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_15 = 3'h2 == state ? $signed(_partial_res2_T) : $signed({{20{_GEN_66[63]}},_GEN_66}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_17 = 3'h2 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_10); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_23 = 3'h1 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_14); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_24 = 3'h1 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_15); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_25 = 3'h1 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_17); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_29 = 3'h0 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_23); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_30 = 3'h0 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_24); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_31 = 3'h0 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_25); // @[MonteCarlo.scala 66:19 60:27]
  reg [2:0] state_1; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_6 = $signed(io_request_1_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_7 = io_request_1_ready & io_request_1_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1_1; // @[Reg.scala 16:16]
  reg [31:0] c2_1; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_4 = io_request_1_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step_1; // @[Reg.scala 16:16]
  reg [31:0] price_1; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1_1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2_1; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3_1; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter_1; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T_1 = $signed(price_1) * $signed(c1_1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T_1 = $signed(rng_io_g2_bits) * $signed(c2_1); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T_1 = $signed(price_1) * $signed(partial_res2_1); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_5 = $signed(partial_res3_1) + $signed(partial_res1_1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_35 = counter_1 == last_step_1 ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_36 = counter_1 == last_step_1 ? counter_1 : _counter_T_3; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_15 = io_response_1_ready & io_response_1_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_37 = _T_15 ? 3'h1 : state_1; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_38 = 3'h5 == state_1 ? _GEN_37 : state_1; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_39 = 3'h4 == state_1 ? $signed(_price_T_5) : $signed(price_1); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_40 = 3'h4 == state_1 ? _GEN_35 : _GEN_38; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_41 = 3'h4 == state_1 ? _GEN_36 : counter_1; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_74 = {$signed(partial_res3_1), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_42 = 3'h3 == state_1 ? $signed(_partial_res3_T_1) : $signed({{12{_GEN_74[51]}},_GEN_74}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_43 = 3'h3 == state_1 ? 3'h4 : _GEN_40; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_75 = {$signed(partial_res1_1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_46 = 3'h2 == state_1 ? $signed(_partial_res1_T_1) : $signed({{12{_GEN_75[51]}},_GEN_75}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_76 = {$signed(partial_res2_1), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_47 = 3'h2 == state_1 ? $signed(_partial_res2_T_1) : $signed({{20{_GEN_76[63]}},_GEN_76}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_49 = 3'h2 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_42); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_55 = 3'h1 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_46); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_56 = 3'h1 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_47); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_57 = 3'h1 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_49); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_61 = 3'h0 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_55); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_62 = 3'h0 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_56); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_63 = 3'h0 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_57); // @[MonteCarlo.scala 66:19 60:27]
  wire [43:0] _GEN_84 = _GEN_29[63:20];
  wire [51:0] _GEN_86 = _GEN_30[83:32];
  wire [43:0] _GEN_88 = _GEN_31[63:20];
  wire [43:0] _GEN_90 = _GEN_61[63:20];
  wire [51:0] _GEN_92 = _GEN_62[83:32];
  wire [43:0] _GEN_94 = _GEN_63[63:20];
  BoxMuller_3 rng ( // @[MonteCarlo.scala 42:19]
    .clock(rng_clock),
    .reset(rng_reset),
    .io_g1_valid(rng_io_g1_valid),
    .io_g1_bits(rng_io_g1_bits),
    .io_g2_valid(rng_io_g2_valid),
    .io_g2_bits(rng_io_g2_bits)
  );
  assign io_request_0_ready = state == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_request_1_ready = state_1 == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_response_0_valid = state == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_0_bits = price; // @[MonteCarlo.scala 65:16]
  assign io_response_1_valid = state_1 == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_1_bits = price_1; // @[MonteCarlo.scala 65:16]
  assign rng_clock = clock;
  assign rng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state <= 3'h1;
      end else begin
        state <= 3'h0;
      end
    end else if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_3) begin // @[MonteCarlo.scala 71:23]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[MonteCarlo.scala 66:19]
      state <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state <= _GEN_11;
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c1 <= _c1_T_2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c2 <= io_request_0_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      last_step <= _last_step_T_1; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        price <= io_request_0_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          price <= _GEN_7;
        end
      end
    end
    partial_res1 <= _GEN_84[31:0];
    partial_res2 <= _GEN_86[31:0];
    partial_res3 <= _GEN_88[31:0];
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        counter <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          counter <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state_1 <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state_1 <= 3'h1;
      end else begin
        state_1 <= 3'h0;
      end
    end else if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_7) begin // @[MonteCarlo.scala 71:23]
        state_1 <= 3'h2;
      end else begin
        state_1 <= 3'h1;
      end
    end else if (3'h2 == state_1) begin // @[MonteCarlo.scala 66:19]
      state_1 <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state_1 <= _GEN_43;
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c1_1 <= _c1_T_6; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c2_1 <= io_request_1_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      last_step_1 <= _last_step_T_4; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        price_1 <= io_request_1_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          price_1 <= _GEN_39;
        end
      end
    end
    partial_res1_1 <= _GEN_90[31:0];
    partial_res2_1 <= _GEN_92[31:0];
    partial_res3_1 <= _GEN_94[31:0];
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        counter_1 <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          counter_1 <= _GEN_41;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  c1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_step = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  price = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  partial_res1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  partial_res2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  partial_res3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  c1_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_step_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  price_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  partial_res1_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  partial_res2_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  partial_res3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  counter_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_8(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h961ebe6 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h2d21954e : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h17cbbc7 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_9(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h16b82d : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h22fdc8c2 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h9723d7 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoxMuller_4(
  input         clock,
  input         reset,
  output        io_g1_valid,
  output [51:0] io_g1_bits,
  output        io_g2_valid,
  output [51:0] io_g2_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [95:0] _RAND_77;
`endif // RANDOMIZE_REG_INIT
  wire  rng1_clock; // @[BoxMuller.scala 51:20]
  wire  rng1_reset; // @[BoxMuller.scala 51:20]
  wire  rng1_io_rand_valid; // @[BoxMuller.scala 51:20]
  wire [31:0] rng1_io_rand_bits; // @[BoxMuller.scala 51:20]
  wire  rng2_clock; // @[BoxMuller.scala 52:20]
  wire  rng2_reset; // @[BoxMuller.scala 52:20]
  wire  rng2_io_rand_valid; // @[BoxMuller.scala 52:20]
  wire [31:0] rng2_io_rand_bits; // @[BoxMuller.scala 52:20]
  wire  trigonometric_clock; // @[BoxMuller.scala 55:29]
  wire  trigonometric_reset; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_theta_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_theta_bits; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_result_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_sine; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_cosine; // @[BoxMuller.scala 55:29]
  wire  sqrt_log_clock; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_reset; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_uniform_valid; // @[BoxMuller.scala 84:24]
  wire [31:0] sqrt_log_io_uniform_bits; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_result_valid; // @[BoxMuller.scala 84:24]
  wire [51:0] sqrt_log_io_result_bits; // @[BoxMuller.scala 84:24]
  wire [30:0] _theta_T_3 = {2'h0,rng1_io_rand_bits[28:0]}; // @[BoxMuller.scala 62:18]
  wire [62:0] _theta_T_4 = $signed(_theta_T_3) * 32'sh6487ed51; // @[BoxMuller.scala 62:26]
  reg  quadrantPipe_valid; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_1; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_1; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_2; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_2; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_3; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_3; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_4; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_4; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_5; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_5; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_6; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_6; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_7; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_7; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_8; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_8; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_9; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_9; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_10; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_10; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_11; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_11; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_12; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_12; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_13; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_13; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_14; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_14; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_15; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_15; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_16; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_16; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_17; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_17; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_18; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_18; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_19; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_19; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_20; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_20; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_21; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_21; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_22; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_22; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_23; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_23; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_24; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_24; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_25; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_25; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_26; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_26; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_27; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_27; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_28; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_28; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_29; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_29; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_30; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_30; // @[Reg.scala 16:16]
  reg [1:0] quadrantPipe_bits_31; // @[Reg.scala 16:16]
  reg  trigonometric_io_theta_v; // @[Valid.scala 127:22]
  reg [31:0] trigonometric_io_theta_b; // @[Reg.scala 16:16]
  wire [33:0] _GEN_40 = _theta_T_4[62:29]; // @[BoxMuller.scala 59:19 61:9]
  wire [31:0] theta = _GEN_40[31:0]; // @[BoxMuller.scala 59:19 61:9]
  wire  _cosine_T = quadrantPipe_bits_31 == 2'h0; // @[BoxMuller.scala 70:21]
  wire  _cosine_T_2 = quadrantPipe_bits_31 == 2'h0 | quadrantPipe_bits_31 == 2'h3; // @[BoxMuller.scala 70:29]
  wire [31:0] _cosine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_cosine); // @[BoxMuller.scala 72:7]
  reg  cosinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] cosinePipe_bits; // @[Reg.scala 16:16]
  wire  _sine_T_2 = _cosine_T | quadrantPipe_bits_31 == 2'h2; // @[BoxMuller.scala 78:29]
  wire [31:0] _sine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_sine); // @[BoxMuller.scala 80:7]
  reg  sinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] sinePipe_bits; // @[Reg.scala 16:16]
  reg  signPipe_bits; // @[Reg.scala 16:16]
  wire [28:0] _sqrt_log_io_uniform_T_1 = rng2_io_rand_bits[28:0]; // @[BoxMuller.scala 87:89]
  reg  sqrt_log_io_uniform_v; // @[Valid.scala 127:22]
  reg [28:0] sqrt_log_io_uniform_b; // @[Reg.scala 16:16]
  wire [51:0] _sign_adjusted_T_3 = 52'sh0 - $signed(sqrt_log_io_result_bits); // @[BoxMuller.scala 93:7]
  reg  sign_adjustedPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] sign_adjustedPipe_bits; // @[Reg.scala 16:16]
  wire  _io_g1_T = sign_adjustedPipe_valid & cosinePipe_valid; // @[BoxMuller.scala 99:25]
  wire [83:0] _io_g1_T_1 = $signed(cosinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 100:17]
  reg  io_g1_v; // @[Valid.scala 127:22]
  reg [83:0] io_g1_b; // @[Reg.scala 16:16]
  wire  _io_g2_T = sign_adjustedPipe_valid & sinePipe_valid; // @[BoxMuller.scala 103:25]
  wire [83:0] _io_g2_T_1 = $signed(sinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 104:15]
  reg  io_g2_v; // @[Valid.scala 127:22]
  reg [83:0] io_g2_b; // @[Reg.scala 16:16]
  wire [53:0] _GEN_42 = io_g1_b[83:30]; // @[BoxMuller.scala 98:9]
  wire [53:0] _GEN_44 = io_g2_b[83:30]; // @[BoxMuller.scala 102:9]
  wire [32:0] _GEN_46 = {$signed(trigonometric_io_theta_b), 1'h0}; // @[BoxMuller.scala 65:26]
  TauswortheUniform_8 rng1 ( // @[BoxMuller.scala 51:20]
    .clock(rng1_clock),
    .reset(rng1_reset),
    .io_rand_valid(rng1_io_rand_valid),
    .io_rand_bits(rng1_io_rand_bits)
  );
  TauswortheUniform_9 rng2 ( // @[BoxMuller.scala 52:20]
    .clock(rng2_clock),
    .reset(rng2_reset),
    .io_rand_valid(rng2_io_rand_valid),
    .io_rand_bits(rng2_io_rand_bits)
  );
  Trigonometric trigonometric ( // @[BoxMuller.scala 55:29]
    .clock(trigonometric_clock),
    .reset(trigonometric_reset),
    .io_theta_valid(trigonometric_io_theta_valid),
    .io_theta_bits(trigonometric_io_theta_bits),
    .io_result_valid(trigonometric_io_result_valid),
    .io_result_bits_sine(trigonometric_io_result_bits_sine),
    .io_result_bits_cosine(trigonometric_io_result_bits_cosine)
  );
  SquareRootLog sqrt_log ( // @[BoxMuller.scala 84:24]
    .clock(sqrt_log_clock),
    .reset(sqrt_log_reset),
    .io_uniform_valid(sqrt_log_io_uniform_valid),
    .io_uniform_bits(sqrt_log_io_uniform_bits),
    .io_result_valid(sqrt_log_io_result_valid),
    .io_result_bits(sqrt_log_io_result_bits)
  );
  assign io_g1_valid = io_g1_v; // @[Valid.scala 122:21 123:17]
  assign io_g1_bits = _GEN_42[51:0]; // @[BoxMuller.scala 98:9]
  assign io_g2_valid = io_g2_v; // @[Valid.scala 122:21 123:17]
  assign io_g2_bits = _GEN_44[51:0]; // @[BoxMuller.scala 102:9]
  assign rng1_clock = clock;
  assign rng1_reset = reset;
  assign rng2_clock = clock;
  assign rng2_reset = reset;
  assign trigonometric_clock = clock;
  assign trigonometric_reset = reset;
  assign trigonometric_io_theta_valid = trigonometric_io_theta_v; // @[Valid.scala 122:21 123:17]
  assign trigonometric_io_theta_bits = _GEN_46[31:0]; // @[BoxMuller.scala 65:26]
  assign sqrt_log_clock = clock;
  assign sqrt_log_reset = reset;
  assign sqrt_log_io_uniform_valid = sqrt_log_io_uniform_v; // @[Valid.scala 122:21 123:17]
  assign sqrt_log_io_uniform_bits = {{3{sqrt_log_io_uniform_b[28]}},sqrt_log_io_uniform_b}; // @[BoxMuller.scala 87:23]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits <= rng1_io_rand_bits[31:30]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_1 <= quadrantPipe_valid; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_1 <= quadrantPipe_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_2 <= quadrantPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_1) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_2 <= quadrantPipe_bits_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_3 <= quadrantPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_2) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_3 <= quadrantPipe_bits_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_4 <= quadrantPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_3) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_4 <= quadrantPipe_bits_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_5 <= quadrantPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_4) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_5 <= quadrantPipe_bits_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_6 <= quadrantPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_5) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_6 <= quadrantPipe_bits_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_7 <= quadrantPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_6) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_7 <= quadrantPipe_bits_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_8 <= quadrantPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_7) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_8 <= quadrantPipe_bits_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_9 <= quadrantPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_8) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_9 <= quadrantPipe_bits_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_10 <= quadrantPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_9) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_10 <= quadrantPipe_bits_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_11 <= quadrantPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_10) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_11 <= quadrantPipe_bits_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_12 <= quadrantPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_11) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_12 <= quadrantPipe_bits_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_13 <= quadrantPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_12) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_13 <= quadrantPipe_bits_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_14 <= quadrantPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_13) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_14 <= quadrantPipe_bits_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_15 <= quadrantPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_14) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_15 <= quadrantPipe_bits_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_16 <= quadrantPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_15) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_16 <= quadrantPipe_bits_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_17 <= quadrantPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_16) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_17 <= quadrantPipe_bits_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_18 <= quadrantPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_17) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_18 <= quadrantPipe_bits_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_19 <= quadrantPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_18) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_19 <= quadrantPipe_bits_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_20 <= quadrantPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_19) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_20 <= quadrantPipe_bits_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_21 <= quadrantPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_20) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_21 <= quadrantPipe_bits_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_22 <= quadrantPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_21) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_22 <= quadrantPipe_bits_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_23 <= quadrantPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_22) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_23 <= quadrantPipe_bits_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_24 <= quadrantPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_23) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_24 <= quadrantPipe_bits_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_25 <= quadrantPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_24) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_25 <= quadrantPipe_bits_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_26 <= quadrantPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_25) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_26 <= quadrantPipe_bits_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_27 <= quadrantPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_26) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_27 <= quadrantPipe_bits_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_28 <= quadrantPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_27) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_28 <= quadrantPipe_bits_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_29 <= quadrantPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_28) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_29 <= quadrantPipe_bits_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_30 <= quadrantPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_29) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_30 <= quadrantPipe_bits_29; // @[Reg.scala 17:22]
    end
    if (quadrantPipe_valid_30) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_31 <= quadrantPipe_bits_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      trigonometric_io_theta_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      trigonometric_io_theta_v <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      trigonometric_io_theta_b <= theta; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      cosinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      cosinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_cosine_T_2) begin // @[BoxMuller.scala 69:8]
        cosinePipe_bits <= trigonometric_io_result_bits_cosine;
      end else begin
        cosinePipe_bits <= _cosine_T_5;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      sinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_sine_T_2) begin // @[BoxMuller.scala 77:8]
        sinePipe_bits <= trigonometric_io_result_bits_sine;
      end else begin
        sinePipe_bits <= _sine_T_5;
      end
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      signPipe_bits <= rng2_io_rand_bits[31]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sqrt_log_io_uniform_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sqrt_log_io_uniform_v <= rng2_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      sqrt_log_io_uniform_b <= _sqrt_log_io_uniform_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sign_adjustedPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sign_adjustedPipe_valid <= sqrt_log_io_result_valid; // @[Valid.scala 127:22]
    end
    if (sqrt_log_io_result_valid) begin // @[Reg.scala 17:18]
      if (signPipe_bits) begin // @[BoxMuller.scala 91:8]
        sign_adjustedPipe_bits <= _sign_adjusted_T_3;
      end else begin
        sign_adjustedPipe_bits <= sqrt_log_io_result_bits;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g1_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g1_v <= _io_g1_T; // @[Valid.scala 127:22]
    end
    if (_io_g1_T) begin // @[Reg.scala 17:18]
      io_g1_b <= _io_g1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g2_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g2_v <= _io_g2_T; // @[Valid.scala 127:22]
    end
    if (_io_g2_T) begin // @[Reg.scala 17:18]
      io_g2_b <= _io_g2_T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quadrantPipe_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  quadrantPipe_bits = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  quadrantPipe_valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  quadrantPipe_bits_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  quadrantPipe_valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  quadrantPipe_bits_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  quadrantPipe_valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quadrantPipe_bits_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  quadrantPipe_valid_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  quadrantPipe_bits_4 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  quadrantPipe_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  quadrantPipe_bits_5 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  quadrantPipe_valid_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  quadrantPipe_bits_6 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  quadrantPipe_valid_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  quadrantPipe_bits_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  quadrantPipe_valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  quadrantPipe_bits_8 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  quadrantPipe_valid_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  quadrantPipe_bits_9 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  quadrantPipe_valid_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  quadrantPipe_bits_10 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  quadrantPipe_valid_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  quadrantPipe_bits_11 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  quadrantPipe_valid_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  quadrantPipe_bits_12 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  quadrantPipe_valid_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  quadrantPipe_bits_13 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  quadrantPipe_valid_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  quadrantPipe_bits_14 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  quadrantPipe_valid_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  quadrantPipe_bits_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  quadrantPipe_valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  quadrantPipe_bits_16 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  quadrantPipe_valid_17 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  quadrantPipe_bits_17 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  quadrantPipe_valid_18 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  quadrantPipe_bits_18 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  quadrantPipe_valid_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  quadrantPipe_bits_19 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  quadrantPipe_valid_20 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  quadrantPipe_bits_20 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  quadrantPipe_valid_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  quadrantPipe_bits_21 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  quadrantPipe_valid_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  quadrantPipe_bits_22 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  quadrantPipe_valid_23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  quadrantPipe_bits_23 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  quadrantPipe_valid_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  quadrantPipe_bits_24 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  quadrantPipe_valid_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  quadrantPipe_bits_25 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  quadrantPipe_valid_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  quadrantPipe_bits_26 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  quadrantPipe_valid_27 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  quadrantPipe_bits_27 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  quadrantPipe_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  quadrantPipe_bits_28 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  quadrantPipe_valid_29 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  quadrantPipe_bits_29 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  quadrantPipe_valid_30 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  quadrantPipe_bits_30 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  quadrantPipe_bits_31 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  trigonometric_io_theta_v = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  trigonometric_io_theta_b = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cosinePipe_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cosinePipe_bits = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sinePipe_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sinePipe_bits = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  signPipe_bits = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sqrt_log_io_uniform_v = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sqrt_log_io_uniform_b = _RAND_71[28:0];
  _RAND_72 = {1{`RANDOM}};
  sign_adjustedPipe_valid = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  sign_adjustedPipe_bits = _RAND_73[51:0];
  _RAND_74 = {1{`RANDOM}};
  io_g1_v = _RAND_74[0:0];
  _RAND_75 = {3{`RANDOM}};
  io_g1_b = _RAND_75[83:0];
  _RAND_76 = {1{`RANDOM}};
  io_g2_v = _RAND_76[0:0];
  _RAND_77 = {3{`RANDOM}};
  io_g2_b = _RAND_77[83:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MonteCarlo_4(
  input         clock,
  input         reset,
  output        io_request_0_ready,
  input         io_request_0_valid,
  input  [31:0] io_request_0_bits_time_steps,
  input  [31:0] io_request_0_bits_start_value,
  input  [31:0] io_request_0_bits_coefficient1,
  input  [31:0] io_request_0_bits_coefficient2,
  output        io_request_1_ready,
  input         io_request_1_valid,
  input  [31:0] io_request_1_bits_time_steps,
  input  [31:0] io_request_1_bits_start_value,
  input  [31:0] io_request_1_bits_coefficient1,
  input  [31:0] io_request_1_bits_coefficient2,
  input         io_response_0_ready,
  output        io_response_0_valid,
  output [31:0] io_response_0_bits,
  input         io_response_1_ready,
  output        io_response_1_valid,
  output [31:0] io_response_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rng_clock; // @[MonteCarlo.scala 42:19]
  wire  rng_reset; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g1_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g1_bits; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g2_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g2_bits; // @[MonteCarlo.scala 42:19]
  wire  initialized = rng_io_g1_valid & rng_io_g2_valid; // @[MonteCarlo.scala 47:37]
  reg [2:0] state; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_2 = $signed(io_request_0_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_3 = io_request_0_ready & io_request_0_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1; // @[Reg.scala 16:16]
  reg [31:0] c2; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_1 = io_request_0_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step; // @[Reg.scala 16:16]
  reg [31:0] price; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T = $signed(price) * $signed(c1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T = $signed(rng_io_g1_bits) * $signed(c2); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T = $signed(price) * $signed(partial_res2); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_2 = $signed(partial_res3) + $signed(partial_res1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_3 = counter == last_step ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_4 = counter == last_step ? counter : _counter_T_1; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_7 = io_response_0_ready & io_response_0_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_5 = _T_7 ? 3'h1 : state; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_6 = 3'h5 == state ? _GEN_5 : state; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_7 = 3'h4 == state ? $signed(_price_T_2) : $signed(price); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_3 : _GEN_6; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_9 = 3'h4 == state ? _GEN_4 : counter; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_64 = {$signed(partial_res3), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_10 = 3'h3 == state ? $signed(_partial_res3_T) : $signed({{12{_GEN_64[51]}},_GEN_64}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_11 = 3'h3 == state ? 3'h4 : _GEN_8; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_65 = {$signed(partial_res1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_14 = 3'h2 == state ? $signed(_partial_res1_T) : $signed({{12{_GEN_65[51]}},_GEN_65}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_66 = {$signed(partial_res2), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_15 = 3'h2 == state ? $signed(_partial_res2_T) : $signed({{20{_GEN_66[63]}},_GEN_66}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_17 = 3'h2 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_10); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_23 = 3'h1 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_14); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_24 = 3'h1 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_15); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_25 = 3'h1 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_17); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_29 = 3'h0 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_23); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_30 = 3'h0 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_24); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_31 = 3'h0 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_25); // @[MonteCarlo.scala 66:19 60:27]
  reg [2:0] state_1; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_6 = $signed(io_request_1_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_7 = io_request_1_ready & io_request_1_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1_1; // @[Reg.scala 16:16]
  reg [31:0] c2_1; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_4 = io_request_1_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step_1; // @[Reg.scala 16:16]
  reg [31:0] price_1; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1_1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2_1; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3_1; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter_1; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T_1 = $signed(price_1) * $signed(c1_1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T_1 = $signed(rng_io_g2_bits) * $signed(c2_1); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T_1 = $signed(price_1) * $signed(partial_res2_1); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_5 = $signed(partial_res3_1) + $signed(partial_res1_1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_35 = counter_1 == last_step_1 ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_36 = counter_1 == last_step_1 ? counter_1 : _counter_T_3; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_15 = io_response_1_ready & io_response_1_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_37 = _T_15 ? 3'h1 : state_1; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_38 = 3'h5 == state_1 ? _GEN_37 : state_1; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_39 = 3'h4 == state_1 ? $signed(_price_T_5) : $signed(price_1); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_40 = 3'h4 == state_1 ? _GEN_35 : _GEN_38; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_41 = 3'h4 == state_1 ? _GEN_36 : counter_1; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_74 = {$signed(partial_res3_1), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_42 = 3'h3 == state_1 ? $signed(_partial_res3_T_1) : $signed({{12{_GEN_74[51]}},_GEN_74}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_43 = 3'h3 == state_1 ? 3'h4 : _GEN_40; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_75 = {$signed(partial_res1_1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_46 = 3'h2 == state_1 ? $signed(_partial_res1_T_1) : $signed({{12{_GEN_75[51]}},_GEN_75}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_76 = {$signed(partial_res2_1), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_47 = 3'h2 == state_1 ? $signed(_partial_res2_T_1) : $signed({{20{_GEN_76[63]}},_GEN_76}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_49 = 3'h2 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_42); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_55 = 3'h1 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_46); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_56 = 3'h1 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_47); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_57 = 3'h1 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_49); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_61 = 3'h0 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_55); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_62 = 3'h0 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_56); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_63 = 3'h0 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_57); // @[MonteCarlo.scala 66:19 60:27]
  wire [43:0] _GEN_84 = _GEN_29[63:20];
  wire [51:0] _GEN_86 = _GEN_30[83:32];
  wire [43:0] _GEN_88 = _GEN_31[63:20];
  wire [43:0] _GEN_90 = _GEN_61[63:20];
  wire [51:0] _GEN_92 = _GEN_62[83:32];
  wire [43:0] _GEN_94 = _GEN_63[63:20];
  BoxMuller_4 rng ( // @[MonteCarlo.scala 42:19]
    .clock(rng_clock),
    .reset(rng_reset),
    .io_g1_valid(rng_io_g1_valid),
    .io_g1_bits(rng_io_g1_bits),
    .io_g2_valid(rng_io_g2_valid),
    .io_g2_bits(rng_io_g2_bits)
  );
  assign io_request_0_ready = state == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_request_1_ready = state_1 == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_response_0_valid = state == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_0_bits = price; // @[MonteCarlo.scala 65:16]
  assign io_response_1_valid = state_1 == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_1_bits = price_1; // @[MonteCarlo.scala 65:16]
  assign rng_clock = clock;
  assign rng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state <= 3'h1;
      end else begin
        state <= 3'h0;
      end
    end else if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_3) begin // @[MonteCarlo.scala 71:23]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[MonteCarlo.scala 66:19]
      state <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state <= _GEN_11;
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c1 <= _c1_T_2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c2 <= io_request_0_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      last_step <= _last_step_T_1; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        price <= io_request_0_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          price <= _GEN_7;
        end
      end
    end
    partial_res1 <= _GEN_84[31:0];
    partial_res2 <= _GEN_86[31:0];
    partial_res3 <= _GEN_88[31:0];
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        counter <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          counter <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state_1 <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state_1 <= 3'h1;
      end else begin
        state_1 <= 3'h0;
      end
    end else if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_7) begin // @[MonteCarlo.scala 71:23]
        state_1 <= 3'h2;
      end else begin
        state_1 <= 3'h1;
      end
    end else if (3'h2 == state_1) begin // @[MonteCarlo.scala 66:19]
      state_1 <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state_1 <= _GEN_43;
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c1_1 <= _c1_T_6; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c2_1 <= io_request_1_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      last_step_1 <= _last_step_T_4; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        price_1 <= io_request_1_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          price_1 <= _GEN_39;
        end
      end
    end
    partial_res1_1 <= _GEN_90[31:0];
    partial_res2_1 <= _GEN_92[31:0];
    partial_res3_1 <= _GEN_94[31:0];
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        counter_1 <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          counter_1 <= _GEN_41;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  c1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_step = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  price = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  partial_res1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  partial_res2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  partial_res3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  c1_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_step_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  price_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  partial_res1_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  partial_res2_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  partial_res3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  counter_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_10(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h3dba2710 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h24075e1e : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h6aff9b2 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_11(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h102f3cb9 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h280265e9 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h124c439b : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoxMuller_5(
  input         clock,
  input         reset,
  output        io_g1_valid,
  output [51:0] io_g1_bits,
  output        io_g2_valid,
  output [51:0] io_g2_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [95:0] _RAND_77;
`endif // RANDOMIZE_REG_INIT
  wire  rng1_clock; // @[BoxMuller.scala 51:20]
  wire  rng1_reset; // @[BoxMuller.scala 51:20]
  wire  rng1_io_rand_valid; // @[BoxMuller.scala 51:20]
  wire [31:0] rng1_io_rand_bits; // @[BoxMuller.scala 51:20]
  wire  rng2_clock; // @[BoxMuller.scala 52:20]
  wire  rng2_reset; // @[BoxMuller.scala 52:20]
  wire  rng2_io_rand_valid; // @[BoxMuller.scala 52:20]
  wire [31:0] rng2_io_rand_bits; // @[BoxMuller.scala 52:20]
  wire  trigonometric_clock; // @[BoxMuller.scala 55:29]
  wire  trigonometric_reset; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_theta_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_theta_bits; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_result_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_sine; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_cosine; // @[BoxMuller.scala 55:29]
  wire  sqrt_log_clock; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_reset; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_uniform_valid; // @[BoxMuller.scala 84:24]
  wire [31:0] sqrt_log_io_uniform_bits; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_result_valid; // @[BoxMuller.scala 84:24]
  wire [51:0] sqrt_log_io_result_bits; // @[BoxMuller.scala 84:24]
  wire [30:0] _theta_T_3 = {2'h0,rng1_io_rand_bits[28:0]}; // @[BoxMuller.scala 62:18]
  wire [62:0] _theta_T_4 = $signed(_theta_T_3) * 32'sh6487ed51; // @[BoxMuller.scala 62:26]
  reg  quadrantPipe_valid; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_1; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_1; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_2; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_2; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_3; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_3; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_4; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_4; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_5; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_5; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_6; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_6; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_7; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_7; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_8; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_8; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_9; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_9; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_10; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_10; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_11; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_11; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_12; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_12; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_13; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_13; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_14; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_14; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_15; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_15; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_16; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_16; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_17; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_17; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_18; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_18; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_19; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_19; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_20; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_20; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_21; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_21; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_22; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_22; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_23; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_23; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_24; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_24; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_25; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_25; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_26; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_26; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_27; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_27; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_28; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_28; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_29; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_29; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_30; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_30; // @[Reg.scala 16:16]
  reg [1:0] quadrantPipe_bits_31; // @[Reg.scala 16:16]
  reg  trigonometric_io_theta_v; // @[Valid.scala 127:22]
  reg [31:0] trigonometric_io_theta_b; // @[Reg.scala 16:16]
  wire [33:0] _GEN_40 = _theta_T_4[62:29]; // @[BoxMuller.scala 59:19 61:9]
  wire [31:0] theta = _GEN_40[31:0]; // @[BoxMuller.scala 59:19 61:9]
  wire  _cosine_T = quadrantPipe_bits_31 == 2'h0; // @[BoxMuller.scala 70:21]
  wire  _cosine_T_2 = quadrantPipe_bits_31 == 2'h0 | quadrantPipe_bits_31 == 2'h3; // @[BoxMuller.scala 70:29]
  wire [31:0] _cosine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_cosine); // @[BoxMuller.scala 72:7]
  reg  cosinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] cosinePipe_bits; // @[Reg.scala 16:16]
  wire  _sine_T_2 = _cosine_T | quadrantPipe_bits_31 == 2'h2; // @[BoxMuller.scala 78:29]
  wire [31:0] _sine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_sine); // @[BoxMuller.scala 80:7]
  reg  sinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] sinePipe_bits; // @[Reg.scala 16:16]
  reg  signPipe_bits; // @[Reg.scala 16:16]
  wire [28:0] _sqrt_log_io_uniform_T_1 = rng2_io_rand_bits[28:0]; // @[BoxMuller.scala 87:89]
  reg  sqrt_log_io_uniform_v; // @[Valid.scala 127:22]
  reg [28:0] sqrt_log_io_uniform_b; // @[Reg.scala 16:16]
  wire [51:0] _sign_adjusted_T_3 = 52'sh0 - $signed(sqrt_log_io_result_bits); // @[BoxMuller.scala 93:7]
  reg  sign_adjustedPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] sign_adjustedPipe_bits; // @[Reg.scala 16:16]
  wire  _io_g1_T = sign_adjustedPipe_valid & cosinePipe_valid; // @[BoxMuller.scala 99:25]
  wire [83:0] _io_g1_T_1 = $signed(cosinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 100:17]
  reg  io_g1_v; // @[Valid.scala 127:22]
  reg [83:0] io_g1_b; // @[Reg.scala 16:16]
  wire  _io_g2_T = sign_adjustedPipe_valid & sinePipe_valid; // @[BoxMuller.scala 103:25]
  wire [83:0] _io_g2_T_1 = $signed(sinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 104:15]
  reg  io_g2_v; // @[Valid.scala 127:22]
  reg [83:0] io_g2_b; // @[Reg.scala 16:16]
  wire [53:0] _GEN_42 = io_g1_b[83:30]; // @[BoxMuller.scala 98:9]
  wire [53:0] _GEN_44 = io_g2_b[83:30]; // @[BoxMuller.scala 102:9]
  wire [32:0] _GEN_46 = {$signed(trigonometric_io_theta_b), 1'h0}; // @[BoxMuller.scala 65:26]
  TauswortheUniform_10 rng1 ( // @[BoxMuller.scala 51:20]
    .clock(rng1_clock),
    .reset(rng1_reset),
    .io_rand_valid(rng1_io_rand_valid),
    .io_rand_bits(rng1_io_rand_bits)
  );
  TauswortheUniform_11 rng2 ( // @[BoxMuller.scala 52:20]
    .clock(rng2_clock),
    .reset(rng2_reset),
    .io_rand_valid(rng2_io_rand_valid),
    .io_rand_bits(rng2_io_rand_bits)
  );
  Trigonometric trigonometric ( // @[BoxMuller.scala 55:29]
    .clock(trigonometric_clock),
    .reset(trigonometric_reset),
    .io_theta_valid(trigonometric_io_theta_valid),
    .io_theta_bits(trigonometric_io_theta_bits),
    .io_result_valid(trigonometric_io_result_valid),
    .io_result_bits_sine(trigonometric_io_result_bits_sine),
    .io_result_bits_cosine(trigonometric_io_result_bits_cosine)
  );
  SquareRootLog sqrt_log ( // @[BoxMuller.scala 84:24]
    .clock(sqrt_log_clock),
    .reset(sqrt_log_reset),
    .io_uniform_valid(sqrt_log_io_uniform_valid),
    .io_uniform_bits(sqrt_log_io_uniform_bits),
    .io_result_valid(sqrt_log_io_result_valid),
    .io_result_bits(sqrt_log_io_result_bits)
  );
  assign io_g1_valid = io_g1_v; // @[Valid.scala 122:21 123:17]
  assign io_g1_bits = _GEN_42[51:0]; // @[BoxMuller.scala 98:9]
  assign io_g2_valid = io_g2_v; // @[Valid.scala 122:21 123:17]
  assign io_g2_bits = _GEN_44[51:0]; // @[BoxMuller.scala 102:9]
  assign rng1_clock = clock;
  assign rng1_reset = reset;
  assign rng2_clock = clock;
  assign rng2_reset = reset;
  assign trigonometric_clock = clock;
  assign trigonometric_reset = reset;
  assign trigonometric_io_theta_valid = trigonometric_io_theta_v; // @[Valid.scala 122:21 123:17]
  assign trigonometric_io_theta_bits = _GEN_46[31:0]; // @[BoxMuller.scala 65:26]
  assign sqrt_log_clock = clock;
  assign sqrt_log_reset = reset;
  assign sqrt_log_io_uniform_valid = sqrt_log_io_uniform_v; // @[Valid.scala 122:21 123:17]
  assign sqrt_log_io_uniform_bits = {{3{sqrt_log_io_uniform_b[28]}},sqrt_log_io_uniform_b}; // @[BoxMuller.scala 87:23]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits <= rng1_io_rand_bits[31:30]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_1 <= quadrantPipe_valid; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_1 <= quadrantPipe_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_2 <= quadrantPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_1) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_2 <= quadrantPipe_bits_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_3 <= quadrantPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_2) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_3 <= quadrantPipe_bits_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_4 <= quadrantPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_3) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_4 <= quadrantPipe_bits_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_5 <= quadrantPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_4) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_5 <= quadrantPipe_bits_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_6 <= quadrantPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_5) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_6 <= quadrantPipe_bits_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_7 <= quadrantPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_6) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_7 <= quadrantPipe_bits_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_8 <= quadrantPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_7) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_8 <= quadrantPipe_bits_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_9 <= quadrantPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_8) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_9 <= quadrantPipe_bits_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_10 <= quadrantPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_9) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_10 <= quadrantPipe_bits_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_11 <= quadrantPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_10) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_11 <= quadrantPipe_bits_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_12 <= quadrantPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_11) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_12 <= quadrantPipe_bits_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_13 <= quadrantPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_12) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_13 <= quadrantPipe_bits_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_14 <= quadrantPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_13) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_14 <= quadrantPipe_bits_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_15 <= quadrantPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_14) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_15 <= quadrantPipe_bits_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_16 <= quadrantPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_15) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_16 <= quadrantPipe_bits_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_17 <= quadrantPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_16) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_17 <= quadrantPipe_bits_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_18 <= quadrantPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_17) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_18 <= quadrantPipe_bits_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_19 <= quadrantPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_18) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_19 <= quadrantPipe_bits_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_20 <= quadrantPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_19) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_20 <= quadrantPipe_bits_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_21 <= quadrantPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_20) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_21 <= quadrantPipe_bits_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_22 <= quadrantPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_21) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_22 <= quadrantPipe_bits_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_23 <= quadrantPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_22) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_23 <= quadrantPipe_bits_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_24 <= quadrantPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_23) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_24 <= quadrantPipe_bits_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_25 <= quadrantPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_24) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_25 <= quadrantPipe_bits_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_26 <= quadrantPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_25) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_26 <= quadrantPipe_bits_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_27 <= quadrantPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_26) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_27 <= quadrantPipe_bits_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_28 <= quadrantPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_27) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_28 <= quadrantPipe_bits_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_29 <= quadrantPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_28) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_29 <= quadrantPipe_bits_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_30 <= quadrantPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_29) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_30 <= quadrantPipe_bits_29; // @[Reg.scala 17:22]
    end
    if (quadrantPipe_valid_30) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_31 <= quadrantPipe_bits_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      trigonometric_io_theta_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      trigonometric_io_theta_v <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      trigonometric_io_theta_b <= theta; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      cosinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      cosinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_cosine_T_2) begin // @[BoxMuller.scala 69:8]
        cosinePipe_bits <= trigonometric_io_result_bits_cosine;
      end else begin
        cosinePipe_bits <= _cosine_T_5;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      sinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_sine_T_2) begin // @[BoxMuller.scala 77:8]
        sinePipe_bits <= trigonometric_io_result_bits_sine;
      end else begin
        sinePipe_bits <= _sine_T_5;
      end
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      signPipe_bits <= rng2_io_rand_bits[31]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sqrt_log_io_uniform_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sqrt_log_io_uniform_v <= rng2_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      sqrt_log_io_uniform_b <= _sqrt_log_io_uniform_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sign_adjustedPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sign_adjustedPipe_valid <= sqrt_log_io_result_valid; // @[Valid.scala 127:22]
    end
    if (sqrt_log_io_result_valid) begin // @[Reg.scala 17:18]
      if (signPipe_bits) begin // @[BoxMuller.scala 91:8]
        sign_adjustedPipe_bits <= _sign_adjusted_T_3;
      end else begin
        sign_adjustedPipe_bits <= sqrt_log_io_result_bits;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g1_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g1_v <= _io_g1_T; // @[Valid.scala 127:22]
    end
    if (_io_g1_T) begin // @[Reg.scala 17:18]
      io_g1_b <= _io_g1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g2_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g2_v <= _io_g2_T; // @[Valid.scala 127:22]
    end
    if (_io_g2_T) begin // @[Reg.scala 17:18]
      io_g2_b <= _io_g2_T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quadrantPipe_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  quadrantPipe_bits = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  quadrantPipe_valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  quadrantPipe_bits_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  quadrantPipe_valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  quadrantPipe_bits_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  quadrantPipe_valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quadrantPipe_bits_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  quadrantPipe_valid_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  quadrantPipe_bits_4 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  quadrantPipe_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  quadrantPipe_bits_5 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  quadrantPipe_valid_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  quadrantPipe_bits_6 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  quadrantPipe_valid_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  quadrantPipe_bits_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  quadrantPipe_valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  quadrantPipe_bits_8 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  quadrantPipe_valid_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  quadrantPipe_bits_9 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  quadrantPipe_valid_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  quadrantPipe_bits_10 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  quadrantPipe_valid_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  quadrantPipe_bits_11 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  quadrantPipe_valid_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  quadrantPipe_bits_12 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  quadrantPipe_valid_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  quadrantPipe_bits_13 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  quadrantPipe_valid_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  quadrantPipe_bits_14 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  quadrantPipe_valid_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  quadrantPipe_bits_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  quadrantPipe_valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  quadrantPipe_bits_16 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  quadrantPipe_valid_17 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  quadrantPipe_bits_17 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  quadrantPipe_valid_18 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  quadrantPipe_bits_18 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  quadrantPipe_valid_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  quadrantPipe_bits_19 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  quadrantPipe_valid_20 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  quadrantPipe_bits_20 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  quadrantPipe_valid_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  quadrantPipe_bits_21 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  quadrantPipe_valid_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  quadrantPipe_bits_22 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  quadrantPipe_valid_23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  quadrantPipe_bits_23 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  quadrantPipe_valid_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  quadrantPipe_bits_24 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  quadrantPipe_valid_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  quadrantPipe_bits_25 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  quadrantPipe_valid_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  quadrantPipe_bits_26 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  quadrantPipe_valid_27 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  quadrantPipe_bits_27 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  quadrantPipe_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  quadrantPipe_bits_28 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  quadrantPipe_valid_29 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  quadrantPipe_bits_29 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  quadrantPipe_valid_30 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  quadrantPipe_bits_30 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  quadrantPipe_bits_31 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  trigonometric_io_theta_v = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  trigonometric_io_theta_b = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cosinePipe_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cosinePipe_bits = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sinePipe_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sinePipe_bits = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  signPipe_bits = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sqrt_log_io_uniform_v = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sqrt_log_io_uniform_b = _RAND_71[28:0];
  _RAND_72 = {1{`RANDOM}};
  sign_adjustedPipe_valid = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  sign_adjustedPipe_bits = _RAND_73[51:0];
  _RAND_74 = {1{`RANDOM}};
  io_g1_v = _RAND_74[0:0];
  _RAND_75 = {3{`RANDOM}};
  io_g1_b = _RAND_75[83:0];
  _RAND_76 = {1{`RANDOM}};
  io_g2_v = _RAND_76[0:0];
  _RAND_77 = {3{`RANDOM}};
  io_g2_b = _RAND_77[83:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MonteCarlo_5(
  input         clock,
  input         reset,
  output        io_request_0_ready,
  input         io_request_0_valid,
  input  [31:0] io_request_0_bits_time_steps,
  input  [31:0] io_request_0_bits_start_value,
  input  [31:0] io_request_0_bits_coefficient1,
  input  [31:0] io_request_0_bits_coefficient2,
  output        io_request_1_ready,
  input         io_request_1_valid,
  input  [31:0] io_request_1_bits_time_steps,
  input  [31:0] io_request_1_bits_start_value,
  input  [31:0] io_request_1_bits_coefficient1,
  input  [31:0] io_request_1_bits_coefficient2,
  input         io_response_0_ready,
  output        io_response_0_valid,
  output [31:0] io_response_0_bits,
  input         io_response_1_ready,
  output        io_response_1_valid,
  output [31:0] io_response_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rng_clock; // @[MonteCarlo.scala 42:19]
  wire  rng_reset; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g1_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g1_bits; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g2_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g2_bits; // @[MonteCarlo.scala 42:19]
  wire  initialized = rng_io_g1_valid & rng_io_g2_valid; // @[MonteCarlo.scala 47:37]
  reg [2:0] state; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_2 = $signed(io_request_0_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_3 = io_request_0_ready & io_request_0_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1; // @[Reg.scala 16:16]
  reg [31:0] c2; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_1 = io_request_0_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step; // @[Reg.scala 16:16]
  reg [31:0] price; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T = $signed(price) * $signed(c1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T = $signed(rng_io_g1_bits) * $signed(c2); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T = $signed(price) * $signed(partial_res2); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_2 = $signed(partial_res3) + $signed(partial_res1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_3 = counter == last_step ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_4 = counter == last_step ? counter : _counter_T_1; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_7 = io_response_0_ready & io_response_0_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_5 = _T_7 ? 3'h1 : state; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_6 = 3'h5 == state ? _GEN_5 : state; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_7 = 3'h4 == state ? $signed(_price_T_2) : $signed(price); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_3 : _GEN_6; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_9 = 3'h4 == state ? _GEN_4 : counter; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_64 = {$signed(partial_res3), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_10 = 3'h3 == state ? $signed(_partial_res3_T) : $signed({{12{_GEN_64[51]}},_GEN_64}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_11 = 3'h3 == state ? 3'h4 : _GEN_8; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_65 = {$signed(partial_res1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_14 = 3'h2 == state ? $signed(_partial_res1_T) : $signed({{12{_GEN_65[51]}},_GEN_65}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_66 = {$signed(partial_res2), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_15 = 3'h2 == state ? $signed(_partial_res2_T) : $signed({{20{_GEN_66[63]}},_GEN_66}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_17 = 3'h2 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_10); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_23 = 3'h1 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_14); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_24 = 3'h1 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_15); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_25 = 3'h1 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_17); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_29 = 3'h0 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_23); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_30 = 3'h0 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_24); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_31 = 3'h0 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_25); // @[MonteCarlo.scala 66:19 60:27]
  reg [2:0] state_1; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_6 = $signed(io_request_1_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_7 = io_request_1_ready & io_request_1_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1_1; // @[Reg.scala 16:16]
  reg [31:0] c2_1; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_4 = io_request_1_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step_1; // @[Reg.scala 16:16]
  reg [31:0] price_1; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1_1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2_1; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3_1; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter_1; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T_1 = $signed(price_1) * $signed(c1_1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T_1 = $signed(rng_io_g2_bits) * $signed(c2_1); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T_1 = $signed(price_1) * $signed(partial_res2_1); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_5 = $signed(partial_res3_1) + $signed(partial_res1_1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_35 = counter_1 == last_step_1 ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_36 = counter_1 == last_step_1 ? counter_1 : _counter_T_3; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_15 = io_response_1_ready & io_response_1_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_37 = _T_15 ? 3'h1 : state_1; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_38 = 3'h5 == state_1 ? _GEN_37 : state_1; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_39 = 3'h4 == state_1 ? $signed(_price_T_5) : $signed(price_1); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_40 = 3'h4 == state_1 ? _GEN_35 : _GEN_38; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_41 = 3'h4 == state_1 ? _GEN_36 : counter_1; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_74 = {$signed(partial_res3_1), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_42 = 3'h3 == state_1 ? $signed(_partial_res3_T_1) : $signed({{12{_GEN_74[51]}},_GEN_74}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_43 = 3'h3 == state_1 ? 3'h4 : _GEN_40; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_75 = {$signed(partial_res1_1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_46 = 3'h2 == state_1 ? $signed(_partial_res1_T_1) : $signed({{12{_GEN_75[51]}},_GEN_75}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_76 = {$signed(partial_res2_1), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_47 = 3'h2 == state_1 ? $signed(_partial_res2_T_1) : $signed({{20{_GEN_76[63]}},_GEN_76}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_49 = 3'h2 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_42); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_55 = 3'h1 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_46); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_56 = 3'h1 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_47); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_57 = 3'h1 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_49); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_61 = 3'h0 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_55); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_62 = 3'h0 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_56); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_63 = 3'h0 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_57); // @[MonteCarlo.scala 66:19 60:27]
  wire [43:0] _GEN_84 = _GEN_29[63:20];
  wire [51:0] _GEN_86 = _GEN_30[83:32];
  wire [43:0] _GEN_88 = _GEN_31[63:20];
  wire [43:0] _GEN_90 = _GEN_61[63:20];
  wire [51:0] _GEN_92 = _GEN_62[83:32];
  wire [43:0] _GEN_94 = _GEN_63[63:20];
  BoxMuller_5 rng ( // @[MonteCarlo.scala 42:19]
    .clock(rng_clock),
    .reset(rng_reset),
    .io_g1_valid(rng_io_g1_valid),
    .io_g1_bits(rng_io_g1_bits),
    .io_g2_valid(rng_io_g2_valid),
    .io_g2_bits(rng_io_g2_bits)
  );
  assign io_request_0_ready = state == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_request_1_ready = state_1 == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_response_0_valid = state == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_0_bits = price; // @[MonteCarlo.scala 65:16]
  assign io_response_1_valid = state_1 == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_1_bits = price_1; // @[MonteCarlo.scala 65:16]
  assign rng_clock = clock;
  assign rng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state <= 3'h1;
      end else begin
        state <= 3'h0;
      end
    end else if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_3) begin // @[MonteCarlo.scala 71:23]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[MonteCarlo.scala 66:19]
      state <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state <= _GEN_11;
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c1 <= _c1_T_2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c2 <= io_request_0_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      last_step <= _last_step_T_1; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        price <= io_request_0_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          price <= _GEN_7;
        end
      end
    end
    partial_res1 <= _GEN_84[31:0];
    partial_res2 <= _GEN_86[31:0];
    partial_res3 <= _GEN_88[31:0];
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        counter <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          counter <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state_1 <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state_1 <= 3'h1;
      end else begin
        state_1 <= 3'h0;
      end
    end else if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_7) begin // @[MonteCarlo.scala 71:23]
        state_1 <= 3'h2;
      end else begin
        state_1 <= 3'h1;
      end
    end else if (3'h2 == state_1) begin // @[MonteCarlo.scala 66:19]
      state_1 <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state_1 <= _GEN_43;
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c1_1 <= _c1_T_6; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c2_1 <= io_request_1_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      last_step_1 <= _last_step_T_4; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        price_1 <= io_request_1_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          price_1 <= _GEN_39;
        end
      end
    end
    partial_res1_1 <= _GEN_90[31:0];
    partial_res2_1 <= _GEN_92[31:0];
    partial_res3_1 <= _GEN_94[31:0];
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        counter_1 <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          counter_1 <= _GEN_41;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  c1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_step = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  price = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  partial_res1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  partial_res2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  partial_res3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  c1_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_step_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  price_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  partial_res1_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  partial_res2_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  partial_res3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  counter_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_12(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h1a4a7c26 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'hf490b2 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h31af19b9 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_13(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h3e8237a5 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h3f680080 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h2c0c08cb : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoxMuller_6(
  input         clock,
  input         reset,
  output        io_g1_valid,
  output [51:0] io_g1_bits,
  output        io_g2_valid,
  output [51:0] io_g2_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [95:0] _RAND_77;
`endif // RANDOMIZE_REG_INIT
  wire  rng1_clock; // @[BoxMuller.scala 51:20]
  wire  rng1_reset; // @[BoxMuller.scala 51:20]
  wire  rng1_io_rand_valid; // @[BoxMuller.scala 51:20]
  wire [31:0] rng1_io_rand_bits; // @[BoxMuller.scala 51:20]
  wire  rng2_clock; // @[BoxMuller.scala 52:20]
  wire  rng2_reset; // @[BoxMuller.scala 52:20]
  wire  rng2_io_rand_valid; // @[BoxMuller.scala 52:20]
  wire [31:0] rng2_io_rand_bits; // @[BoxMuller.scala 52:20]
  wire  trigonometric_clock; // @[BoxMuller.scala 55:29]
  wire  trigonometric_reset; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_theta_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_theta_bits; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_result_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_sine; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_cosine; // @[BoxMuller.scala 55:29]
  wire  sqrt_log_clock; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_reset; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_uniform_valid; // @[BoxMuller.scala 84:24]
  wire [31:0] sqrt_log_io_uniform_bits; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_result_valid; // @[BoxMuller.scala 84:24]
  wire [51:0] sqrt_log_io_result_bits; // @[BoxMuller.scala 84:24]
  wire [30:0] _theta_T_3 = {2'h0,rng1_io_rand_bits[28:0]}; // @[BoxMuller.scala 62:18]
  wire [62:0] _theta_T_4 = $signed(_theta_T_3) * 32'sh6487ed51; // @[BoxMuller.scala 62:26]
  reg  quadrantPipe_valid; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_1; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_1; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_2; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_2; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_3; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_3; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_4; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_4; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_5; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_5; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_6; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_6; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_7; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_7; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_8; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_8; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_9; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_9; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_10; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_10; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_11; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_11; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_12; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_12; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_13; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_13; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_14; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_14; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_15; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_15; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_16; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_16; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_17; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_17; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_18; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_18; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_19; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_19; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_20; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_20; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_21; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_21; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_22; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_22; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_23; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_23; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_24; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_24; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_25; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_25; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_26; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_26; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_27; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_27; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_28; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_28; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_29; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_29; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_30; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_30; // @[Reg.scala 16:16]
  reg [1:0] quadrantPipe_bits_31; // @[Reg.scala 16:16]
  reg  trigonometric_io_theta_v; // @[Valid.scala 127:22]
  reg [31:0] trigonometric_io_theta_b; // @[Reg.scala 16:16]
  wire [33:0] _GEN_40 = _theta_T_4[62:29]; // @[BoxMuller.scala 59:19 61:9]
  wire [31:0] theta = _GEN_40[31:0]; // @[BoxMuller.scala 59:19 61:9]
  wire  _cosine_T = quadrantPipe_bits_31 == 2'h0; // @[BoxMuller.scala 70:21]
  wire  _cosine_T_2 = quadrantPipe_bits_31 == 2'h0 | quadrantPipe_bits_31 == 2'h3; // @[BoxMuller.scala 70:29]
  wire [31:0] _cosine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_cosine); // @[BoxMuller.scala 72:7]
  reg  cosinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] cosinePipe_bits; // @[Reg.scala 16:16]
  wire  _sine_T_2 = _cosine_T | quadrantPipe_bits_31 == 2'h2; // @[BoxMuller.scala 78:29]
  wire [31:0] _sine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_sine); // @[BoxMuller.scala 80:7]
  reg  sinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] sinePipe_bits; // @[Reg.scala 16:16]
  reg  signPipe_bits; // @[Reg.scala 16:16]
  wire [28:0] _sqrt_log_io_uniform_T_1 = rng2_io_rand_bits[28:0]; // @[BoxMuller.scala 87:89]
  reg  sqrt_log_io_uniform_v; // @[Valid.scala 127:22]
  reg [28:0] sqrt_log_io_uniform_b; // @[Reg.scala 16:16]
  wire [51:0] _sign_adjusted_T_3 = 52'sh0 - $signed(sqrt_log_io_result_bits); // @[BoxMuller.scala 93:7]
  reg  sign_adjustedPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] sign_adjustedPipe_bits; // @[Reg.scala 16:16]
  wire  _io_g1_T = sign_adjustedPipe_valid & cosinePipe_valid; // @[BoxMuller.scala 99:25]
  wire [83:0] _io_g1_T_1 = $signed(cosinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 100:17]
  reg  io_g1_v; // @[Valid.scala 127:22]
  reg [83:0] io_g1_b; // @[Reg.scala 16:16]
  wire  _io_g2_T = sign_adjustedPipe_valid & sinePipe_valid; // @[BoxMuller.scala 103:25]
  wire [83:0] _io_g2_T_1 = $signed(sinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 104:15]
  reg  io_g2_v; // @[Valid.scala 127:22]
  reg [83:0] io_g2_b; // @[Reg.scala 16:16]
  wire [53:0] _GEN_42 = io_g1_b[83:30]; // @[BoxMuller.scala 98:9]
  wire [53:0] _GEN_44 = io_g2_b[83:30]; // @[BoxMuller.scala 102:9]
  wire [32:0] _GEN_46 = {$signed(trigonometric_io_theta_b), 1'h0}; // @[BoxMuller.scala 65:26]
  TauswortheUniform_12 rng1 ( // @[BoxMuller.scala 51:20]
    .clock(rng1_clock),
    .reset(rng1_reset),
    .io_rand_valid(rng1_io_rand_valid),
    .io_rand_bits(rng1_io_rand_bits)
  );
  TauswortheUniform_13 rng2 ( // @[BoxMuller.scala 52:20]
    .clock(rng2_clock),
    .reset(rng2_reset),
    .io_rand_valid(rng2_io_rand_valid),
    .io_rand_bits(rng2_io_rand_bits)
  );
  Trigonometric trigonometric ( // @[BoxMuller.scala 55:29]
    .clock(trigonometric_clock),
    .reset(trigonometric_reset),
    .io_theta_valid(trigonometric_io_theta_valid),
    .io_theta_bits(trigonometric_io_theta_bits),
    .io_result_valid(trigonometric_io_result_valid),
    .io_result_bits_sine(trigonometric_io_result_bits_sine),
    .io_result_bits_cosine(trigonometric_io_result_bits_cosine)
  );
  SquareRootLog sqrt_log ( // @[BoxMuller.scala 84:24]
    .clock(sqrt_log_clock),
    .reset(sqrt_log_reset),
    .io_uniform_valid(sqrt_log_io_uniform_valid),
    .io_uniform_bits(sqrt_log_io_uniform_bits),
    .io_result_valid(sqrt_log_io_result_valid),
    .io_result_bits(sqrt_log_io_result_bits)
  );
  assign io_g1_valid = io_g1_v; // @[Valid.scala 122:21 123:17]
  assign io_g1_bits = _GEN_42[51:0]; // @[BoxMuller.scala 98:9]
  assign io_g2_valid = io_g2_v; // @[Valid.scala 122:21 123:17]
  assign io_g2_bits = _GEN_44[51:0]; // @[BoxMuller.scala 102:9]
  assign rng1_clock = clock;
  assign rng1_reset = reset;
  assign rng2_clock = clock;
  assign rng2_reset = reset;
  assign trigonometric_clock = clock;
  assign trigonometric_reset = reset;
  assign trigonometric_io_theta_valid = trigonometric_io_theta_v; // @[Valid.scala 122:21 123:17]
  assign trigonometric_io_theta_bits = _GEN_46[31:0]; // @[BoxMuller.scala 65:26]
  assign sqrt_log_clock = clock;
  assign sqrt_log_reset = reset;
  assign sqrt_log_io_uniform_valid = sqrt_log_io_uniform_v; // @[Valid.scala 122:21 123:17]
  assign sqrt_log_io_uniform_bits = {{3{sqrt_log_io_uniform_b[28]}},sqrt_log_io_uniform_b}; // @[BoxMuller.scala 87:23]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits <= rng1_io_rand_bits[31:30]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_1 <= quadrantPipe_valid; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_1 <= quadrantPipe_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_2 <= quadrantPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_1) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_2 <= quadrantPipe_bits_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_3 <= quadrantPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_2) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_3 <= quadrantPipe_bits_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_4 <= quadrantPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_3) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_4 <= quadrantPipe_bits_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_5 <= quadrantPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_4) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_5 <= quadrantPipe_bits_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_6 <= quadrantPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_5) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_6 <= quadrantPipe_bits_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_7 <= quadrantPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_6) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_7 <= quadrantPipe_bits_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_8 <= quadrantPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_7) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_8 <= quadrantPipe_bits_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_9 <= quadrantPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_8) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_9 <= quadrantPipe_bits_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_10 <= quadrantPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_9) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_10 <= quadrantPipe_bits_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_11 <= quadrantPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_10) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_11 <= quadrantPipe_bits_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_12 <= quadrantPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_11) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_12 <= quadrantPipe_bits_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_13 <= quadrantPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_12) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_13 <= quadrantPipe_bits_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_14 <= quadrantPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_13) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_14 <= quadrantPipe_bits_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_15 <= quadrantPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_14) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_15 <= quadrantPipe_bits_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_16 <= quadrantPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_15) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_16 <= quadrantPipe_bits_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_17 <= quadrantPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_16) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_17 <= quadrantPipe_bits_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_18 <= quadrantPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_17) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_18 <= quadrantPipe_bits_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_19 <= quadrantPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_18) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_19 <= quadrantPipe_bits_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_20 <= quadrantPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_19) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_20 <= quadrantPipe_bits_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_21 <= quadrantPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_20) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_21 <= quadrantPipe_bits_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_22 <= quadrantPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_21) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_22 <= quadrantPipe_bits_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_23 <= quadrantPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_22) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_23 <= quadrantPipe_bits_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_24 <= quadrantPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_23) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_24 <= quadrantPipe_bits_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_25 <= quadrantPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_24) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_25 <= quadrantPipe_bits_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_26 <= quadrantPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_25) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_26 <= quadrantPipe_bits_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_27 <= quadrantPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_26) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_27 <= quadrantPipe_bits_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_28 <= quadrantPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_27) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_28 <= quadrantPipe_bits_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_29 <= quadrantPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_28) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_29 <= quadrantPipe_bits_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_30 <= quadrantPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_29) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_30 <= quadrantPipe_bits_29; // @[Reg.scala 17:22]
    end
    if (quadrantPipe_valid_30) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_31 <= quadrantPipe_bits_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      trigonometric_io_theta_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      trigonometric_io_theta_v <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      trigonometric_io_theta_b <= theta; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      cosinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      cosinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_cosine_T_2) begin // @[BoxMuller.scala 69:8]
        cosinePipe_bits <= trigonometric_io_result_bits_cosine;
      end else begin
        cosinePipe_bits <= _cosine_T_5;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      sinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_sine_T_2) begin // @[BoxMuller.scala 77:8]
        sinePipe_bits <= trigonometric_io_result_bits_sine;
      end else begin
        sinePipe_bits <= _sine_T_5;
      end
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      signPipe_bits <= rng2_io_rand_bits[31]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sqrt_log_io_uniform_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sqrt_log_io_uniform_v <= rng2_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      sqrt_log_io_uniform_b <= _sqrt_log_io_uniform_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sign_adjustedPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sign_adjustedPipe_valid <= sqrt_log_io_result_valid; // @[Valid.scala 127:22]
    end
    if (sqrt_log_io_result_valid) begin // @[Reg.scala 17:18]
      if (signPipe_bits) begin // @[BoxMuller.scala 91:8]
        sign_adjustedPipe_bits <= _sign_adjusted_T_3;
      end else begin
        sign_adjustedPipe_bits <= sqrt_log_io_result_bits;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g1_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g1_v <= _io_g1_T; // @[Valid.scala 127:22]
    end
    if (_io_g1_T) begin // @[Reg.scala 17:18]
      io_g1_b <= _io_g1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g2_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g2_v <= _io_g2_T; // @[Valid.scala 127:22]
    end
    if (_io_g2_T) begin // @[Reg.scala 17:18]
      io_g2_b <= _io_g2_T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quadrantPipe_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  quadrantPipe_bits = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  quadrantPipe_valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  quadrantPipe_bits_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  quadrantPipe_valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  quadrantPipe_bits_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  quadrantPipe_valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quadrantPipe_bits_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  quadrantPipe_valid_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  quadrantPipe_bits_4 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  quadrantPipe_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  quadrantPipe_bits_5 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  quadrantPipe_valid_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  quadrantPipe_bits_6 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  quadrantPipe_valid_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  quadrantPipe_bits_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  quadrantPipe_valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  quadrantPipe_bits_8 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  quadrantPipe_valid_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  quadrantPipe_bits_9 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  quadrantPipe_valid_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  quadrantPipe_bits_10 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  quadrantPipe_valid_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  quadrantPipe_bits_11 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  quadrantPipe_valid_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  quadrantPipe_bits_12 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  quadrantPipe_valid_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  quadrantPipe_bits_13 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  quadrantPipe_valid_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  quadrantPipe_bits_14 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  quadrantPipe_valid_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  quadrantPipe_bits_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  quadrantPipe_valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  quadrantPipe_bits_16 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  quadrantPipe_valid_17 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  quadrantPipe_bits_17 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  quadrantPipe_valid_18 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  quadrantPipe_bits_18 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  quadrantPipe_valid_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  quadrantPipe_bits_19 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  quadrantPipe_valid_20 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  quadrantPipe_bits_20 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  quadrantPipe_valid_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  quadrantPipe_bits_21 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  quadrantPipe_valid_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  quadrantPipe_bits_22 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  quadrantPipe_valid_23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  quadrantPipe_bits_23 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  quadrantPipe_valid_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  quadrantPipe_bits_24 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  quadrantPipe_valid_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  quadrantPipe_bits_25 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  quadrantPipe_valid_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  quadrantPipe_bits_26 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  quadrantPipe_valid_27 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  quadrantPipe_bits_27 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  quadrantPipe_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  quadrantPipe_bits_28 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  quadrantPipe_valid_29 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  quadrantPipe_bits_29 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  quadrantPipe_valid_30 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  quadrantPipe_bits_30 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  quadrantPipe_bits_31 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  trigonometric_io_theta_v = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  trigonometric_io_theta_b = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cosinePipe_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cosinePipe_bits = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sinePipe_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sinePipe_bits = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  signPipe_bits = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sqrt_log_io_uniform_v = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sqrt_log_io_uniform_b = _RAND_71[28:0];
  _RAND_72 = {1{`RANDOM}};
  sign_adjustedPipe_valid = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  sign_adjustedPipe_bits = _RAND_73[51:0];
  _RAND_74 = {1{`RANDOM}};
  io_g1_v = _RAND_74[0:0];
  _RAND_75 = {3{`RANDOM}};
  io_g1_b = _RAND_75[83:0];
  _RAND_76 = {1{`RANDOM}};
  io_g2_v = _RAND_76[0:0];
  _RAND_77 = {3{`RANDOM}};
  io_g2_b = _RAND_77[83:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MonteCarlo_6(
  input         clock,
  input         reset,
  output        io_request_0_ready,
  input         io_request_0_valid,
  input  [31:0] io_request_0_bits_time_steps,
  input  [31:0] io_request_0_bits_start_value,
  input  [31:0] io_request_0_bits_coefficient1,
  input  [31:0] io_request_0_bits_coefficient2,
  output        io_request_1_ready,
  input         io_request_1_valid,
  input  [31:0] io_request_1_bits_time_steps,
  input  [31:0] io_request_1_bits_start_value,
  input  [31:0] io_request_1_bits_coefficient1,
  input  [31:0] io_request_1_bits_coefficient2,
  input         io_response_0_ready,
  output        io_response_0_valid,
  output [31:0] io_response_0_bits,
  input         io_response_1_ready,
  output        io_response_1_valid,
  output [31:0] io_response_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rng_clock; // @[MonteCarlo.scala 42:19]
  wire  rng_reset; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g1_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g1_bits; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g2_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g2_bits; // @[MonteCarlo.scala 42:19]
  wire  initialized = rng_io_g1_valid & rng_io_g2_valid; // @[MonteCarlo.scala 47:37]
  reg [2:0] state; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_2 = $signed(io_request_0_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_3 = io_request_0_ready & io_request_0_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1; // @[Reg.scala 16:16]
  reg [31:0] c2; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_1 = io_request_0_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step; // @[Reg.scala 16:16]
  reg [31:0] price; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T = $signed(price) * $signed(c1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T = $signed(rng_io_g1_bits) * $signed(c2); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T = $signed(price) * $signed(partial_res2); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_2 = $signed(partial_res3) + $signed(partial_res1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_3 = counter == last_step ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_4 = counter == last_step ? counter : _counter_T_1; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_7 = io_response_0_ready & io_response_0_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_5 = _T_7 ? 3'h1 : state; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_6 = 3'h5 == state ? _GEN_5 : state; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_7 = 3'h4 == state ? $signed(_price_T_2) : $signed(price); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_3 : _GEN_6; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_9 = 3'h4 == state ? _GEN_4 : counter; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_64 = {$signed(partial_res3), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_10 = 3'h3 == state ? $signed(_partial_res3_T) : $signed({{12{_GEN_64[51]}},_GEN_64}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_11 = 3'h3 == state ? 3'h4 : _GEN_8; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_65 = {$signed(partial_res1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_14 = 3'h2 == state ? $signed(_partial_res1_T) : $signed({{12{_GEN_65[51]}},_GEN_65}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_66 = {$signed(partial_res2), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_15 = 3'h2 == state ? $signed(_partial_res2_T) : $signed({{20{_GEN_66[63]}},_GEN_66}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_17 = 3'h2 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_10); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_23 = 3'h1 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_14); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_24 = 3'h1 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_15); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_25 = 3'h1 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_17); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_29 = 3'h0 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_23); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_30 = 3'h0 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_24); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_31 = 3'h0 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_25); // @[MonteCarlo.scala 66:19 60:27]
  reg [2:0] state_1; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_6 = $signed(io_request_1_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_7 = io_request_1_ready & io_request_1_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1_1; // @[Reg.scala 16:16]
  reg [31:0] c2_1; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_4 = io_request_1_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step_1; // @[Reg.scala 16:16]
  reg [31:0] price_1; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1_1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2_1; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3_1; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter_1; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T_1 = $signed(price_1) * $signed(c1_1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T_1 = $signed(rng_io_g2_bits) * $signed(c2_1); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T_1 = $signed(price_1) * $signed(partial_res2_1); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_5 = $signed(partial_res3_1) + $signed(partial_res1_1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_35 = counter_1 == last_step_1 ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_36 = counter_1 == last_step_1 ? counter_1 : _counter_T_3; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_15 = io_response_1_ready & io_response_1_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_37 = _T_15 ? 3'h1 : state_1; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_38 = 3'h5 == state_1 ? _GEN_37 : state_1; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_39 = 3'h4 == state_1 ? $signed(_price_T_5) : $signed(price_1); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_40 = 3'h4 == state_1 ? _GEN_35 : _GEN_38; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_41 = 3'h4 == state_1 ? _GEN_36 : counter_1; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_74 = {$signed(partial_res3_1), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_42 = 3'h3 == state_1 ? $signed(_partial_res3_T_1) : $signed({{12{_GEN_74[51]}},_GEN_74}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_43 = 3'h3 == state_1 ? 3'h4 : _GEN_40; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_75 = {$signed(partial_res1_1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_46 = 3'h2 == state_1 ? $signed(_partial_res1_T_1) : $signed({{12{_GEN_75[51]}},_GEN_75}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_76 = {$signed(partial_res2_1), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_47 = 3'h2 == state_1 ? $signed(_partial_res2_T_1) : $signed({{20{_GEN_76[63]}},_GEN_76}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_49 = 3'h2 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_42); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_55 = 3'h1 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_46); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_56 = 3'h1 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_47); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_57 = 3'h1 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_49); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_61 = 3'h0 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_55); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_62 = 3'h0 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_56); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_63 = 3'h0 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_57); // @[MonteCarlo.scala 66:19 60:27]
  wire [43:0] _GEN_84 = _GEN_29[63:20];
  wire [51:0] _GEN_86 = _GEN_30[83:32];
  wire [43:0] _GEN_88 = _GEN_31[63:20];
  wire [43:0] _GEN_90 = _GEN_61[63:20];
  wire [51:0] _GEN_92 = _GEN_62[83:32];
  wire [43:0] _GEN_94 = _GEN_63[63:20];
  BoxMuller_6 rng ( // @[MonteCarlo.scala 42:19]
    .clock(rng_clock),
    .reset(rng_reset),
    .io_g1_valid(rng_io_g1_valid),
    .io_g1_bits(rng_io_g1_bits),
    .io_g2_valid(rng_io_g2_valid),
    .io_g2_bits(rng_io_g2_bits)
  );
  assign io_request_0_ready = state == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_request_1_ready = state_1 == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_response_0_valid = state == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_0_bits = price; // @[MonteCarlo.scala 65:16]
  assign io_response_1_valid = state_1 == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_1_bits = price_1; // @[MonteCarlo.scala 65:16]
  assign rng_clock = clock;
  assign rng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state <= 3'h1;
      end else begin
        state <= 3'h0;
      end
    end else if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_3) begin // @[MonteCarlo.scala 71:23]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[MonteCarlo.scala 66:19]
      state <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state <= _GEN_11;
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c1 <= _c1_T_2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c2 <= io_request_0_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      last_step <= _last_step_T_1; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        price <= io_request_0_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          price <= _GEN_7;
        end
      end
    end
    partial_res1 <= _GEN_84[31:0];
    partial_res2 <= _GEN_86[31:0];
    partial_res3 <= _GEN_88[31:0];
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        counter <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          counter <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state_1 <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state_1 <= 3'h1;
      end else begin
        state_1 <= 3'h0;
      end
    end else if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_7) begin // @[MonteCarlo.scala 71:23]
        state_1 <= 3'h2;
      end else begin
        state_1 <= 3'h1;
      end
    end else if (3'h2 == state_1) begin // @[MonteCarlo.scala 66:19]
      state_1 <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state_1 <= _GEN_43;
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c1_1 <= _c1_T_6; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c2_1 <= io_request_1_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      last_step_1 <= _last_step_T_4; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        price_1 <= io_request_1_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          price_1 <= _GEN_39;
        end
      end
    end
    partial_res1_1 <= _GEN_90[31:0];
    partial_res2_1 <= _GEN_92[31:0];
    partial_res3_1 <= _GEN_94[31:0];
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        counter_1 <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          counter_1 <= _GEN_41;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  c1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_step = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  price = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  partial_res1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  partial_res2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  partial_res3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  c1_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_step_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  price_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  partial_res1_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  partial_res2_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  partial_res3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  counter_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_14(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h1f2ed2a5 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h37880c11 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h2fc26b47 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_15(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h3ec7ce35 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h2eebf6a5 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h247b7124 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoxMuller_7(
  input         clock,
  input         reset,
  output        io_g1_valid,
  output [51:0] io_g1_bits,
  output        io_g2_valid,
  output [51:0] io_g2_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [95:0] _RAND_77;
`endif // RANDOMIZE_REG_INIT
  wire  rng1_clock; // @[BoxMuller.scala 51:20]
  wire  rng1_reset; // @[BoxMuller.scala 51:20]
  wire  rng1_io_rand_valid; // @[BoxMuller.scala 51:20]
  wire [31:0] rng1_io_rand_bits; // @[BoxMuller.scala 51:20]
  wire  rng2_clock; // @[BoxMuller.scala 52:20]
  wire  rng2_reset; // @[BoxMuller.scala 52:20]
  wire  rng2_io_rand_valid; // @[BoxMuller.scala 52:20]
  wire [31:0] rng2_io_rand_bits; // @[BoxMuller.scala 52:20]
  wire  trigonometric_clock; // @[BoxMuller.scala 55:29]
  wire  trigonometric_reset; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_theta_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_theta_bits; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_result_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_sine; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_cosine; // @[BoxMuller.scala 55:29]
  wire  sqrt_log_clock; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_reset; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_uniform_valid; // @[BoxMuller.scala 84:24]
  wire [31:0] sqrt_log_io_uniform_bits; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_result_valid; // @[BoxMuller.scala 84:24]
  wire [51:0] sqrt_log_io_result_bits; // @[BoxMuller.scala 84:24]
  wire [30:0] _theta_T_3 = {2'h0,rng1_io_rand_bits[28:0]}; // @[BoxMuller.scala 62:18]
  wire [62:0] _theta_T_4 = $signed(_theta_T_3) * 32'sh6487ed51; // @[BoxMuller.scala 62:26]
  reg  quadrantPipe_valid; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_1; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_1; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_2; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_2; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_3; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_3; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_4; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_4; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_5; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_5; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_6; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_6; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_7; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_7; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_8; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_8; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_9; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_9; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_10; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_10; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_11; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_11; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_12; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_12; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_13; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_13; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_14; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_14; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_15; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_15; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_16; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_16; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_17; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_17; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_18; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_18; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_19; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_19; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_20; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_20; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_21; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_21; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_22; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_22; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_23; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_23; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_24; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_24; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_25; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_25; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_26; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_26; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_27; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_27; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_28; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_28; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_29; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_29; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_30; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_30; // @[Reg.scala 16:16]
  reg [1:0] quadrantPipe_bits_31; // @[Reg.scala 16:16]
  reg  trigonometric_io_theta_v; // @[Valid.scala 127:22]
  reg [31:0] trigonometric_io_theta_b; // @[Reg.scala 16:16]
  wire [33:0] _GEN_40 = _theta_T_4[62:29]; // @[BoxMuller.scala 59:19 61:9]
  wire [31:0] theta = _GEN_40[31:0]; // @[BoxMuller.scala 59:19 61:9]
  wire  _cosine_T = quadrantPipe_bits_31 == 2'h0; // @[BoxMuller.scala 70:21]
  wire  _cosine_T_2 = quadrantPipe_bits_31 == 2'h0 | quadrantPipe_bits_31 == 2'h3; // @[BoxMuller.scala 70:29]
  wire [31:0] _cosine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_cosine); // @[BoxMuller.scala 72:7]
  reg  cosinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] cosinePipe_bits; // @[Reg.scala 16:16]
  wire  _sine_T_2 = _cosine_T | quadrantPipe_bits_31 == 2'h2; // @[BoxMuller.scala 78:29]
  wire [31:0] _sine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_sine); // @[BoxMuller.scala 80:7]
  reg  sinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] sinePipe_bits; // @[Reg.scala 16:16]
  reg  signPipe_bits; // @[Reg.scala 16:16]
  wire [28:0] _sqrt_log_io_uniform_T_1 = rng2_io_rand_bits[28:0]; // @[BoxMuller.scala 87:89]
  reg  sqrt_log_io_uniform_v; // @[Valid.scala 127:22]
  reg [28:0] sqrt_log_io_uniform_b; // @[Reg.scala 16:16]
  wire [51:0] _sign_adjusted_T_3 = 52'sh0 - $signed(sqrt_log_io_result_bits); // @[BoxMuller.scala 93:7]
  reg  sign_adjustedPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] sign_adjustedPipe_bits; // @[Reg.scala 16:16]
  wire  _io_g1_T = sign_adjustedPipe_valid & cosinePipe_valid; // @[BoxMuller.scala 99:25]
  wire [83:0] _io_g1_T_1 = $signed(cosinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 100:17]
  reg  io_g1_v; // @[Valid.scala 127:22]
  reg [83:0] io_g1_b; // @[Reg.scala 16:16]
  wire  _io_g2_T = sign_adjustedPipe_valid & sinePipe_valid; // @[BoxMuller.scala 103:25]
  wire [83:0] _io_g2_T_1 = $signed(sinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 104:15]
  reg  io_g2_v; // @[Valid.scala 127:22]
  reg [83:0] io_g2_b; // @[Reg.scala 16:16]
  wire [53:0] _GEN_42 = io_g1_b[83:30]; // @[BoxMuller.scala 98:9]
  wire [53:0] _GEN_44 = io_g2_b[83:30]; // @[BoxMuller.scala 102:9]
  wire [32:0] _GEN_46 = {$signed(trigonometric_io_theta_b), 1'h0}; // @[BoxMuller.scala 65:26]
  TauswortheUniform_14 rng1 ( // @[BoxMuller.scala 51:20]
    .clock(rng1_clock),
    .reset(rng1_reset),
    .io_rand_valid(rng1_io_rand_valid),
    .io_rand_bits(rng1_io_rand_bits)
  );
  TauswortheUniform_15 rng2 ( // @[BoxMuller.scala 52:20]
    .clock(rng2_clock),
    .reset(rng2_reset),
    .io_rand_valid(rng2_io_rand_valid),
    .io_rand_bits(rng2_io_rand_bits)
  );
  Trigonometric trigonometric ( // @[BoxMuller.scala 55:29]
    .clock(trigonometric_clock),
    .reset(trigonometric_reset),
    .io_theta_valid(trigonometric_io_theta_valid),
    .io_theta_bits(trigonometric_io_theta_bits),
    .io_result_valid(trigonometric_io_result_valid),
    .io_result_bits_sine(trigonometric_io_result_bits_sine),
    .io_result_bits_cosine(trigonometric_io_result_bits_cosine)
  );
  SquareRootLog sqrt_log ( // @[BoxMuller.scala 84:24]
    .clock(sqrt_log_clock),
    .reset(sqrt_log_reset),
    .io_uniform_valid(sqrt_log_io_uniform_valid),
    .io_uniform_bits(sqrt_log_io_uniform_bits),
    .io_result_valid(sqrt_log_io_result_valid),
    .io_result_bits(sqrt_log_io_result_bits)
  );
  assign io_g1_valid = io_g1_v; // @[Valid.scala 122:21 123:17]
  assign io_g1_bits = _GEN_42[51:0]; // @[BoxMuller.scala 98:9]
  assign io_g2_valid = io_g2_v; // @[Valid.scala 122:21 123:17]
  assign io_g2_bits = _GEN_44[51:0]; // @[BoxMuller.scala 102:9]
  assign rng1_clock = clock;
  assign rng1_reset = reset;
  assign rng2_clock = clock;
  assign rng2_reset = reset;
  assign trigonometric_clock = clock;
  assign trigonometric_reset = reset;
  assign trigonometric_io_theta_valid = trigonometric_io_theta_v; // @[Valid.scala 122:21 123:17]
  assign trigonometric_io_theta_bits = _GEN_46[31:0]; // @[BoxMuller.scala 65:26]
  assign sqrt_log_clock = clock;
  assign sqrt_log_reset = reset;
  assign sqrt_log_io_uniform_valid = sqrt_log_io_uniform_v; // @[Valid.scala 122:21 123:17]
  assign sqrt_log_io_uniform_bits = {{3{sqrt_log_io_uniform_b[28]}},sqrt_log_io_uniform_b}; // @[BoxMuller.scala 87:23]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits <= rng1_io_rand_bits[31:30]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_1 <= quadrantPipe_valid; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_1 <= quadrantPipe_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_2 <= quadrantPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_1) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_2 <= quadrantPipe_bits_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_3 <= quadrantPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_2) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_3 <= quadrantPipe_bits_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_4 <= quadrantPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_3) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_4 <= quadrantPipe_bits_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_5 <= quadrantPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_4) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_5 <= quadrantPipe_bits_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_6 <= quadrantPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_5) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_6 <= quadrantPipe_bits_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_7 <= quadrantPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_6) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_7 <= quadrantPipe_bits_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_8 <= quadrantPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_7) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_8 <= quadrantPipe_bits_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_9 <= quadrantPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_8) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_9 <= quadrantPipe_bits_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_10 <= quadrantPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_9) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_10 <= quadrantPipe_bits_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_11 <= quadrantPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_10) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_11 <= quadrantPipe_bits_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_12 <= quadrantPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_11) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_12 <= quadrantPipe_bits_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_13 <= quadrantPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_12) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_13 <= quadrantPipe_bits_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_14 <= quadrantPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_13) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_14 <= quadrantPipe_bits_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_15 <= quadrantPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_14) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_15 <= quadrantPipe_bits_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_16 <= quadrantPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_15) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_16 <= quadrantPipe_bits_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_17 <= quadrantPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_16) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_17 <= quadrantPipe_bits_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_18 <= quadrantPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_17) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_18 <= quadrantPipe_bits_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_19 <= quadrantPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_18) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_19 <= quadrantPipe_bits_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_20 <= quadrantPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_19) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_20 <= quadrantPipe_bits_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_21 <= quadrantPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_20) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_21 <= quadrantPipe_bits_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_22 <= quadrantPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_21) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_22 <= quadrantPipe_bits_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_23 <= quadrantPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_22) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_23 <= quadrantPipe_bits_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_24 <= quadrantPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_23) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_24 <= quadrantPipe_bits_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_25 <= quadrantPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_24) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_25 <= quadrantPipe_bits_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_26 <= quadrantPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_25) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_26 <= quadrantPipe_bits_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_27 <= quadrantPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_26) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_27 <= quadrantPipe_bits_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_28 <= quadrantPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_27) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_28 <= quadrantPipe_bits_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_29 <= quadrantPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_28) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_29 <= quadrantPipe_bits_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_30 <= quadrantPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_29) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_30 <= quadrantPipe_bits_29; // @[Reg.scala 17:22]
    end
    if (quadrantPipe_valid_30) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_31 <= quadrantPipe_bits_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      trigonometric_io_theta_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      trigonometric_io_theta_v <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      trigonometric_io_theta_b <= theta; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      cosinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      cosinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_cosine_T_2) begin // @[BoxMuller.scala 69:8]
        cosinePipe_bits <= trigonometric_io_result_bits_cosine;
      end else begin
        cosinePipe_bits <= _cosine_T_5;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      sinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_sine_T_2) begin // @[BoxMuller.scala 77:8]
        sinePipe_bits <= trigonometric_io_result_bits_sine;
      end else begin
        sinePipe_bits <= _sine_T_5;
      end
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      signPipe_bits <= rng2_io_rand_bits[31]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sqrt_log_io_uniform_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sqrt_log_io_uniform_v <= rng2_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      sqrt_log_io_uniform_b <= _sqrt_log_io_uniform_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sign_adjustedPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sign_adjustedPipe_valid <= sqrt_log_io_result_valid; // @[Valid.scala 127:22]
    end
    if (sqrt_log_io_result_valid) begin // @[Reg.scala 17:18]
      if (signPipe_bits) begin // @[BoxMuller.scala 91:8]
        sign_adjustedPipe_bits <= _sign_adjusted_T_3;
      end else begin
        sign_adjustedPipe_bits <= sqrt_log_io_result_bits;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g1_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g1_v <= _io_g1_T; // @[Valid.scala 127:22]
    end
    if (_io_g1_T) begin // @[Reg.scala 17:18]
      io_g1_b <= _io_g1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g2_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g2_v <= _io_g2_T; // @[Valid.scala 127:22]
    end
    if (_io_g2_T) begin // @[Reg.scala 17:18]
      io_g2_b <= _io_g2_T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quadrantPipe_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  quadrantPipe_bits = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  quadrantPipe_valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  quadrantPipe_bits_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  quadrantPipe_valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  quadrantPipe_bits_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  quadrantPipe_valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quadrantPipe_bits_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  quadrantPipe_valid_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  quadrantPipe_bits_4 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  quadrantPipe_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  quadrantPipe_bits_5 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  quadrantPipe_valid_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  quadrantPipe_bits_6 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  quadrantPipe_valid_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  quadrantPipe_bits_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  quadrantPipe_valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  quadrantPipe_bits_8 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  quadrantPipe_valid_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  quadrantPipe_bits_9 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  quadrantPipe_valid_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  quadrantPipe_bits_10 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  quadrantPipe_valid_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  quadrantPipe_bits_11 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  quadrantPipe_valid_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  quadrantPipe_bits_12 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  quadrantPipe_valid_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  quadrantPipe_bits_13 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  quadrantPipe_valid_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  quadrantPipe_bits_14 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  quadrantPipe_valid_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  quadrantPipe_bits_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  quadrantPipe_valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  quadrantPipe_bits_16 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  quadrantPipe_valid_17 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  quadrantPipe_bits_17 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  quadrantPipe_valid_18 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  quadrantPipe_bits_18 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  quadrantPipe_valid_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  quadrantPipe_bits_19 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  quadrantPipe_valid_20 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  quadrantPipe_bits_20 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  quadrantPipe_valid_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  quadrantPipe_bits_21 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  quadrantPipe_valid_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  quadrantPipe_bits_22 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  quadrantPipe_valid_23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  quadrantPipe_bits_23 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  quadrantPipe_valid_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  quadrantPipe_bits_24 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  quadrantPipe_valid_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  quadrantPipe_bits_25 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  quadrantPipe_valid_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  quadrantPipe_bits_26 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  quadrantPipe_valid_27 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  quadrantPipe_bits_27 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  quadrantPipe_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  quadrantPipe_bits_28 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  quadrantPipe_valid_29 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  quadrantPipe_bits_29 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  quadrantPipe_valid_30 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  quadrantPipe_bits_30 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  quadrantPipe_bits_31 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  trigonometric_io_theta_v = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  trigonometric_io_theta_b = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cosinePipe_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cosinePipe_bits = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sinePipe_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sinePipe_bits = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  signPipe_bits = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sqrt_log_io_uniform_v = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sqrt_log_io_uniform_b = _RAND_71[28:0];
  _RAND_72 = {1{`RANDOM}};
  sign_adjustedPipe_valid = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  sign_adjustedPipe_bits = _RAND_73[51:0];
  _RAND_74 = {1{`RANDOM}};
  io_g1_v = _RAND_74[0:0];
  _RAND_75 = {3{`RANDOM}};
  io_g1_b = _RAND_75[83:0];
  _RAND_76 = {1{`RANDOM}};
  io_g2_v = _RAND_76[0:0];
  _RAND_77 = {3{`RANDOM}};
  io_g2_b = _RAND_77[83:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MonteCarlo_7(
  input         clock,
  input         reset,
  output        io_request_0_ready,
  input         io_request_0_valid,
  input  [31:0] io_request_0_bits_time_steps,
  input  [31:0] io_request_0_bits_start_value,
  input  [31:0] io_request_0_bits_coefficient1,
  input  [31:0] io_request_0_bits_coefficient2,
  output        io_request_1_ready,
  input         io_request_1_valid,
  input  [31:0] io_request_1_bits_time_steps,
  input  [31:0] io_request_1_bits_start_value,
  input  [31:0] io_request_1_bits_coefficient1,
  input  [31:0] io_request_1_bits_coefficient2,
  input         io_response_0_ready,
  output        io_response_0_valid,
  output [31:0] io_response_0_bits,
  input         io_response_1_ready,
  output        io_response_1_valid,
  output [31:0] io_response_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rng_clock; // @[MonteCarlo.scala 42:19]
  wire  rng_reset; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g1_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g1_bits; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g2_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g2_bits; // @[MonteCarlo.scala 42:19]
  wire  initialized = rng_io_g1_valid & rng_io_g2_valid; // @[MonteCarlo.scala 47:37]
  reg [2:0] state; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_2 = $signed(io_request_0_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_3 = io_request_0_ready & io_request_0_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1; // @[Reg.scala 16:16]
  reg [31:0] c2; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_1 = io_request_0_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step; // @[Reg.scala 16:16]
  reg [31:0] price; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T = $signed(price) * $signed(c1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T = $signed(rng_io_g1_bits) * $signed(c2); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T = $signed(price) * $signed(partial_res2); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_2 = $signed(partial_res3) + $signed(partial_res1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_3 = counter == last_step ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_4 = counter == last_step ? counter : _counter_T_1; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_7 = io_response_0_ready & io_response_0_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_5 = _T_7 ? 3'h1 : state; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_6 = 3'h5 == state ? _GEN_5 : state; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_7 = 3'h4 == state ? $signed(_price_T_2) : $signed(price); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_3 : _GEN_6; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_9 = 3'h4 == state ? _GEN_4 : counter; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_64 = {$signed(partial_res3), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_10 = 3'h3 == state ? $signed(_partial_res3_T) : $signed({{12{_GEN_64[51]}},_GEN_64}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_11 = 3'h3 == state ? 3'h4 : _GEN_8; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_65 = {$signed(partial_res1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_14 = 3'h2 == state ? $signed(_partial_res1_T) : $signed({{12{_GEN_65[51]}},_GEN_65}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_66 = {$signed(partial_res2), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_15 = 3'h2 == state ? $signed(_partial_res2_T) : $signed({{20{_GEN_66[63]}},_GEN_66}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_17 = 3'h2 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_10); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_23 = 3'h1 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_14); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_24 = 3'h1 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_15); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_25 = 3'h1 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_17); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_29 = 3'h0 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_23); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_30 = 3'h0 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_24); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_31 = 3'h0 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_25); // @[MonteCarlo.scala 66:19 60:27]
  reg [2:0] state_1; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_6 = $signed(io_request_1_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_7 = io_request_1_ready & io_request_1_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1_1; // @[Reg.scala 16:16]
  reg [31:0] c2_1; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_4 = io_request_1_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step_1; // @[Reg.scala 16:16]
  reg [31:0] price_1; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1_1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2_1; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3_1; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter_1; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T_1 = $signed(price_1) * $signed(c1_1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T_1 = $signed(rng_io_g2_bits) * $signed(c2_1); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T_1 = $signed(price_1) * $signed(partial_res2_1); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_5 = $signed(partial_res3_1) + $signed(partial_res1_1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_35 = counter_1 == last_step_1 ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_36 = counter_1 == last_step_1 ? counter_1 : _counter_T_3; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_15 = io_response_1_ready & io_response_1_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_37 = _T_15 ? 3'h1 : state_1; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_38 = 3'h5 == state_1 ? _GEN_37 : state_1; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_39 = 3'h4 == state_1 ? $signed(_price_T_5) : $signed(price_1); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_40 = 3'h4 == state_1 ? _GEN_35 : _GEN_38; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_41 = 3'h4 == state_1 ? _GEN_36 : counter_1; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_74 = {$signed(partial_res3_1), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_42 = 3'h3 == state_1 ? $signed(_partial_res3_T_1) : $signed({{12{_GEN_74[51]}},_GEN_74}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_43 = 3'h3 == state_1 ? 3'h4 : _GEN_40; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_75 = {$signed(partial_res1_1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_46 = 3'h2 == state_1 ? $signed(_partial_res1_T_1) : $signed({{12{_GEN_75[51]}},_GEN_75}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_76 = {$signed(partial_res2_1), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_47 = 3'h2 == state_1 ? $signed(_partial_res2_T_1) : $signed({{20{_GEN_76[63]}},_GEN_76}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_49 = 3'h2 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_42); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_55 = 3'h1 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_46); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_56 = 3'h1 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_47); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_57 = 3'h1 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_49); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_61 = 3'h0 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_55); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_62 = 3'h0 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_56); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_63 = 3'h0 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_57); // @[MonteCarlo.scala 66:19 60:27]
  wire [43:0] _GEN_84 = _GEN_29[63:20];
  wire [51:0] _GEN_86 = _GEN_30[83:32];
  wire [43:0] _GEN_88 = _GEN_31[63:20];
  wire [43:0] _GEN_90 = _GEN_61[63:20];
  wire [51:0] _GEN_92 = _GEN_62[83:32];
  wire [43:0] _GEN_94 = _GEN_63[63:20];
  BoxMuller_7 rng ( // @[MonteCarlo.scala 42:19]
    .clock(rng_clock),
    .reset(rng_reset),
    .io_g1_valid(rng_io_g1_valid),
    .io_g1_bits(rng_io_g1_bits),
    .io_g2_valid(rng_io_g2_valid),
    .io_g2_bits(rng_io_g2_bits)
  );
  assign io_request_0_ready = state == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_request_1_ready = state_1 == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_response_0_valid = state == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_0_bits = price; // @[MonteCarlo.scala 65:16]
  assign io_response_1_valid = state_1 == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_1_bits = price_1; // @[MonteCarlo.scala 65:16]
  assign rng_clock = clock;
  assign rng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state <= 3'h1;
      end else begin
        state <= 3'h0;
      end
    end else if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_3) begin // @[MonteCarlo.scala 71:23]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[MonteCarlo.scala 66:19]
      state <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state <= _GEN_11;
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c1 <= _c1_T_2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c2 <= io_request_0_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      last_step <= _last_step_T_1; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        price <= io_request_0_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          price <= _GEN_7;
        end
      end
    end
    partial_res1 <= _GEN_84[31:0];
    partial_res2 <= _GEN_86[31:0];
    partial_res3 <= _GEN_88[31:0];
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        counter <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          counter <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state_1 <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state_1 <= 3'h1;
      end else begin
        state_1 <= 3'h0;
      end
    end else if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_7) begin // @[MonteCarlo.scala 71:23]
        state_1 <= 3'h2;
      end else begin
        state_1 <= 3'h1;
      end
    end else if (3'h2 == state_1) begin // @[MonteCarlo.scala 66:19]
      state_1 <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state_1 <= _GEN_43;
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c1_1 <= _c1_T_6; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c2_1 <= io_request_1_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      last_step_1 <= _last_step_T_4; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        price_1 <= io_request_1_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          price_1 <= _GEN_39;
        end
      end
    end
    partial_res1_1 <= _GEN_90[31:0];
    partial_res2_1 <= _GEN_92[31:0];
    partial_res3_1 <= _GEN_94[31:0];
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        counter_1 <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          counter_1 <= _GEN_41;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  c1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_step = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  price = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  partial_res1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  partial_res2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  partial_res3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  c1_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_step_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  price_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  partial_res1_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  partial_res2_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  partial_res3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  counter_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_16(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h344e9868 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'hd1d2f7 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h35b0612b : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_17(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h1a61c68e : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h21b57188 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h2e731867 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoxMuller_8(
  input         clock,
  input         reset,
  output        io_g1_valid,
  output [51:0] io_g1_bits,
  output        io_g2_valid,
  output [51:0] io_g2_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [95:0] _RAND_77;
`endif // RANDOMIZE_REG_INIT
  wire  rng1_clock; // @[BoxMuller.scala 51:20]
  wire  rng1_reset; // @[BoxMuller.scala 51:20]
  wire  rng1_io_rand_valid; // @[BoxMuller.scala 51:20]
  wire [31:0] rng1_io_rand_bits; // @[BoxMuller.scala 51:20]
  wire  rng2_clock; // @[BoxMuller.scala 52:20]
  wire  rng2_reset; // @[BoxMuller.scala 52:20]
  wire  rng2_io_rand_valid; // @[BoxMuller.scala 52:20]
  wire [31:0] rng2_io_rand_bits; // @[BoxMuller.scala 52:20]
  wire  trigonometric_clock; // @[BoxMuller.scala 55:29]
  wire  trigonometric_reset; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_theta_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_theta_bits; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_result_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_sine; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_cosine; // @[BoxMuller.scala 55:29]
  wire  sqrt_log_clock; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_reset; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_uniform_valid; // @[BoxMuller.scala 84:24]
  wire [31:0] sqrt_log_io_uniform_bits; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_result_valid; // @[BoxMuller.scala 84:24]
  wire [51:0] sqrt_log_io_result_bits; // @[BoxMuller.scala 84:24]
  wire [30:0] _theta_T_3 = {2'h0,rng1_io_rand_bits[28:0]}; // @[BoxMuller.scala 62:18]
  wire [62:0] _theta_T_4 = $signed(_theta_T_3) * 32'sh6487ed51; // @[BoxMuller.scala 62:26]
  reg  quadrantPipe_valid; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_1; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_1; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_2; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_2; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_3; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_3; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_4; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_4; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_5; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_5; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_6; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_6; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_7; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_7; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_8; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_8; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_9; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_9; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_10; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_10; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_11; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_11; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_12; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_12; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_13; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_13; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_14; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_14; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_15; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_15; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_16; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_16; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_17; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_17; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_18; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_18; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_19; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_19; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_20; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_20; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_21; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_21; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_22; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_22; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_23; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_23; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_24; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_24; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_25; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_25; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_26; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_26; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_27; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_27; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_28; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_28; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_29; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_29; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_30; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_30; // @[Reg.scala 16:16]
  reg [1:0] quadrantPipe_bits_31; // @[Reg.scala 16:16]
  reg  trigonometric_io_theta_v; // @[Valid.scala 127:22]
  reg [31:0] trigonometric_io_theta_b; // @[Reg.scala 16:16]
  wire [33:0] _GEN_40 = _theta_T_4[62:29]; // @[BoxMuller.scala 59:19 61:9]
  wire [31:0] theta = _GEN_40[31:0]; // @[BoxMuller.scala 59:19 61:9]
  wire  _cosine_T = quadrantPipe_bits_31 == 2'h0; // @[BoxMuller.scala 70:21]
  wire  _cosine_T_2 = quadrantPipe_bits_31 == 2'h0 | quadrantPipe_bits_31 == 2'h3; // @[BoxMuller.scala 70:29]
  wire [31:0] _cosine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_cosine); // @[BoxMuller.scala 72:7]
  reg  cosinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] cosinePipe_bits; // @[Reg.scala 16:16]
  wire  _sine_T_2 = _cosine_T | quadrantPipe_bits_31 == 2'h2; // @[BoxMuller.scala 78:29]
  wire [31:0] _sine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_sine); // @[BoxMuller.scala 80:7]
  reg  sinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] sinePipe_bits; // @[Reg.scala 16:16]
  reg  signPipe_bits; // @[Reg.scala 16:16]
  wire [28:0] _sqrt_log_io_uniform_T_1 = rng2_io_rand_bits[28:0]; // @[BoxMuller.scala 87:89]
  reg  sqrt_log_io_uniform_v; // @[Valid.scala 127:22]
  reg [28:0] sqrt_log_io_uniform_b; // @[Reg.scala 16:16]
  wire [51:0] _sign_adjusted_T_3 = 52'sh0 - $signed(sqrt_log_io_result_bits); // @[BoxMuller.scala 93:7]
  reg  sign_adjustedPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] sign_adjustedPipe_bits; // @[Reg.scala 16:16]
  wire  _io_g1_T = sign_adjustedPipe_valid & cosinePipe_valid; // @[BoxMuller.scala 99:25]
  wire [83:0] _io_g1_T_1 = $signed(cosinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 100:17]
  reg  io_g1_v; // @[Valid.scala 127:22]
  reg [83:0] io_g1_b; // @[Reg.scala 16:16]
  wire  _io_g2_T = sign_adjustedPipe_valid & sinePipe_valid; // @[BoxMuller.scala 103:25]
  wire [83:0] _io_g2_T_1 = $signed(sinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 104:15]
  reg  io_g2_v; // @[Valid.scala 127:22]
  reg [83:0] io_g2_b; // @[Reg.scala 16:16]
  wire [53:0] _GEN_42 = io_g1_b[83:30]; // @[BoxMuller.scala 98:9]
  wire [53:0] _GEN_44 = io_g2_b[83:30]; // @[BoxMuller.scala 102:9]
  wire [32:0] _GEN_46 = {$signed(trigonometric_io_theta_b), 1'h0}; // @[BoxMuller.scala 65:26]
  TauswortheUniform_16 rng1 ( // @[BoxMuller.scala 51:20]
    .clock(rng1_clock),
    .reset(rng1_reset),
    .io_rand_valid(rng1_io_rand_valid),
    .io_rand_bits(rng1_io_rand_bits)
  );
  TauswortheUniform_17 rng2 ( // @[BoxMuller.scala 52:20]
    .clock(rng2_clock),
    .reset(rng2_reset),
    .io_rand_valid(rng2_io_rand_valid),
    .io_rand_bits(rng2_io_rand_bits)
  );
  Trigonometric trigonometric ( // @[BoxMuller.scala 55:29]
    .clock(trigonometric_clock),
    .reset(trigonometric_reset),
    .io_theta_valid(trigonometric_io_theta_valid),
    .io_theta_bits(trigonometric_io_theta_bits),
    .io_result_valid(trigonometric_io_result_valid),
    .io_result_bits_sine(trigonometric_io_result_bits_sine),
    .io_result_bits_cosine(trigonometric_io_result_bits_cosine)
  );
  SquareRootLog sqrt_log ( // @[BoxMuller.scala 84:24]
    .clock(sqrt_log_clock),
    .reset(sqrt_log_reset),
    .io_uniform_valid(sqrt_log_io_uniform_valid),
    .io_uniform_bits(sqrt_log_io_uniform_bits),
    .io_result_valid(sqrt_log_io_result_valid),
    .io_result_bits(sqrt_log_io_result_bits)
  );
  assign io_g1_valid = io_g1_v; // @[Valid.scala 122:21 123:17]
  assign io_g1_bits = _GEN_42[51:0]; // @[BoxMuller.scala 98:9]
  assign io_g2_valid = io_g2_v; // @[Valid.scala 122:21 123:17]
  assign io_g2_bits = _GEN_44[51:0]; // @[BoxMuller.scala 102:9]
  assign rng1_clock = clock;
  assign rng1_reset = reset;
  assign rng2_clock = clock;
  assign rng2_reset = reset;
  assign trigonometric_clock = clock;
  assign trigonometric_reset = reset;
  assign trigonometric_io_theta_valid = trigonometric_io_theta_v; // @[Valid.scala 122:21 123:17]
  assign trigonometric_io_theta_bits = _GEN_46[31:0]; // @[BoxMuller.scala 65:26]
  assign sqrt_log_clock = clock;
  assign sqrt_log_reset = reset;
  assign sqrt_log_io_uniform_valid = sqrt_log_io_uniform_v; // @[Valid.scala 122:21 123:17]
  assign sqrt_log_io_uniform_bits = {{3{sqrt_log_io_uniform_b[28]}},sqrt_log_io_uniform_b}; // @[BoxMuller.scala 87:23]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits <= rng1_io_rand_bits[31:30]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_1 <= quadrantPipe_valid; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_1 <= quadrantPipe_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_2 <= quadrantPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_1) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_2 <= quadrantPipe_bits_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_3 <= quadrantPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_2) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_3 <= quadrantPipe_bits_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_4 <= quadrantPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_3) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_4 <= quadrantPipe_bits_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_5 <= quadrantPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_4) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_5 <= quadrantPipe_bits_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_6 <= quadrantPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_5) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_6 <= quadrantPipe_bits_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_7 <= quadrantPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_6) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_7 <= quadrantPipe_bits_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_8 <= quadrantPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_7) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_8 <= quadrantPipe_bits_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_9 <= quadrantPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_8) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_9 <= quadrantPipe_bits_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_10 <= quadrantPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_9) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_10 <= quadrantPipe_bits_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_11 <= quadrantPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_10) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_11 <= quadrantPipe_bits_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_12 <= quadrantPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_11) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_12 <= quadrantPipe_bits_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_13 <= quadrantPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_12) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_13 <= quadrantPipe_bits_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_14 <= quadrantPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_13) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_14 <= quadrantPipe_bits_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_15 <= quadrantPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_14) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_15 <= quadrantPipe_bits_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_16 <= quadrantPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_15) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_16 <= quadrantPipe_bits_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_17 <= quadrantPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_16) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_17 <= quadrantPipe_bits_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_18 <= quadrantPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_17) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_18 <= quadrantPipe_bits_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_19 <= quadrantPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_18) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_19 <= quadrantPipe_bits_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_20 <= quadrantPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_19) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_20 <= quadrantPipe_bits_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_21 <= quadrantPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_20) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_21 <= quadrantPipe_bits_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_22 <= quadrantPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_21) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_22 <= quadrantPipe_bits_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_23 <= quadrantPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_22) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_23 <= quadrantPipe_bits_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_24 <= quadrantPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_23) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_24 <= quadrantPipe_bits_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_25 <= quadrantPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_24) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_25 <= quadrantPipe_bits_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_26 <= quadrantPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_25) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_26 <= quadrantPipe_bits_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_27 <= quadrantPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_26) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_27 <= quadrantPipe_bits_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_28 <= quadrantPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_27) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_28 <= quadrantPipe_bits_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_29 <= quadrantPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_28) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_29 <= quadrantPipe_bits_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_30 <= quadrantPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_29) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_30 <= quadrantPipe_bits_29; // @[Reg.scala 17:22]
    end
    if (quadrantPipe_valid_30) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_31 <= quadrantPipe_bits_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      trigonometric_io_theta_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      trigonometric_io_theta_v <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      trigonometric_io_theta_b <= theta; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      cosinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      cosinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_cosine_T_2) begin // @[BoxMuller.scala 69:8]
        cosinePipe_bits <= trigonometric_io_result_bits_cosine;
      end else begin
        cosinePipe_bits <= _cosine_T_5;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      sinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_sine_T_2) begin // @[BoxMuller.scala 77:8]
        sinePipe_bits <= trigonometric_io_result_bits_sine;
      end else begin
        sinePipe_bits <= _sine_T_5;
      end
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      signPipe_bits <= rng2_io_rand_bits[31]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sqrt_log_io_uniform_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sqrt_log_io_uniform_v <= rng2_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      sqrt_log_io_uniform_b <= _sqrt_log_io_uniform_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sign_adjustedPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sign_adjustedPipe_valid <= sqrt_log_io_result_valid; // @[Valid.scala 127:22]
    end
    if (sqrt_log_io_result_valid) begin // @[Reg.scala 17:18]
      if (signPipe_bits) begin // @[BoxMuller.scala 91:8]
        sign_adjustedPipe_bits <= _sign_adjusted_T_3;
      end else begin
        sign_adjustedPipe_bits <= sqrt_log_io_result_bits;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g1_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g1_v <= _io_g1_T; // @[Valid.scala 127:22]
    end
    if (_io_g1_T) begin // @[Reg.scala 17:18]
      io_g1_b <= _io_g1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g2_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g2_v <= _io_g2_T; // @[Valid.scala 127:22]
    end
    if (_io_g2_T) begin // @[Reg.scala 17:18]
      io_g2_b <= _io_g2_T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quadrantPipe_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  quadrantPipe_bits = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  quadrantPipe_valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  quadrantPipe_bits_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  quadrantPipe_valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  quadrantPipe_bits_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  quadrantPipe_valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quadrantPipe_bits_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  quadrantPipe_valid_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  quadrantPipe_bits_4 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  quadrantPipe_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  quadrantPipe_bits_5 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  quadrantPipe_valid_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  quadrantPipe_bits_6 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  quadrantPipe_valid_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  quadrantPipe_bits_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  quadrantPipe_valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  quadrantPipe_bits_8 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  quadrantPipe_valid_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  quadrantPipe_bits_9 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  quadrantPipe_valid_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  quadrantPipe_bits_10 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  quadrantPipe_valid_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  quadrantPipe_bits_11 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  quadrantPipe_valid_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  quadrantPipe_bits_12 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  quadrantPipe_valid_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  quadrantPipe_bits_13 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  quadrantPipe_valid_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  quadrantPipe_bits_14 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  quadrantPipe_valid_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  quadrantPipe_bits_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  quadrantPipe_valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  quadrantPipe_bits_16 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  quadrantPipe_valid_17 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  quadrantPipe_bits_17 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  quadrantPipe_valid_18 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  quadrantPipe_bits_18 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  quadrantPipe_valid_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  quadrantPipe_bits_19 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  quadrantPipe_valid_20 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  quadrantPipe_bits_20 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  quadrantPipe_valid_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  quadrantPipe_bits_21 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  quadrantPipe_valid_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  quadrantPipe_bits_22 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  quadrantPipe_valid_23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  quadrantPipe_bits_23 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  quadrantPipe_valid_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  quadrantPipe_bits_24 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  quadrantPipe_valid_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  quadrantPipe_bits_25 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  quadrantPipe_valid_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  quadrantPipe_bits_26 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  quadrantPipe_valid_27 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  quadrantPipe_bits_27 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  quadrantPipe_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  quadrantPipe_bits_28 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  quadrantPipe_valid_29 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  quadrantPipe_bits_29 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  quadrantPipe_valid_30 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  quadrantPipe_bits_30 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  quadrantPipe_bits_31 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  trigonometric_io_theta_v = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  trigonometric_io_theta_b = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cosinePipe_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cosinePipe_bits = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sinePipe_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sinePipe_bits = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  signPipe_bits = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sqrt_log_io_uniform_v = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sqrt_log_io_uniform_b = _RAND_71[28:0];
  _RAND_72 = {1{`RANDOM}};
  sign_adjustedPipe_valid = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  sign_adjustedPipe_bits = _RAND_73[51:0];
  _RAND_74 = {1{`RANDOM}};
  io_g1_v = _RAND_74[0:0];
  _RAND_75 = {3{`RANDOM}};
  io_g1_b = _RAND_75[83:0];
  _RAND_76 = {1{`RANDOM}};
  io_g2_v = _RAND_76[0:0];
  _RAND_77 = {3{`RANDOM}};
  io_g2_b = _RAND_77[83:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MonteCarlo_8(
  input         clock,
  input         reset,
  output        io_request_0_ready,
  input         io_request_0_valid,
  input  [31:0] io_request_0_bits_time_steps,
  input  [31:0] io_request_0_bits_start_value,
  input  [31:0] io_request_0_bits_coefficient1,
  input  [31:0] io_request_0_bits_coefficient2,
  output        io_request_1_ready,
  input         io_request_1_valid,
  input  [31:0] io_request_1_bits_time_steps,
  input  [31:0] io_request_1_bits_start_value,
  input  [31:0] io_request_1_bits_coefficient1,
  input  [31:0] io_request_1_bits_coefficient2,
  input         io_response_0_ready,
  output        io_response_0_valid,
  output [31:0] io_response_0_bits,
  input         io_response_1_ready,
  output        io_response_1_valid,
  output [31:0] io_response_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rng_clock; // @[MonteCarlo.scala 42:19]
  wire  rng_reset; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g1_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g1_bits; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g2_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g2_bits; // @[MonteCarlo.scala 42:19]
  wire  initialized = rng_io_g1_valid & rng_io_g2_valid; // @[MonteCarlo.scala 47:37]
  reg [2:0] state; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_2 = $signed(io_request_0_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_3 = io_request_0_ready & io_request_0_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1; // @[Reg.scala 16:16]
  reg [31:0] c2; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_1 = io_request_0_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step; // @[Reg.scala 16:16]
  reg [31:0] price; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T = $signed(price) * $signed(c1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T = $signed(rng_io_g1_bits) * $signed(c2); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T = $signed(price) * $signed(partial_res2); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_2 = $signed(partial_res3) + $signed(partial_res1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_3 = counter == last_step ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_4 = counter == last_step ? counter : _counter_T_1; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_7 = io_response_0_ready & io_response_0_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_5 = _T_7 ? 3'h1 : state; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_6 = 3'h5 == state ? _GEN_5 : state; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_7 = 3'h4 == state ? $signed(_price_T_2) : $signed(price); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_3 : _GEN_6; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_9 = 3'h4 == state ? _GEN_4 : counter; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_64 = {$signed(partial_res3), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_10 = 3'h3 == state ? $signed(_partial_res3_T) : $signed({{12{_GEN_64[51]}},_GEN_64}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_11 = 3'h3 == state ? 3'h4 : _GEN_8; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_65 = {$signed(partial_res1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_14 = 3'h2 == state ? $signed(_partial_res1_T) : $signed({{12{_GEN_65[51]}},_GEN_65}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_66 = {$signed(partial_res2), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_15 = 3'h2 == state ? $signed(_partial_res2_T) : $signed({{20{_GEN_66[63]}},_GEN_66}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_17 = 3'h2 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_10); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_23 = 3'h1 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_14); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_24 = 3'h1 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_15); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_25 = 3'h1 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_17); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_29 = 3'h0 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_23); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_30 = 3'h0 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_24); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_31 = 3'h0 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_25); // @[MonteCarlo.scala 66:19 60:27]
  reg [2:0] state_1; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_6 = $signed(io_request_1_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_7 = io_request_1_ready & io_request_1_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1_1; // @[Reg.scala 16:16]
  reg [31:0] c2_1; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_4 = io_request_1_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step_1; // @[Reg.scala 16:16]
  reg [31:0] price_1; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1_1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2_1; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3_1; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter_1; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T_1 = $signed(price_1) * $signed(c1_1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T_1 = $signed(rng_io_g2_bits) * $signed(c2_1); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T_1 = $signed(price_1) * $signed(partial_res2_1); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_5 = $signed(partial_res3_1) + $signed(partial_res1_1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_35 = counter_1 == last_step_1 ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_36 = counter_1 == last_step_1 ? counter_1 : _counter_T_3; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_15 = io_response_1_ready & io_response_1_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_37 = _T_15 ? 3'h1 : state_1; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_38 = 3'h5 == state_1 ? _GEN_37 : state_1; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_39 = 3'h4 == state_1 ? $signed(_price_T_5) : $signed(price_1); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_40 = 3'h4 == state_1 ? _GEN_35 : _GEN_38; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_41 = 3'h4 == state_1 ? _GEN_36 : counter_1; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_74 = {$signed(partial_res3_1), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_42 = 3'h3 == state_1 ? $signed(_partial_res3_T_1) : $signed({{12{_GEN_74[51]}},_GEN_74}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_43 = 3'h3 == state_1 ? 3'h4 : _GEN_40; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_75 = {$signed(partial_res1_1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_46 = 3'h2 == state_1 ? $signed(_partial_res1_T_1) : $signed({{12{_GEN_75[51]}},_GEN_75}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_76 = {$signed(partial_res2_1), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_47 = 3'h2 == state_1 ? $signed(_partial_res2_T_1) : $signed({{20{_GEN_76[63]}},_GEN_76}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_49 = 3'h2 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_42); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_55 = 3'h1 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_46); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_56 = 3'h1 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_47); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_57 = 3'h1 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_49); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_61 = 3'h0 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_55); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_62 = 3'h0 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_56); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_63 = 3'h0 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_57); // @[MonteCarlo.scala 66:19 60:27]
  wire [43:0] _GEN_84 = _GEN_29[63:20];
  wire [51:0] _GEN_86 = _GEN_30[83:32];
  wire [43:0] _GEN_88 = _GEN_31[63:20];
  wire [43:0] _GEN_90 = _GEN_61[63:20];
  wire [51:0] _GEN_92 = _GEN_62[83:32];
  wire [43:0] _GEN_94 = _GEN_63[63:20];
  BoxMuller_8 rng ( // @[MonteCarlo.scala 42:19]
    .clock(rng_clock),
    .reset(rng_reset),
    .io_g1_valid(rng_io_g1_valid),
    .io_g1_bits(rng_io_g1_bits),
    .io_g2_valid(rng_io_g2_valid),
    .io_g2_bits(rng_io_g2_bits)
  );
  assign io_request_0_ready = state == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_request_1_ready = state_1 == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_response_0_valid = state == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_0_bits = price; // @[MonteCarlo.scala 65:16]
  assign io_response_1_valid = state_1 == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_1_bits = price_1; // @[MonteCarlo.scala 65:16]
  assign rng_clock = clock;
  assign rng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state <= 3'h1;
      end else begin
        state <= 3'h0;
      end
    end else if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_3) begin // @[MonteCarlo.scala 71:23]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[MonteCarlo.scala 66:19]
      state <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state <= _GEN_11;
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c1 <= _c1_T_2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c2 <= io_request_0_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      last_step <= _last_step_T_1; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        price <= io_request_0_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          price <= _GEN_7;
        end
      end
    end
    partial_res1 <= _GEN_84[31:0];
    partial_res2 <= _GEN_86[31:0];
    partial_res3 <= _GEN_88[31:0];
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        counter <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          counter <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state_1 <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state_1 <= 3'h1;
      end else begin
        state_1 <= 3'h0;
      end
    end else if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_7) begin // @[MonteCarlo.scala 71:23]
        state_1 <= 3'h2;
      end else begin
        state_1 <= 3'h1;
      end
    end else if (3'h2 == state_1) begin // @[MonteCarlo.scala 66:19]
      state_1 <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state_1 <= _GEN_43;
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c1_1 <= _c1_T_6; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c2_1 <= io_request_1_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      last_step_1 <= _last_step_T_4; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        price_1 <= io_request_1_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          price_1 <= _GEN_39;
        end
      end
    end
    partial_res1_1 <= _GEN_90[31:0];
    partial_res2_1 <= _GEN_92[31:0];
    partial_res3_1 <= _GEN_94[31:0];
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        counter_1 <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          counter_1 <= _GEN_41;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  c1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_step = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  price = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  partial_res1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  partial_res2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  partial_res3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  c1_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_step_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  price_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  partial_res1_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  partial_res2_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  partial_res3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  counter_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_18(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h398eb463 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h3f04e6b0 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h8927864 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_19(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h22f3c07c : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h550e4f3 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'hbe74129 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoxMuller_9(
  input         clock,
  input         reset,
  output        io_g1_valid,
  output [51:0] io_g1_bits,
  output        io_g2_valid,
  output [51:0] io_g2_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [95:0] _RAND_77;
`endif // RANDOMIZE_REG_INIT
  wire  rng1_clock; // @[BoxMuller.scala 51:20]
  wire  rng1_reset; // @[BoxMuller.scala 51:20]
  wire  rng1_io_rand_valid; // @[BoxMuller.scala 51:20]
  wire [31:0] rng1_io_rand_bits; // @[BoxMuller.scala 51:20]
  wire  rng2_clock; // @[BoxMuller.scala 52:20]
  wire  rng2_reset; // @[BoxMuller.scala 52:20]
  wire  rng2_io_rand_valid; // @[BoxMuller.scala 52:20]
  wire [31:0] rng2_io_rand_bits; // @[BoxMuller.scala 52:20]
  wire  trigonometric_clock; // @[BoxMuller.scala 55:29]
  wire  trigonometric_reset; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_theta_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_theta_bits; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_result_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_sine; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_cosine; // @[BoxMuller.scala 55:29]
  wire  sqrt_log_clock; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_reset; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_uniform_valid; // @[BoxMuller.scala 84:24]
  wire [31:0] sqrt_log_io_uniform_bits; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_result_valid; // @[BoxMuller.scala 84:24]
  wire [51:0] sqrt_log_io_result_bits; // @[BoxMuller.scala 84:24]
  wire [30:0] _theta_T_3 = {2'h0,rng1_io_rand_bits[28:0]}; // @[BoxMuller.scala 62:18]
  wire [62:0] _theta_T_4 = $signed(_theta_T_3) * 32'sh6487ed51; // @[BoxMuller.scala 62:26]
  reg  quadrantPipe_valid; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_1; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_1; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_2; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_2; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_3; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_3; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_4; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_4; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_5; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_5; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_6; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_6; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_7; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_7; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_8; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_8; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_9; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_9; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_10; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_10; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_11; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_11; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_12; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_12; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_13; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_13; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_14; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_14; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_15; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_15; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_16; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_16; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_17; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_17; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_18; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_18; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_19; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_19; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_20; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_20; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_21; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_21; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_22; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_22; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_23; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_23; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_24; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_24; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_25; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_25; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_26; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_26; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_27; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_27; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_28; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_28; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_29; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_29; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_30; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_30; // @[Reg.scala 16:16]
  reg [1:0] quadrantPipe_bits_31; // @[Reg.scala 16:16]
  reg  trigonometric_io_theta_v; // @[Valid.scala 127:22]
  reg [31:0] trigonometric_io_theta_b; // @[Reg.scala 16:16]
  wire [33:0] _GEN_40 = _theta_T_4[62:29]; // @[BoxMuller.scala 59:19 61:9]
  wire [31:0] theta = _GEN_40[31:0]; // @[BoxMuller.scala 59:19 61:9]
  wire  _cosine_T = quadrantPipe_bits_31 == 2'h0; // @[BoxMuller.scala 70:21]
  wire  _cosine_T_2 = quadrantPipe_bits_31 == 2'h0 | quadrantPipe_bits_31 == 2'h3; // @[BoxMuller.scala 70:29]
  wire [31:0] _cosine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_cosine); // @[BoxMuller.scala 72:7]
  reg  cosinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] cosinePipe_bits; // @[Reg.scala 16:16]
  wire  _sine_T_2 = _cosine_T | quadrantPipe_bits_31 == 2'h2; // @[BoxMuller.scala 78:29]
  wire [31:0] _sine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_sine); // @[BoxMuller.scala 80:7]
  reg  sinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] sinePipe_bits; // @[Reg.scala 16:16]
  reg  signPipe_bits; // @[Reg.scala 16:16]
  wire [28:0] _sqrt_log_io_uniform_T_1 = rng2_io_rand_bits[28:0]; // @[BoxMuller.scala 87:89]
  reg  sqrt_log_io_uniform_v; // @[Valid.scala 127:22]
  reg [28:0] sqrt_log_io_uniform_b; // @[Reg.scala 16:16]
  wire [51:0] _sign_adjusted_T_3 = 52'sh0 - $signed(sqrt_log_io_result_bits); // @[BoxMuller.scala 93:7]
  reg  sign_adjustedPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] sign_adjustedPipe_bits; // @[Reg.scala 16:16]
  wire  _io_g1_T = sign_adjustedPipe_valid & cosinePipe_valid; // @[BoxMuller.scala 99:25]
  wire [83:0] _io_g1_T_1 = $signed(cosinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 100:17]
  reg  io_g1_v; // @[Valid.scala 127:22]
  reg [83:0] io_g1_b; // @[Reg.scala 16:16]
  wire  _io_g2_T = sign_adjustedPipe_valid & sinePipe_valid; // @[BoxMuller.scala 103:25]
  wire [83:0] _io_g2_T_1 = $signed(sinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 104:15]
  reg  io_g2_v; // @[Valid.scala 127:22]
  reg [83:0] io_g2_b; // @[Reg.scala 16:16]
  wire [53:0] _GEN_42 = io_g1_b[83:30]; // @[BoxMuller.scala 98:9]
  wire [53:0] _GEN_44 = io_g2_b[83:30]; // @[BoxMuller.scala 102:9]
  wire [32:0] _GEN_46 = {$signed(trigonometric_io_theta_b), 1'h0}; // @[BoxMuller.scala 65:26]
  TauswortheUniform_18 rng1 ( // @[BoxMuller.scala 51:20]
    .clock(rng1_clock),
    .reset(rng1_reset),
    .io_rand_valid(rng1_io_rand_valid),
    .io_rand_bits(rng1_io_rand_bits)
  );
  TauswortheUniform_19 rng2 ( // @[BoxMuller.scala 52:20]
    .clock(rng2_clock),
    .reset(rng2_reset),
    .io_rand_valid(rng2_io_rand_valid),
    .io_rand_bits(rng2_io_rand_bits)
  );
  Trigonometric trigonometric ( // @[BoxMuller.scala 55:29]
    .clock(trigonometric_clock),
    .reset(trigonometric_reset),
    .io_theta_valid(trigonometric_io_theta_valid),
    .io_theta_bits(trigonometric_io_theta_bits),
    .io_result_valid(trigonometric_io_result_valid),
    .io_result_bits_sine(trigonometric_io_result_bits_sine),
    .io_result_bits_cosine(trigonometric_io_result_bits_cosine)
  );
  SquareRootLog sqrt_log ( // @[BoxMuller.scala 84:24]
    .clock(sqrt_log_clock),
    .reset(sqrt_log_reset),
    .io_uniform_valid(sqrt_log_io_uniform_valid),
    .io_uniform_bits(sqrt_log_io_uniform_bits),
    .io_result_valid(sqrt_log_io_result_valid),
    .io_result_bits(sqrt_log_io_result_bits)
  );
  assign io_g1_valid = io_g1_v; // @[Valid.scala 122:21 123:17]
  assign io_g1_bits = _GEN_42[51:0]; // @[BoxMuller.scala 98:9]
  assign io_g2_valid = io_g2_v; // @[Valid.scala 122:21 123:17]
  assign io_g2_bits = _GEN_44[51:0]; // @[BoxMuller.scala 102:9]
  assign rng1_clock = clock;
  assign rng1_reset = reset;
  assign rng2_clock = clock;
  assign rng2_reset = reset;
  assign trigonometric_clock = clock;
  assign trigonometric_reset = reset;
  assign trigonometric_io_theta_valid = trigonometric_io_theta_v; // @[Valid.scala 122:21 123:17]
  assign trigonometric_io_theta_bits = _GEN_46[31:0]; // @[BoxMuller.scala 65:26]
  assign sqrt_log_clock = clock;
  assign sqrt_log_reset = reset;
  assign sqrt_log_io_uniform_valid = sqrt_log_io_uniform_v; // @[Valid.scala 122:21 123:17]
  assign sqrt_log_io_uniform_bits = {{3{sqrt_log_io_uniform_b[28]}},sqrt_log_io_uniform_b}; // @[BoxMuller.scala 87:23]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits <= rng1_io_rand_bits[31:30]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_1 <= quadrantPipe_valid; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_1 <= quadrantPipe_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_2 <= quadrantPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_1) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_2 <= quadrantPipe_bits_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_3 <= quadrantPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_2) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_3 <= quadrantPipe_bits_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_4 <= quadrantPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_3) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_4 <= quadrantPipe_bits_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_5 <= quadrantPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_4) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_5 <= quadrantPipe_bits_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_6 <= quadrantPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_5) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_6 <= quadrantPipe_bits_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_7 <= quadrantPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_6) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_7 <= quadrantPipe_bits_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_8 <= quadrantPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_7) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_8 <= quadrantPipe_bits_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_9 <= quadrantPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_8) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_9 <= quadrantPipe_bits_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_10 <= quadrantPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_9) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_10 <= quadrantPipe_bits_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_11 <= quadrantPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_10) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_11 <= quadrantPipe_bits_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_12 <= quadrantPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_11) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_12 <= quadrantPipe_bits_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_13 <= quadrantPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_12) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_13 <= quadrantPipe_bits_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_14 <= quadrantPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_13) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_14 <= quadrantPipe_bits_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_15 <= quadrantPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_14) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_15 <= quadrantPipe_bits_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_16 <= quadrantPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_15) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_16 <= quadrantPipe_bits_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_17 <= quadrantPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_16) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_17 <= quadrantPipe_bits_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_18 <= quadrantPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_17) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_18 <= quadrantPipe_bits_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_19 <= quadrantPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_18) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_19 <= quadrantPipe_bits_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_20 <= quadrantPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_19) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_20 <= quadrantPipe_bits_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_21 <= quadrantPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_20) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_21 <= quadrantPipe_bits_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_22 <= quadrantPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_21) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_22 <= quadrantPipe_bits_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_23 <= quadrantPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_22) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_23 <= quadrantPipe_bits_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_24 <= quadrantPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_23) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_24 <= quadrantPipe_bits_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_25 <= quadrantPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_24) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_25 <= quadrantPipe_bits_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_26 <= quadrantPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_25) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_26 <= quadrantPipe_bits_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_27 <= quadrantPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_26) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_27 <= quadrantPipe_bits_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_28 <= quadrantPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_27) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_28 <= quadrantPipe_bits_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_29 <= quadrantPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_28) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_29 <= quadrantPipe_bits_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_30 <= quadrantPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_29) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_30 <= quadrantPipe_bits_29; // @[Reg.scala 17:22]
    end
    if (quadrantPipe_valid_30) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_31 <= quadrantPipe_bits_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      trigonometric_io_theta_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      trigonometric_io_theta_v <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      trigonometric_io_theta_b <= theta; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      cosinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      cosinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_cosine_T_2) begin // @[BoxMuller.scala 69:8]
        cosinePipe_bits <= trigonometric_io_result_bits_cosine;
      end else begin
        cosinePipe_bits <= _cosine_T_5;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      sinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_sine_T_2) begin // @[BoxMuller.scala 77:8]
        sinePipe_bits <= trigonometric_io_result_bits_sine;
      end else begin
        sinePipe_bits <= _sine_T_5;
      end
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      signPipe_bits <= rng2_io_rand_bits[31]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sqrt_log_io_uniform_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sqrt_log_io_uniform_v <= rng2_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      sqrt_log_io_uniform_b <= _sqrt_log_io_uniform_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sign_adjustedPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sign_adjustedPipe_valid <= sqrt_log_io_result_valid; // @[Valid.scala 127:22]
    end
    if (sqrt_log_io_result_valid) begin // @[Reg.scala 17:18]
      if (signPipe_bits) begin // @[BoxMuller.scala 91:8]
        sign_adjustedPipe_bits <= _sign_adjusted_T_3;
      end else begin
        sign_adjustedPipe_bits <= sqrt_log_io_result_bits;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g1_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g1_v <= _io_g1_T; // @[Valid.scala 127:22]
    end
    if (_io_g1_T) begin // @[Reg.scala 17:18]
      io_g1_b <= _io_g1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g2_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g2_v <= _io_g2_T; // @[Valid.scala 127:22]
    end
    if (_io_g2_T) begin // @[Reg.scala 17:18]
      io_g2_b <= _io_g2_T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quadrantPipe_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  quadrantPipe_bits = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  quadrantPipe_valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  quadrantPipe_bits_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  quadrantPipe_valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  quadrantPipe_bits_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  quadrantPipe_valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quadrantPipe_bits_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  quadrantPipe_valid_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  quadrantPipe_bits_4 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  quadrantPipe_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  quadrantPipe_bits_5 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  quadrantPipe_valid_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  quadrantPipe_bits_6 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  quadrantPipe_valid_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  quadrantPipe_bits_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  quadrantPipe_valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  quadrantPipe_bits_8 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  quadrantPipe_valid_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  quadrantPipe_bits_9 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  quadrantPipe_valid_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  quadrantPipe_bits_10 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  quadrantPipe_valid_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  quadrantPipe_bits_11 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  quadrantPipe_valid_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  quadrantPipe_bits_12 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  quadrantPipe_valid_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  quadrantPipe_bits_13 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  quadrantPipe_valid_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  quadrantPipe_bits_14 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  quadrantPipe_valid_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  quadrantPipe_bits_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  quadrantPipe_valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  quadrantPipe_bits_16 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  quadrantPipe_valid_17 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  quadrantPipe_bits_17 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  quadrantPipe_valid_18 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  quadrantPipe_bits_18 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  quadrantPipe_valid_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  quadrantPipe_bits_19 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  quadrantPipe_valid_20 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  quadrantPipe_bits_20 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  quadrantPipe_valid_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  quadrantPipe_bits_21 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  quadrantPipe_valid_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  quadrantPipe_bits_22 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  quadrantPipe_valid_23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  quadrantPipe_bits_23 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  quadrantPipe_valid_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  quadrantPipe_bits_24 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  quadrantPipe_valid_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  quadrantPipe_bits_25 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  quadrantPipe_valid_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  quadrantPipe_bits_26 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  quadrantPipe_valid_27 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  quadrantPipe_bits_27 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  quadrantPipe_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  quadrantPipe_bits_28 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  quadrantPipe_valid_29 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  quadrantPipe_bits_29 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  quadrantPipe_valid_30 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  quadrantPipe_bits_30 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  quadrantPipe_bits_31 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  trigonometric_io_theta_v = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  trigonometric_io_theta_b = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cosinePipe_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cosinePipe_bits = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sinePipe_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sinePipe_bits = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  signPipe_bits = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sqrt_log_io_uniform_v = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sqrt_log_io_uniform_b = _RAND_71[28:0];
  _RAND_72 = {1{`RANDOM}};
  sign_adjustedPipe_valid = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  sign_adjustedPipe_bits = _RAND_73[51:0];
  _RAND_74 = {1{`RANDOM}};
  io_g1_v = _RAND_74[0:0];
  _RAND_75 = {3{`RANDOM}};
  io_g1_b = _RAND_75[83:0];
  _RAND_76 = {1{`RANDOM}};
  io_g2_v = _RAND_76[0:0];
  _RAND_77 = {3{`RANDOM}};
  io_g2_b = _RAND_77[83:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MonteCarlo_9(
  input         clock,
  input         reset,
  output        io_request_0_ready,
  input         io_request_0_valid,
  input  [31:0] io_request_0_bits_time_steps,
  input  [31:0] io_request_0_bits_start_value,
  input  [31:0] io_request_0_bits_coefficient1,
  input  [31:0] io_request_0_bits_coefficient2,
  output        io_request_1_ready,
  input         io_request_1_valid,
  input  [31:0] io_request_1_bits_time_steps,
  input  [31:0] io_request_1_bits_start_value,
  input  [31:0] io_request_1_bits_coefficient1,
  input  [31:0] io_request_1_bits_coefficient2,
  input         io_response_0_ready,
  output        io_response_0_valid,
  output [31:0] io_response_0_bits,
  input         io_response_1_ready,
  output        io_response_1_valid,
  output [31:0] io_response_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rng_clock; // @[MonteCarlo.scala 42:19]
  wire  rng_reset; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g1_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g1_bits; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g2_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g2_bits; // @[MonteCarlo.scala 42:19]
  wire  initialized = rng_io_g1_valid & rng_io_g2_valid; // @[MonteCarlo.scala 47:37]
  reg [2:0] state; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_2 = $signed(io_request_0_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_3 = io_request_0_ready & io_request_0_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1; // @[Reg.scala 16:16]
  reg [31:0] c2; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_1 = io_request_0_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step; // @[Reg.scala 16:16]
  reg [31:0] price; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T = $signed(price) * $signed(c1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T = $signed(rng_io_g1_bits) * $signed(c2); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T = $signed(price) * $signed(partial_res2); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_2 = $signed(partial_res3) + $signed(partial_res1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_3 = counter == last_step ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_4 = counter == last_step ? counter : _counter_T_1; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_7 = io_response_0_ready & io_response_0_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_5 = _T_7 ? 3'h1 : state; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_6 = 3'h5 == state ? _GEN_5 : state; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_7 = 3'h4 == state ? $signed(_price_T_2) : $signed(price); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_3 : _GEN_6; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_9 = 3'h4 == state ? _GEN_4 : counter; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_64 = {$signed(partial_res3), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_10 = 3'h3 == state ? $signed(_partial_res3_T) : $signed({{12{_GEN_64[51]}},_GEN_64}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_11 = 3'h3 == state ? 3'h4 : _GEN_8; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_65 = {$signed(partial_res1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_14 = 3'h2 == state ? $signed(_partial_res1_T) : $signed({{12{_GEN_65[51]}},_GEN_65}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_66 = {$signed(partial_res2), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_15 = 3'h2 == state ? $signed(_partial_res2_T) : $signed({{20{_GEN_66[63]}},_GEN_66}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_17 = 3'h2 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_10); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_23 = 3'h1 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_14); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_24 = 3'h1 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_15); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_25 = 3'h1 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_17); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_29 = 3'h0 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_23); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_30 = 3'h0 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_24); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_31 = 3'h0 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_25); // @[MonteCarlo.scala 66:19 60:27]
  reg [2:0] state_1; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_6 = $signed(io_request_1_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_7 = io_request_1_ready & io_request_1_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1_1; // @[Reg.scala 16:16]
  reg [31:0] c2_1; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_4 = io_request_1_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step_1; // @[Reg.scala 16:16]
  reg [31:0] price_1; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1_1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2_1; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3_1; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter_1; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T_1 = $signed(price_1) * $signed(c1_1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T_1 = $signed(rng_io_g2_bits) * $signed(c2_1); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T_1 = $signed(price_1) * $signed(partial_res2_1); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_5 = $signed(partial_res3_1) + $signed(partial_res1_1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_35 = counter_1 == last_step_1 ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_36 = counter_1 == last_step_1 ? counter_1 : _counter_T_3; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_15 = io_response_1_ready & io_response_1_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_37 = _T_15 ? 3'h1 : state_1; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_38 = 3'h5 == state_1 ? _GEN_37 : state_1; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_39 = 3'h4 == state_1 ? $signed(_price_T_5) : $signed(price_1); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_40 = 3'h4 == state_1 ? _GEN_35 : _GEN_38; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_41 = 3'h4 == state_1 ? _GEN_36 : counter_1; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_74 = {$signed(partial_res3_1), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_42 = 3'h3 == state_1 ? $signed(_partial_res3_T_1) : $signed({{12{_GEN_74[51]}},_GEN_74}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_43 = 3'h3 == state_1 ? 3'h4 : _GEN_40; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_75 = {$signed(partial_res1_1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_46 = 3'h2 == state_1 ? $signed(_partial_res1_T_1) : $signed({{12{_GEN_75[51]}},_GEN_75}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_76 = {$signed(partial_res2_1), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_47 = 3'h2 == state_1 ? $signed(_partial_res2_T_1) : $signed({{20{_GEN_76[63]}},_GEN_76}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_49 = 3'h2 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_42); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_55 = 3'h1 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_46); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_56 = 3'h1 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_47); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_57 = 3'h1 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_49); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_61 = 3'h0 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_55); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_62 = 3'h0 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_56); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_63 = 3'h0 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_57); // @[MonteCarlo.scala 66:19 60:27]
  wire [43:0] _GEN_84 = _GEN_29[63:20];
  wire [51:0] _GEN_86 = _GEN_30[83:32];
  wire [43:0] _GEN_88 = _GEN_31[63:20];
  wire [43:0] _GEN_90 = _GEN_61[63:20];
  wire [51:0] _GEN_92 = _GEN_62[83:32];
  wire [43:0] _GEN_94 = _GEN_63[63:20];
  BoxMuller_9 rng ( // @[MonteCarlo.scala 42:19]
    .clock(rng_clock),
    .reset(rng_reset),
    .io_g1_valid(rng_io_g1_valid),
    .io_g1_bits(rng_io_g1_bits),
    .io_g2_valid(rng_io_g2_valid),
    .io_g2_bits(rng_io_g2_bits)
  );
  assign io_request_0_ready = state == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_request_1_ready = state_1 == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_response_0_valid = state == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_0_bits = price; // @[MonteCarlo.scala 65:16]
  assign io_response_1_valid = state_1 == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_1_bits = price_1; // @[MonteCarlo.scala 65:16]
  assign rng_clock = clock;
  assign rng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state <= 3'h1;
      end else begin
        state <= 3'h0;
      end
    end else if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_3) begin // @[MonteCarlo.scala 71:23]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[MonteCarlo.scala 66:19]
      state <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state <= _GEN_11;
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c1 <= _c1_T_2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c2 <= io_request_0_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      last_step <= _last_step_T_1; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        price <= io_request_0_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          price <= _GEN_7;
        end
      end
    end
    partial_res1 <= _GEN_84[31:0];
    partial_res2 <= _GEN_86[31:0];
    partial_res3 <= _GEN_88[31:0];
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        counter <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          counter <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state_1 <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state_1 <= 3'h1;
      end else begin
        state_1 <= 3'h0;
      end
    end else if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_7) begin // @[MonteCarlo.scala 71:23]
        state_1 <= 3'h2;
      end else begin
        state_1 <= 3'h1;
      end
    end else if (3'h2 == state_1) begin // @[MonteCarlo.scala 66:19]
      state_1 <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state_1 <= _GEN_43;
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c1_1 <= _c1_T_6; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c2_1 <= io_request_1_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      last_step_1 <= _last_step_T_4; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        price_1 <= io_request_1_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          price_1 <= _GEN_39;
        end
      end
    end
    partial_res1_1 <= _GEN_90[31:0];
    partial_res2_1 <= _GEN_92[31:0];
    partial_res3_1 <= _GEN_94[31:0];
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        counter_1 <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          counter_1 <= _GEN_41;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  c1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_step = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  price = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  partial_res1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  partial_res2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  partial_res3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  c1_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_step_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  price_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  partial_res1_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  partial_res2_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  partial_res3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  counter_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_20(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h3ea0f641 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h13a3c6ea : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h2e3b195c : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_21(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h2af2e9c5 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h2dc31170 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h41d0f0a : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoxMuller_10(
  input         clock,
  input         reset,
  output        io_g1_valid,
  output [51:0] io_g1_bits,
  output        io_g2_valid,
  output [51:0] io_g2_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [95:0] _RAND_77;
`endif // RANDOMIZE_REG_INIT
  wire  rng1_clock; // @[BoxMuller.scala 51:20]
  wire  rng1_reset; // @[BoxMuller.scala 51:20]
  wire  rng1_io_rand_valid; // @[BoxMuller.scala 51:20]
  wire [31:0] rng1_io_rand_bits; // @[BoxMuller.scala 51:20]
  wire  rng2_clock; // @[BoxMuller.scala 52:20]
  wire  rng2_reset; // @[BoxMuller.scala 52:20]
  wire  rng2_io_rand_valid; // @[BoxMuller.scala 52:20]
  wire [31:0] rng2_io_rand_bits; // @[BoxMuller.scala 52:20]
  wire  trigonometric_clock; // @[BoxMuller.scala 55:29]
  wire  trigonometric_reset; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_theta_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_theta_bits; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_result_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_sine; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_cosine; // @[BoxMuller.scala 55:29]
  wire  sqrt_log_clock; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_reset; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_uniform_valid; // @[BoxMuller.scala 84:24]
  wire [31:0] sqrt_log_io_uniform_bits; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_result_valid; // @[BoxMuller.scala 84:24]
  wire [51:0] sqrt_log_io_result_bits; // @[BoxMuller.scala 84:24]
  wire [30:0] _theta_T_3 = {2'h0,rng1_io_rand_bits[28:0]}; // @[BoxMuller.scala 62:18]
  wire [62:0] _theta_T_4 = $signed(_theta_T_3) * 32'sh6487ed51; // @[BoxMuller.scala 62:26]
  reg  quadrantPipe_valid; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_1; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_1; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_2; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_2; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_3; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_3; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_4; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_4; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_5; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_5; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_6; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_6; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_7; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_7; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_8; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_8; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_9; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_9; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_10; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_10; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_11; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_11; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_12; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_12; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_13; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_13; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_14; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_14; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_15; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_15; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_16; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_16; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_17; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_17; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_18; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_18; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_19; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_19; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_20; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_20; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_21; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_21; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_22; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_22; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_23; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_23; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_24; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_24; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_25; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_25; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_26; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_26; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_27; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_27; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_28; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_28; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_29; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_29; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_30; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_30; // @[Reg.scala 16:16]
  reg [1:0] quadrantPipe_bits_31; // @[Reg.scala 16:16]
  reg  trigonometric_io_theta_v; // @[Valid.scala 127:22]
  reg [31:0] trigonometric_io_theta_b; // @[Reg.scala 16:16]
  wire [33:0] _GEN_40 = _theta_T_4[62:29]; // @[BoxMuller.scala 59:19 61:9]
  wire [31:0] theta = _GEN_40[31:0]; // @[BoxMuller.scala 59:19 61:9]
  wire  _cosine_T = quadrantPipe_bits_31 == 2'h0; // @[BoxMuller.scala 70:21]
  wire  _cosine_T_2 = quadrantPipe_bits_31 == 2'h0 | quadrantPipe_bits_31 == 2'h3; // @[BoxMuller.scala 70:29]
  wire [31:0] _cosine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_cosine); // @[BoxMuller.scala 72:7]
  reg  cosinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] cosinePipe_bits; // @[Reg.scala 16:16]
  wire  _sine_T_2 = _cosine_T | quadrantPipe_bits_31 == 2'h2; // @[BoxMuller.scala 78:29]
  wire [31:0] _sine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_sine); // @[BoxMuller.scala 80:7]
  reg  sinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] sinePipe_bits; // @[Reg.scala 16:16]
  reg  signPipe_bits; // @[Reg.scala 16:16]
  wire [28:0] _sqrt_log_io_uniform_T_1 = rng2_io_rand_bits[28:0]; // @[BoxMuller.scala 87:89]
  reg  sqrt_log_io_uniform_v; // @[Valid.scala 127:22]
  reg [28:0] sqrt_log_io_uniform_b; // @[Reg.scala 16:16]
  wire [51:0] _sign_adjusted_T_3 = 52'sh0 - $signed(sqrt_log_io_result_bits); // @[BoxMuller.scala 93:7]
  reg  sign_adjustedPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] sign_adjustedPipe_bits; // @[Reg.scala 16:16]
  wire  _io_g1_T = sign_adjustedPipe_valid & cosinePipe_valid; // @[BoxMuller.scala 99:25]
  wire [83:0] _io_g1_T_1 = $signed(cosinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 100:17]
  reg  io_g1_v; // @[Valid.scala 127:22]
  reg [83:0] io_g1_b; // @[Reg.scala 16:16]
  wire  _io_g2_T = sign_adjustedPipe_valid & sinePipe_valid; // @[BoxMuller.scala 103:25]
  wire [83:0] _io_g2_T_1 = $signed(sinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 104:15]
  reg  io_g2_v; // @[Valid.scala 127:22]
  reg [83:0] io_g2_b; // @[Reg.scala 16:16]
  wire [53:0] _GEN_42 = io_g1_b[83:30]; // @[BoxMuller.scala 98:9]
  wire [53:0] _GEN_44 = io_g2_b[83:30]; // @[BoxMuller.scala 102:9]
  wire [32:0] _GEN_46 = {$signed(trigonometric_io_theta_b), 1'h0}; // @[BoxMuller.scala 65:26]
  TauswortheUniform_20 rng1 ( // @[BoxMuller.scala 51:20]
    .clock(rng1_clock),
    .reset(rng1_reset),
    .io_rand_valid(rng1_io_rand_valid),
    .io_rand_bits(rng1_io_rand_bits)
  );
  TauswortheUniform_21 rng2 ( // @[BoxMuller.scala 52:20]
    .clock(rng2_clock),
    .reset(rng2_reset),
    .io_rand_valid(rng2_io_rand_valid),
    .io_rand_bits(rng2_io_rand_bits)
  );
  Trigonometric trigonometric ( // @[BoxMuller.scala 55:29]
    .clock(trigonometric_clock),
    .reset(trigonometric_reset),
    .io_theta_valid(trigonometric_io_theta_valid),
    .io_theta_bits(trigonometric_io_theta_bits),
    .io_result_valid(trigonometric_io_result_valid),
    .io_result_bits_sine(trigonometric_io_result_bits_sine),
    .io_result_bits_cosine(trigonometric_io_result_bits_cosine)
  );
  SquareRootLog sqrt_log ( // @[BoxMuller.scala 84:24]
    .clock(sqrt_log_clock),
    .reset(sqrt_log_reset),
    .io_uniform_valid(sqrt_log_io_uniform_valid),
    .io_uniform_bits(sqrt_log_io_uniform_bits),
    .io_result_valid(sqrt_log_io_result_valid),
    .io_result_bits(sqrt_log_io_result_bits)
  );
  assign io_g1_valid = io_g1_v; // @[Valid.scala 122:21 123:17]
  assign io_g1_bits = _GEN_42[51:0]; // @[BoxMuller.scala 98:9]
  assign io_g2_valid = io_g2_v; // @[Valid.scala 122:21 123:17]
  assign io_g2_bits = _GEN_44[51:0]; // @[BoxMuller.scala 102:9]
  assign rng1_clock = clock;
  assign rng1_reset = reset;
  assign rng2_clock = clock;
  assign rng2_reset = reset;
  assign trigonometric_clock = clock;
  assign trigonometric_reset = reset;
  assign trigonometric_io_theta_valid = trigonometric_io_theta_v; // @[Valid.scala 122:21 123:17]
  assign trigonometric_io_theta_bits = _GEN_46[31:0]; // @[BoxMuller.scala 65:26]
  assign sqrt_log_clock = clock;
  assign sqrt_log_reset = reset;
  assign sqrt_log_io_uniform_valid = sqrt_log_io_uniform_v; // @[Valid.scala 122:21 123:17]
  assign sqrt_log_io_uniform_bits = {{3{sqrt_log_io_uniform_b[28]}},sqrt_log_io_uniform_b}; // @[BoxMuller.scala 87:23]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits <= rng1_io_rand_bits[31:30]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_1 <= quadrantPipe_valid; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_1 <= quadrantPipe_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_2 <= quadrantPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_1) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_2 <= quadrantPipe_bits_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_3 <= quadrantPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_2) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_3 <= quadrantPipe_bits_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_4 <= quadrantPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_3) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_4 <= quadrantPipe_bits_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_5 <= quadrantPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_4) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_5 <= quadrantPipe_bits_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_6 <= quadrantPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_5) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_6 <= quadrantPipe_bits_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_7 <= quadrantPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_6) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_7 <= quadrantPipe_bits_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_8 <= quadrantPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_7) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_8 <= quadrantPipe_bits_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_9 <= quadrantPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_8) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_9 <= quadrantPipe_bits_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_10 <= quadrantPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_9) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_10 <= quadrantPipe_bits_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_11 <= quadrantPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_10) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_11 <= quadrantPipe_bits_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_12 <= quadrantPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_11) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_12 <= quadrantPipe_bits_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_13 <= quadrantPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_12) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_13 <= quadrantPipe_bits_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_14 <= quadrantPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_13) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_14 <= quadrantPipe_bits_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_15 <= quadrantPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_14) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_15 <= quadrantPipe_bits_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_16 <= quadrantPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_15) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_16 <= quadrantPipe_bits_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_17 <= quadrantPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_16) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_17 <= quadrantPipe_bits_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_18 <= quadrantPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_17) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_18 <= quadrantPipe_bits_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_19 <= quadrantPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_18) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_19 <= quadrantPipe_bits_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_20 <= quadrantPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_19) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_20 <= quadrantPipe_bits_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_21 <= quadrantPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_20) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_21 <= quadrantPipe_bits_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_22 <= quadrantPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_21) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_22 <= quadrantPipe_bits_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_23 <= quadrantPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_22) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_23 <= quadrantPipe_bits_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_24 <= quadrantPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_23) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_24 <= quadrantPipe_bits_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_25 <= quadrantPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_24) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_25 <= quadrantPipe_bits_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_26 <= quadrantPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_25) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_26 <= quadrantPipe_bits_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_27 <= quadrantPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_26) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_27 <= quadrantPipe_bits_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_28 <= quadrantPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_27) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_28 <= quadrantPipe_bits_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_29 <= quadrantPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_28) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_29 <= quadrantPipe_bits_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_30 <= quadrantPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_29) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_30 <= quadrantPipe_bits_29; // @[Reg.scala 17:22]
    end
    if (quadrantPipe_valid_30) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_31 <= quadrantPipe_bits_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      trigonometric_io_theta_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      trigonometric_io_theta_v <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      trigonometric_io_theta_b <= theta; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      cosinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      cosinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_cosine_T_2) begin // @[BoxMuller.scala 69:8]
        cosinePipe_bits <= trigonometric_io_result_bits_cosine;
      end else begin
        cosinePipe_bits <= _cosine_T_5;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      sinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_sine_T_2) begin // @[BoxMuller.scala 77:8]
        sinePipe_bits <= trigonometric_io_result_bits_sine;
      end else begin
        sinePipe_bits <= _sine_T_5;
      end
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      signPipe_bits <= rng2_io_rand_bits[31]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sqrt_log_io_uniform_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sqrt_log_io_uniform_v <= rng2_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      sqrt_log_io_uniform_b <= _sqrt_log_io_uniform_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sign_adjustedPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sign_adjustedPipe_valid <= sqrt_log_io_result_valid; // @[Valid.scala 127:22]
    end
    if (sqrt_log_io_result_valid) begin // @[Reg.scala 17:18]
      if (signPipe_bits) begin // @[BoxMuller.scala 91:8]
        sign_adjustedPipe_bits <= _sign_adjusted_T_3;
      end else begin
        sign_adjustedPipe_bits <= sqrt_log_io_result_bits;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g1_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g1_v <= _io_g1_T; // @[Valid.scala 127:22]
    end
    if (_io_g1_T) begin // @[Reg.scala 17:18]
      io_g1_b <= _io_g1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g2_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g2_v <= _io_g2_T; // @[Valid.scala 127:22]
    end
    if (_io_g2_T) begin // @[Reg.scala 17:18]
      io_g2_b <= _io_g2_T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quadrantPipe_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  quadrantPipe_bits = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  quadrantPipe_valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  quadrantPipe_bits_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  quadrantPipe_valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  quadrantPipe_bits_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  quadrantPipe_valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quadrantPipe_bits_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  quadrantPipe_valid_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  quadrantPipe_bits_4 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  quadrantPipe_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  quadrantPipe_bits_5 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  quadrantPipe_valid_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  quadrantPipe_bits_6 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  quadrantPipe_valid_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  quadrantPipe_bits_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  quadrantPipe_valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  quadrantPipe_bits_8 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  quadrantPipe_valid_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  quadrantPipe_bits_9 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  quadrantPipe_valid_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  quadrantPipe_bits_10 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  quadrantPipe_valid_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  quadrantPipe_bits_11 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  quadrantPipe_valid_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  quadrantPipe_bits_12 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  quadrantPipe_valid_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  quadrantPipe_bits_13 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  quadrantPipe_valid_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  quadrantPipe_bits_14 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  quadrantPipe_valid_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  quadrantPipe_bits_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  quadrantPipe_valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  quadrantPipe_bits_16 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  quadrantPipe_valid_17 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  quadrantPipe_bits_17 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  quadrantPipe_valid_18 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  quadrantPipe_bits_18 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  quadrantPipe_valid_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  quadrantPipe_bits_19 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  quadrantPipe_valid_20 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  quadrantPipe_bits_20 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  quadrantPipe_valid_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  quadrantPipe_bits_21 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  quadrantPipe_valid_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  quadrantPipe_bits_22 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  quadrantPipe_valid_23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  quadrantPipe_bits_23 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  quadrantPipe_valid_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  quadrantPipe_bits_24 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  quadrantPipe_valid_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  quadrantPipe_bits_25 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  quadrantPipe_valid_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  quadrantPipe_bits_26 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  quadrantPipe_valid_27 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  quadrantPipe_bits_27 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  quadrantPipe_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  quadrantPipe_bits_28 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  quadrantPipe_valid_29 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  quadrantPipe_bits_29 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  quadrantPipe_valid_30 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  quadrantPipe_bits_30 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  quadrantPipe_bits_31 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  trigonometric_io_theta_v = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  trigonometric_io_theta_b = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cosinePipe_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cosinePipe_bits = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sinePipe_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sinePipe_bits = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  signPipe_bits = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sqrt_log_io_uniform_v = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sqrt_log_io_uniform_b = _RAND_71[28:0];
  _RAND_72 = {1{`RANDOM}};
  sign_adjustedPipe_valid = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  sign_adjustedPipe_bits = _RAND_73[51:0];
  _RAND_74 = {1{`RANDOM}};
  io_g1_v = _RAND_74[0:0];
  _RAND_75 = {3{`RANDOM}};
  io_g1_b = _RAND_75[83:0];
  _RAND_76 = {1{`RANDOM}};
  io_g2_v = _RAND_76[0:0];
  _RAND_77 = {3{`RANDOM}};
  io_g2_b = _RAND_77[83:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MonteCarlo_10(
  input         clock,
  input         reset,
  output        io_request_0_ready,
  input         io_request_0_valid,
  input  [31:0] io_request_0_bits_time_steps,
  input  [31:0] io_request_0_bits_start_value,
  input  [31:0] io_request_0_bits_coefficient1,
  input  [31:0] io_request_0_bits_coefficient2,
  output        io_request_1_ready,
  input         io_request_1_valid,
  input  [31:0] io_request_1_bits_time_steps,
  input  [31:0] io_request_1_bits_start_value,
  input  [31:0] io_request_1_bits_coefficient1,
  input  [31:0] io_request_1_bits_coefficient2,
  input         io_response_0_ready,
  output        io_response_0_valid,
  output [31:0] io_response_0_bits,
  input         io_response_1_ready,
  output        io_response_1_valid,
  output [31:0] io_response_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rng_clock; // @[MonteCarlo.scala 42:19]
  wire  rng_reset; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g1_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g1_bits; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g2_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g2_bits; // @[MonteCarlo.scala 42:19]
  wire  initialized = rng_io_g1_valid & rng_io_g2_valid; // @[MonteCarlo.scala 47:37]
  reg [2:0] state; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_2 = $signed(io_request_0_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_3 = io_request_0_ready & io_request_0_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1; // @[Reg.scala 16:16]
  reg [31:0] c2; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_1 = io_request_0_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step; // @[Reg.scala 16:16]
  reg [31:0] price; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T = $signed(price) * $signed(c1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T = $signed(rng_io_g1_bits) * $signed(c2); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T = $signed(price) * $signed(partial_res2); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_2 = $signed(partial_res3) + $signed(partial_res1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_3 = counter == last_step ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_4 = counter == last_step ? counter : _counter_T_1; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_7 = io_response_0_ready & io_response_0_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_5 = _T_7 ? 3'h1 : state; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_6 = 3'h5 == state ? _GEN_5 : state; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_7 = 3'h4 == state ? $signed(_price_T_2) : $signed(price); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_3 : _GEN_6; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_9 = 3'h4 == state ? _GEN_4 : counter; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_64 = {$signed(partial_res3), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_10 = 3'h3 == state ? $signed(_partial_res3_T) : $signed({{12{_GEN_64[51]}},_GEN_64}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_11 = 3'h3 == state ? 3'h4 : _GEN_8; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_65 = {$signed(partial_res1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_14 = 3'h2 == state ? $signed(_partial_res1_T) : $signed({{12{_GEN_65[51]}},_GEN_65}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_66 = {$signed(partial_res2), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_15 = 3'h2 == state ? $signed(_partial_res2_T) : $signed({{20{_GEN_66[63]}},_GEN_66}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_17 = 3'h2 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_10); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_23 = 3'h1 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_14); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_24 = 3'h1 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_15); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_25 = 3'h1 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_17); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_29 = 3'h0 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_23); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_30 = 3'h0 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_24); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_31 = 3'h0 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_25); // @[MonteCarlo.scala 66:19 60:27]
  reg [2:0] state_1; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_6 = $signed(io_request_1_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_7 = io_request_1_ready & io_request_1_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1_1; // @[Reg.scala 16:16]
  reg [31:0] c2_1; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_4 = io_request_1_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step_1; // @[Reg.scala 16:16]
  reg [31:0] price_1; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1_1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2_1; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3_1; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter_1; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T_1 = $signed(price_1) * $signed(c1_1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T_1 = $signed(rng_io_g2_bits) * $signed(c2_1); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T_1 = $signed(price_1) * $signed(partial_res2_1); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_5 = $signed(partial_res3_1) + $signed(partial_res1_1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_35 = counter_1 == last_step_1 ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_36 = counter_1 == last_step_1 ? counter_1 : _counter_T_3; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_15 = io_response_1_ready & io_response_1_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_37 = _T_15 ? 3'h1 : state_1; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_38 = 3'h5 == state_1 ? _GEN_37 : state_1; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_39 = 3'h4 == state_1 ? $signed(_price_T_5) : $signed(price_1); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_40 = 3'h4 == state_1 ? _GEN_35 : _GEN_38; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_41 = 3'h4 == state_1 ? _GEN_36 : counter_1; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_74 = {$signed(partial_res3_1), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_42 = 3'h3 == state_1 ? $signed(_partial_res3_T_1) : $signed({{12{_GEN_74[51]}},_GEN_74}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_43 = 3'h3 == state_1 ? 3'h4 : _GEN_40; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_75 = {$signed(partial_res1_1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_46 = 3'h2 == state_1 ? $signed(_partial_res1_T_1) : $signed({{12{_GEN_75[51]}},_GEN_75}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_76 = {$signed(partial_res2_1), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_47 = 3'h2 == state_1 ? $signed(_partial_res2_T_1) : $signed({{20{_GEN_76[63]}},_GEN_76}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_49 = 3'h2 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_42); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_55 = 3'h1 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_46); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_56 = 3'h1 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_47); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_57 = 3'h1 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_49); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_61 = 3'h0 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_55); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_62 = 3'h0 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_56); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_63 = 3'h0 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_57); // @[MonteCarlo.scala 66:19 60:27]
  wire [43:0] _GEN_84 = _GEN_29[63:20];
  wire [51:0] _GEN_86 = _GEN_30[83:32];
  wire [43:0] _GEN_88 = _GEN_31[63:20];
  wire [43:0] _GEN_90 = _GEN_61[63:20];
  wire [51:0] _GEN_92 = _GEN_62[83:32];
  wire [43:0] _GEN_94 = _GEN_63[63:20];
  BoxMuller_10 rng ( // @[MonteCarlo.scala 42:19]
    .clock(rng_clock),
    .reset(rng_reset),
    .io_g1_valid(rng_io_g1_valid),
    .io_g1_bits(rng_io_g1_bits),
    .io_g2_valid(rng_io_g2_valid),
    .io_g2_bits(rng_io_g2_bits)
  );
  assign io_request_0_ready = state == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_request_1_ready = state_1 == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_response_0_valid = state == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_0_bits = price; // @[MonteCarlo.scala 65:16]
  assign io_response_1_valid = state_1 == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_1_bits = price_1; // @[MonteCarlo.scala 65:16]
  assign rng_clock = clock;
  assign rng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state <= 3'h1;
      end else begin
        state <= 3'h0;
      end
    end else if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_3) begin // @[MonteCarlo.scala 71:23]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[MonteCarlo.scala 66:19]
      state <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state <= _GEN_11;
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c1 <= _c1_T_2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c2 <= io_request_0_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      last_step <= _last_step_T_1; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        price <= io_request_0_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          price <= _GEN_7;
        end
      end
    end
    partial_res1 <= _GEN_84[31:0];
    partial_res2 <= _GEN_86[31:0];
    partial_res3 <= _GEN_88[31:0];
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        counter <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          counter <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state_1 <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state_1 <= 3'h1;
      end else begin
        state_1 <= 3'h0;
      end
    end else if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_7) begin // @[MonteCarlo.scala 71:23]
        state_1 <= 3'h2;
      end else begin
        state_1 <= 3'h1;
      end
    end else if (3'h2 == state_1) begin // @[MonteCarlo.scala 66:19]
      state_1 <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state_1 <= _GEN_43;
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c1_1 <= _c1_T_6; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c2_1 <= io_request_1_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      last_step_1 <= _last_step_T_4; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        price_1 <= io_request_1_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          price_1 <= _GEN_39;
        end
      end
    end
    partial_res1_1 <= _GEN_90[31:0];
    partial_res2_1 <= _GEN_92[31:0];
    partial_res3_1 <= _GEN_94[31:0];
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        counter_1 <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          counter_1 <= _GEN_41;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  c1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_step = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  price = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  partial_res1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  partial_res2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  partial_res3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  c1_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_step_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  price_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  partial_res1_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  partial_res2_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  partial_res3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  counter_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_22(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h92a85dd : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h16fc90ab : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h1da119db : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_23(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h118d439f : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h497df1 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h2aada8e4 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoxMuller_11(
  input         clock,
  input         reset,
  output        io_g1_valid,
  output [51:0] io_g1_bits,
  output        io_g2_valid,
  output [51:0] io_g2_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [95:0] _RAND_77;
`endif // RANDOMIZE_REG_INIT
  wire  rng1_clock; // @[BoxMuller.scala 51:20]
  wire  rng1_reset; // @[BoxMuller.scala 51:20]
  wire  rng1_io_rand_valid; // @[BoxMuller.scala 51:20]
  wire [31:0] rng1_io_rand_bits; // @[BoxMuller.scala 51:20]
  wire  rng2_clock; // @[BoxMuller.scala 52:20]
  wire  rng2_reset; // @[BoxMuller.scala 52:20]
  wire  rng2_io_rand_valid; // @[BoxMuller.scala 52:20]
  wire [31:0] rng2_io_rand_bits; // @[BoxMuller.scala 52:20]
  wire  trigonometric_clock; // @[BoxMuller.scala 55:29]
  wire  trigonometric_reset; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_theta_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_theta_bits; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_result_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_sine; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_cosine; // @[BoxMuller.scala 55:29]
  wire  sqrt_log_clock; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_reset; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_uniform_valid; // @[BoxMuller.scala 84:24]
  wire [31:0] sqrt_log_io_uniform_bits; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_result_valid; // @[BoxMuller.scala 84:24]
  wire [51:0] sqrt_log_io_result_bits; // @[BoxMuller.scala 84:24]
  wire [30:0] _theta_T_3 = {2'h0,rng1_io_rand_bits[28:0]}; // @[BoxMuller.scala 62:18]
  wire [62:0] _theta_T_4 = $signed(_theta_T_3) * 32'sh6487ed51; // @[BoxMuller.scala 62:26]
  reg  quadrantPipe_valid; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_1; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_1; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_2; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_2; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_3; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_3; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_4; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_4; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_5; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_5; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_6; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_6; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_7; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_7; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_8; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_8; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_9; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_9; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_10; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_10; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_11; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_11; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_12; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_12; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_13; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_13; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_14; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_14; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_15; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_15; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_16; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_16; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_17; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_17; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_18; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_18; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_19; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_19; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_20; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_20; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_21; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_21; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_22; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_22; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_23; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_23; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_24; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_24; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_25; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_25; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_26; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_26; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_27; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_27; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_28; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_28; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_29; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_29; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_30; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_30; // @[Reg.scala 16:16]
  reg [1:0] quadrantPipe_bits_31; // @[Reg.scala 16:16]
  reg  trigonometric_io_theta_v; // @[Valid.scala 127:22]
  reg [31:0] trigonometric_io_theta_b; // @[Reg.scala 16:16]
  wire [33:0] _GEN_40 = _theta_T_4[62:29]; // @[BoxMuller.scala 59:19 61:9]
  wire [31:0] theta = _GEN_40[31:0]; // @[BoxMuller.scala 59:19 61:9]
  wire  _cosine_T = quadrantPipe_bits_31 == 2'h0; // @[BoxMuller.scala 70:21]
  wire  _cosine_T_2 = quadrantPipe_bits_31 == 2'h0 | quadrantPipe_bits_31 == 2'h3; // @[BoxMuller.scala 70:29]
  wire [31:0] _cosine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_cosine); // @[BoxMuller.scala 72:7]
  reg  cosinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] cosinePipe_bits; // @[Reg.scala 16:16]
  wire  _sine_T_2 = _cosine_T | quadrantPipe_bits_31 == 2'h2; // @[BoxMuller.scala 78:29]
  wire [31:0] _sine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_sine); // @[BoxMuller.scala 80:7]
  reg  sinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] sinePipe_bits; // @[Reg.scala 16:16]
  reg  signPipe_bits; // @[Reg.scala 16:16]
  wire [28:0] _sqrt_log_io_uniform_T_1 = rng2_io_rand_bits[28:0]; // @[BoxMuller.scala 87:89]
  reg  sqrt_log_io_uniform_v; // @[Valid.scala 127:22]
  reg [28:0] sqrt_log_io_uniform_b; // @[Reg.scala 16:16]
  wire [51:0] _sign_adjusted_T_3 = 52'sh0 - $signed(sqrt_log_io_result_bits); // @[BoxMuller.scala 93:7]
  reg  sign_adjustedPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] sign_adjustedPipe_bits; // @[Reg.scala 16:16]
  wire  _io_g1_T = sign_adjustedPipe_valid & cosinePipe_valid; // @[BoxMuller.scala 99:25]
  wire [83:0] _io_g1_T_1 = $signed(cosinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 100:17]
  reg  io_g1_v; // @[Valid.scala 127:22]
  reg [83:0] io_g1_b; // @[Reg.scala 16:16]
  wire  _io_g2_T = sign_adjustedPipe_valid & sinePipe_valid; // @[BoxMuller.scala 103:25]
  wire [83:0] _io_g2_T_1 = $signed(sinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 104:15]
  reg  io_g2_v; // @[Valid.scala 127:22]
  reg [83:0] io_g2_b; // @[Reg.scala 16:16]
  wire [53:0] _GEN_42 = io_g1_b[83:30]; // @[BoxMuller.scala 98:9]
  wire [53:0] _GEN_44 = io_g2_b[83:30]; // @[BoxMuller.scala 102:9]
  wire [32:0] _GEN_46 = {$signed(trigonometric_io_theta_b), 1'h0}; // @[BoxMuller.scala 65:26]
  TauswortheUniform_22 rng1 ( // @[BoxMuller.scala 51:20]
    .clock(rng1_clock),
    .reset(rng1_reset),
    .io_rand_valid(rng1_io_rand_valid),
    .io_rand_bits(rng1_io_rand_bits)
  );
  TauswortheUniform_23 rng2 ( // @[BoxMuller.scala 52:20]
    .clock(rng2_clock),
    .reset(rng2_reset),
    .io_rand_valid(rng2_io_rand_valid),
    .io_rand_bits(rng2_io_rand_bits)
  );
  Trigonometric trigonometric ( // @[BoxMuller.scala 55:29]
    .clock(trigonometric_clock),
    .reset(trigonometric_reset),
    .io_theta_valid(trigonometric_io_theta_valid),
    .io_theta_bits(trigonometric_io_theta_bits),
    .io_result_valid(trigonometric_io_result_valid),
    .io_result_bits_sine(trigonometric_io_result_bits_sine),
    .io_result_bits_cosine(trigonometric_io_result_bits_cosine)
  );
  SquareRootLog sqrt_log ( // @[BoxMuller.scala 84:24]
    .clock(sqrt_log_clock),
    .reset(sqrt_log_reset),
    .io_uniform_valid(sqrt_log_io_uniform_valid),
    .io_uniform_bits(sqrt_log_io_uniform_bits),
    .io_result_valid(sqrt_log_io_result_valid),
    .io_result_bits(sqrt_log_io_result_bits)
  );
  assign io_g1_valid = io_g1_v; // @[Valid.scala 122:21 123:17]
  assign io_g1_bits = _GEN_42[51:0]; // @[BoxMuller.scala 98:9]
  assign io_g2_valid = io_g2_v; // @[Valid.scala 122:21 123:17]
  assign io_g2_bits = _GEN_44[51:0]; // @[BoxMuller.scala 102:9]
  assign rng1_clock = clock;
  assign rng1_reset = reset;
  assign rng2_clock = clock;
  assign rng2_reset = reset;
  assign trigonometric_clock = clock;
  assign trigonometric_reset = reset;
  assign trigonometric_io_theta_valid = trigonometric_io_theta_v; // @[Valid.scala 122:21 123:17]
  assign trigonometric_io_theta_bits = _GEN_46[31:0]; // @[BoxMuller.scala 65:26]
  assign sqrt_log_clock = clock;
  assign sqrt_log_reset = reset;
  assign sqrt_log_io_uniform_valid = sqrt_log_io_uniform_v; // @[Valid.scala 122:21 123:17]
  assign sqrt_log_io_uniform_bits = {{3{sqrt_log_io_uniform_b[28]}},sqrt_log_io_uniform_b}; // @[BoxMuller.scala 87:23]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits <= rng1_io_rand_bits[31:30]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_1 <= quadrantPipe_valid; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_1 <= quadrantPipe_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_2 <= quadrantPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_1) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_2 <= quadrantPipe_bits_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_3 <= quadrantPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_2) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_3 <= quadrantPipe_bits_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_4 <= quadrantPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_3) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_4 <= quadrantPipe_bits_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_5 <= quadrantPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_4) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_5 <= quadrantPipe_bits_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_6 <= quadrantPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_5) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_6 <= quadrantPipe_bits_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_7 <= quadrantPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_6) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_7 <= quadrantPipe_bits_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_8 <= quadrantPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_7) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_8 <= quadrantPipe_bits_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_9 <= quadrantPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_8) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_9 <= quadrantPipe_bits_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_10 <= quadrantPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_9) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_10 <= quadrantPipe_bits_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_11 <= quadrantPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_10) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_11 <= quadrantPipe_bits_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_12 <= quadrantPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_11) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_12 <= quadrantPipe_bits_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_13 <= quadrantPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_12) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_13 <= quadrantPipe_bits_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_14 <= quadrantPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_13) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_14 <= quadrantPipe_bits_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_15 <= quadrantPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_14) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_15 <= quadrantPipe_bits_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_16 <= quadrantPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_15) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_16 <= quadrantPipe_bits_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_17 <= quadrantPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_16) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_17 <= quadrantPipe_bits_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_18 <= quadrantPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_17) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_18 <= quadrantPipe_bits_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_19 <= quadrantPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_18) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_19 <= quadrantPipe_bits_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_20 <= quadrantPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_19) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_20 <= quadrantPipe_bits_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_21 <= quadrantPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_20) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_21 <= quadrantPipe_bits_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_22 <= quadrantPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_21) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_22 <= quadrantPipe_bits_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_23 <= quadrantPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_22) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_23 <= quadrantPipe_bits_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_24 <= quadrantPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_23) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_24 <= quadrantPipe_bits_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_25 <= quadrantPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_24) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_25 <= quadrantPipe_bits_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_26 <= quadrantPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_25) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_26 <= quadrantPipe_bits_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_27 <= quadrantPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_26) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_27 <= quadrantPipe_bits_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_28 <= quadrantPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_27) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_28 <= quadrantPipe_bits_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_29 <= quadrantPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_28) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_29 <= quadrantPipe_bits_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_30 <= quadrantPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_29) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_30 <= quadrantPipe_bits_29; // @[Reg.scala 17:22]
    end
    if (quadrantPipe_valid_30) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_31 <= quadrantPipe_bits_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      trigonometric_io_theta_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      trigonometric_io_theta_v <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      trigonometric_io_theta_b <= theta; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      cosinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      cosinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_cosine_T_2) begin // @[BoxMuller.scala 69:8]
        cosinePipe_bits <= trigonometric_io_result_bits_cosine;
      end else begin
        cosinePipe_bits <= _cosine_T_5;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      sinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_sine_T_2) begin // @[BoxMuller.scala 77:8]
        sinePipe_bits <= trigonometric_io_result_bits_sine;
      end else begin
        sinePipe_bits <= _sine_T_5;
      end
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      signPipe_bits <= rng2_io_rand_bits[31]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sqrt_log_io_uniform_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sqrt_log_io_uniform_v <= rng2_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      sqrt_log_io_uniform_b <= _sqrt_log_io_uniform_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sign_adjustedPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sign_adjustedPipe_valid <= sqrt_log_io_result_valid; // @[Valid.scala 127:22]
    end
    if (sqrt_log_io_result_valid) begin // @[Reg.scala 17:18]
      if (signPipe_bits) begin // @[BoxMuller.scala 91:8]
        sign_adjustedPipe_bits <= _sign_adjusted_T_3;
      end else begin
        sign_adjustedPipe_bits <= sqrt_log_io_result_bits;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g1_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g1_v <= _io_g1_T; // @[Valid.scala 127:22]
    end
    if (_io_g1_T) begin // @[Reg.scala 17:18]
      io_g1_b <= _io_g1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g2_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g2_v <= _io_g2_T; // @[Valid.scala 127:22]
    end
    if (_io_g2_T) begin // @[Reg.scala 17:18]
      io_g2_b <= _io_g2_T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quadrantPipe_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  quadrantPipe_bits = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  quadrantPipe_valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  quadrantPipe_bits_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  quadrantPipe_valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  quadrantPipe_bits_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  quadrantPipe_valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quadrantPipe_bits_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  quadrantPipe_valid_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  quadrantPipe_bits_4 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  quadrantPipe_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  quadrantPipe_bits_5 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  quadrantPipe_valid_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  quadrantPipe_bits_6 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  quadrantPipe_valid_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  quadrantPipe_bits_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  quadrantPipe_valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  quadrantPipe_bits_8 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  quadrantPipe_valid_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  quadrantPipe_bits_9 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  quadrantPipe_valid_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  quadrantPipe_bits_10 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  quadrantPipe_valid_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  quadrantPipe_bits_11 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  quadrantPipe_valid_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  quadrantPipe_bits_12 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  quadrantPipe_valid_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  quadrantPipe_bits_13 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  quadrantPipe_valid_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  quadrantPipe_bits_14 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  quadrantPipe_valid_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  quadrantPipe_bits_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  quadrantPipe_valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  quadrantPipe_bits_16 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  quadrantPipe_valid_17 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  quadrantPipe_bits_17 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  quadrantPipe_valid_18 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  quadrantPipe_bits_18 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  quadrantPipe_valid_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  quadrantPipe_bits_19 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  quadrantPipe_valid_20 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  quadrantPipe_bits_20 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  quadrantPipe_valid_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  quadrantPipe_bits_21 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  quadrantPipe_valid_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  quadrantPipe_bits_22 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  quadrantPipe_valid_23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  quadrantPipe_bits_23 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  quadrantPipe_valid_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  quadrantPipe_bits_24 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  quadrantPipe_valid_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  quadrantPipe_bits_25 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  quadrantPipe_valid_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  quadrantPipe_bits_26 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  quadrantPipe_valid_27 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  quadrantPipe_bits_27 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  quadrantPipe_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  quadrantPipe_bits_28 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  quadrantPipe_valid_29 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  quadrantPipe_bits_29 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  quadrantPipe_valid_30 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  quadrantPipe_bits_30 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  quadrantPipe_bits_31 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  trigonometric_io_theta_v = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  trigonometric_io_theta_b = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cosinePipe_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cosinePipe_bits = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sinePipe_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sinePipe_bits = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  signPipe_bits = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sqrt_log_io_uniform_v = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sqrt_log_io_uniform_b = _RAND_71[28:0];
  _RAND_72 = {1{`RANDOM}};
  sign_adjustedPipe_valid = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  sign_adjustedPipe_bits = _RAND_73[51:0];
  _RAND_74 = {1{`RANDOM}};
  io_g1_v = _RAND_74[0:0];
  _RAND_75 = {3{`RANDOM}};
  io_g1_b = _RAND_75[83:0];
  _RAND_76 = {1{`RANDOM}};
  io_g2_v = _RAND_76[0:0];
  _RAND_77 = {3{`RANDOM}};
  io_g2_b = _RAND_77[83:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MonteCarlo_11(
  input         clock,
  input         reset,
  output        io_request_0_ready,
  input         io_request_0_valid,
  input  [31:0] io_request_0_bits_time_steps,
  input  [31:0] io_request_0_bits_start_value,
  input  [31:0] io_request_0_bits_coefficient1,
  input  [31:0] io_request_0_bits_coefficient2,
  output        io_request_1_ready,
  input         io_request_1_valid,
  input  [31:0] io_request_1_bits_time_steps,
  input  [31:0] io_request_1_bits_start_value,
  input  [31:0] io_request_1_bits_coefficient1,
  input  [31:0] io_request_1_bits_coefficient2,
  input         io_response_0_ready,
  output        io_response_0_valid,
  output [31:0] io_response_0_bits,
  input         io_response_1_ready,
  output        io_response_1_valid,
  output [31:0] io_response_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rng_clock; // @[MonteCarlo.scala 42:19]
  wire  rng_reset; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g1_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g1_bits; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g2_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g2_bits; // @[MonteCarlo.scala 42:19]
  wire  initialized = rng_io_g1_valid & rng_io_g2_valid; // @[MonteCarlo.scala 47:37]
  reg [2:0] state; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_2 = $signed(io_request_0_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_3 = io_request_0_ready & io_request_0_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1; // @[Reg.scala 16:16]
  reg [31:0] c2; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_1 = io_request_0_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step; // @[Reg.scala 16:16]
  reg [31:0] price; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T = $signed(price) * $signed(c1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T = $signed(rng_io_g1_bits) * $signed(c2); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T = $signed(price) * $signed(partial_res2); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_2 = $signed(partial_res3) + $signed(partial_res1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_3 = counter == last_step ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_4 = counter == last_step ? counter : _counter_T_1; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_7 = io_response_0_ready & io_response_0_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_5 = _T_7 ? 3'h1 : state; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_6 = 3'h5 == state ? _GEN_5 : state; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_7 = 3'h4 == state ? $signed(_price_T_2) : $signed(price); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_3 : _GEN_6; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_9 = 3'h4 == state ? _GEN_4 : counter; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_64 = {$signed(partial_res3), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_10 = 3'h3 == state ? $signed(_partial_res3_T) : $signed({{12{_GEN_64[51]}},_GEN_64}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_11 = 3'h3 == state ? 3'h4 : _GEN_8; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_65 = {$signed(partial_res1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_14 = 3'h2 == state ? $signed(_partial_res1_T) : $signed({{12{_GEN_65[51]}},_GEN_65}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_66 = {$signed(partial_res2), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_15 = 3'h2 == state ? $signed(_partial_res2_T) : $signed({{20{_GEN_66[63]}},_GEN_66}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_17 = 3'h2 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_10); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_23 = 3'h1 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_14); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_24 = 3'h1 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_15); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_25 = 3'h1 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_17); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_29 = 3'h0 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_23); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_30 = 3'h0 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_24); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_31 = 3'h0 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_25); // @[MonteCarlo.scala 66:19 60:27]
  reg [2:0] state_1; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_6 = $signed(io_request_1_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_7 = io_request_1_ready & io_request_1_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1_1; // @[Reg.scala 16:16]
  reg [31:0] c2_1; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_4 = io_request_1_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step_1; // @[Reg.scala 16:16]
  reg [31:0] price_1; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1_1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2_1; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3_1; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter_1; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T_1 = $signed(price_1) * $signed(c1_1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T_1 = $signed(rng_io_g2_bits) * $signed(c2_1); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T_1 = $signed(price_1) * $signed(partial_res2_1); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_5 = $signed(partial_res3_1) + $signed(partial_res1_1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_35 = counter_1 == last_step_1 ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_36 = counter_1 == last_step_1 ? counter_1 : _counter_T_3; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_15 = io_response_1_ready & io_response_1_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_37 = _T_15 ? 3'h1 : state_1; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_38 = 3'h5 == state_1 ? _GEN_37 : state_1; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_39 = 3'h4 == state_1 ? $signed(_price_T_5) : $signed(price_1); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_40 = 3'h4 == state_1 ? _GEN_35 : _GEN_38; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_41 = 3'h4 == state_1 ? _GEN_36 : counter_1; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_74 = {$signed(partial_res3_1), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_42 = 3'h3 == state_1 ? $signed(_partial_res3_T_1) : $signed({{12{_GEN_74[51]}},_GEN_74}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_43 = 3'h3 == state_1 ? 3'h4 : _GEN_40; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_75 = {$signed(partial_res1_1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_46 = 3'h2 == state_1 ? $signed(_partial_res1_T_1) : $signed({{12{_GEN_75[51]}},_GEN_75}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_76 = {$signed(partial_res2_1), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_47 = 3'h2 == state_1 ? $signed(_partial_res2_T_1) : $signed({{20{_GEN_76[63]}},_GEN_76}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_49 = 3'h2 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_42); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_55 = 3'h1 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_46); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_56 = 3'h1 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_47); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_57 = 3'h1 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_49); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_61 = 3'h0 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_55); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_62 = 3'h0 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_56); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_63 = 3'h0 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_57); // @[MonteCarlo.scala 66:19 60:27]
  wire [43:0] _GEN_84 = _GEN_29[63:20];
  wire [51:0] _GEN_86 = _GEN_30[83:32];
  wire [43:0] _GEN_88 = _GEN_31[63:20];
  wire [43:0] _GEN_90 = _GEN_61[63:20];
  wire [51:0] _GEN_92 = _GEN_62[83:32];
  wire [43:0] _GEN_94 = _GEN_63[63:20];
  BoxMuller_11 rng ( // @[MonteCarlo.scala 42:19]
    .clock(rng_clock),
    .reset(rng_reset),
    .io_g1_valid(rng_io_g1_valid),
    .io_g1_bits(rng_io_g1_bits),
    .io_g2_valid(rng_io_g2_valid),
    .io_g2_bits(rng_io_g2_bits)
  );
  assign io_request_0_ready = state == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_request_1_ready = state_1 == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_response_0_valid = state == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_0_bits = price; // @[MonteCarlo.scala 65:16]
  assign io_response_1_valid = state_1 == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_1_bits = price_1; // @[MonteCarlo.scala 65:16]
  assign rng_clock = clock;
  assign rng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state <= 3'h1;
      end else begin
        state <= 3'h0;
      end
    end else if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_3) begin // @[MonteCarlo.scala 71:23]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[MonteCarlo.scala 66:19]
      state <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state <= _GEN_11;
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c1 <= _c1_T_2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c2 <= io_request_0_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      last_step <= _last_step_T_1; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        price <= io_request_0_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          price <= _GEN_7;
        end
      end
    end
    partial_res1 <= _GEN_84[31:0];
    partial_res2 <= _GEN_86[31:0];
    partial_res3 <= _GEN_88[31:0];
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        counter <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          counter <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state_1 <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state_1 <= 3'h1;
      end else begin
        state_1 <= 3'h0;
      end
    end else if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_7) begin // @[MonteCarlo.scala 71:23]
        state_1 <= 3'h2;
      end else begin
        state_1 <= 3'h1;
      end
    end else if (3'h2 == state_1) begin // @[MonteCarlo.scala 66:19]
      state_1 <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state_1 <= _GEN_43;
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c1_1 <= _c1_T_6; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c2_1 <= io_request_1_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      last_step_1 <= _last_step_T_4; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        price_1 <= io_request_1_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          price_1 <= _GEN_39;
        end
      end
    end
    partial_res1_1 <= _GEN_90[31:0];
    partial_res2_1 <= _GEN_92[31:0];
    partial_res3_1 <= _GEN_94[31:0];
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        counter_1 <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          counter_1 <= _GEN_41;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  c1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_step = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  price = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  partial_res1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  partial_res2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  partial_res3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  c1_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_step_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  price_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  partial_res1_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  partial_res2_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  partial_res3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  counter_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_24(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h4936da8 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h2c20d55b : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h164c8453 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_25(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h34385232 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h15ae66ec : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h26d03543 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoxMuller_12(
  input         clock,
  input         reset,
  output        io_g1_valid,
  output [51:0] io_g1_bits,
  output        io_g2_valid,
  output [51:0] io_g2_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [95:0] _RAND_77;
`endif // RANDOMIZE_REG_INIT
  wire  rng1_clock; // @[BoxMuller.scala 51:20]
  wire  rng1_reset; // @[BoxMuller.scala 51:20]
  wire  rng1_io_rand_valid; // @[BoxMuller.scala 51:20]
  wire [31:0] rng1_io_rand_bits; // @[BoxMuller.scala 51:20]
  wire  rng2_clock; // @[BoxMuller.scala 52:20]
  wire  rng2_reset; // @[BoxMuller.scala 52:20]
  wire  rng2_io_rand_valid; // @[BoxMuller.scala 52:20]
  wire [31:0] rng2_io_rand_bits; // @[BoxMuller.scala 52:20]
  wire  trigonometric_clock; // @[BoxMuller.scala 55:29]
  wire  trigonometric_reset; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_theta_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_theta_bits; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_result_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_sine; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_cosine; // @[BoxMuller.scala 55:29]
  wire  sqrt_log_clock; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_reset; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_uniform_valid; // @[BoxMuller.scala 84:24]
  wire [31:0] sqrt_log_io_uniform_bits; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_result_valid; // @[BoxMuller.scala 84:24]
  wire [51:0] sqrt_log_io_result_bits; // @[BoxMuller.scala 84:24]
  wire [30:0] _theta_T_3 = {2'h0,rng1_io_rand_bits[28:0]}; // @[BoxMuller.scala 62:18]
  wire [62:0] _theta_T_4 = $signed(_theta_T_3) * 32'sh6487ed51; // @[BoxMuller.scala 62:26]
  reg  quadrantPipe_valid; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_1; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_1; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_2; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_2; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_3; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_3; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_4; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_4; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_5; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_5; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_6; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_6; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_7; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_7; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_8; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_8; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_9; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_9; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_10; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_10; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_11; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_11; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_12; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_12; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_13; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_13; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_14; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_14; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_15; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_15; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_16; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_16; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_17; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_17; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_18; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_18; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_19; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_19; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_20; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_20; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_21; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_21; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_22; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_22; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_23; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_23; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_24; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_24; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_25; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_25; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_26; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_26; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_27; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_27; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_28; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_28; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_29; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_29; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_30; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_30; // @[Reg.scala 16:16]
  reg [1:0] quadrantPipe_bits_31; // @[Reg.scala 16:16]
  reg  trigonometric_io_theta_v; // @[Valid.scala 127:22]
  reg [31:0] trigonometric_io_theta_b; // @[Reg.scala 16:16]
  wire [33:0] _GEN_40 = _theta_T_4[62:29]; // @[BoxMuller.scala 59:19 61:9]
  wire [31:0] theta = _GEN_40[31:0]; // @[BoxMuller.scala 59:19 61:9]
  wire  _cosine_T = quadrantPipe_bits_31 == 2'h0; // @[BoxMuller.scala 70:21]
  wire  _cosine_T_2 = quadrantPipe_bits_31 == 2'h0 | quadrantPipe_bits_31 == 2'h3; // @[BoxMuller.scala 70:29]
  wire [31:0] _cosine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_cosine); // @[BoxMuller.scala 72:7]
  reg  cosinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] cosinePipe_bits; // @[Reg.scala 16:16]
  wire  _sine_T_2 = _cosine_T | quadrantPipe_bits_31 == 2'h2; // @[BoxMuller.scala 78:29]
  wire [31:0] _sine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_sine); // @[BoxMuller.scala 80:7]
  reg  sinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] sinePipe_bits; // @[Reg.scala 16:16]
  reg  signPipe_bits; // @[Reg.scala 16:16]
  wire [28:0] _sqrt_log_io_uniform_T_1 = rng2_io_rand_bits[28:0]; // @[BoxMuller.scala 87:89]
  reg  sqrt_log_io_uniform_v; // @[Valid.scala 127:22]
  reg [28:0] sqrt_log_io_uniform_b; // @[Reg.scala 16:16]
  wire [51:0] _sign_adjusted_T_3 = 52'sh0 - $signed(sqrt_log_io_result_bits); // @[BoxMuller.scala 93:7]
  reg  sign_adjustedPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] sign_adjustedPipe_bits; // @[Reg.scala 16:16]
  wire  _io_g1_T = sign_adjustedPipe_valid & cosinePipe_valid; // @[BoxMuller.scala 99:25]
  wire [83:0] _io_g1_T_1 = $signed(cosinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 100:17]
  reg  io_g1_v; // @[Valid.scala 127:22]
  reg [83:0] io_g1_b; // @[Reg.scala 16:16]
  wire  _io_g2_T = sign_adjustedPipe_valid & sinePipe_valid; // @[BoxMuller.scala 103:25]
  wire [83:0] _io_g2_T_1 = $signed(sinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 104:15]
  reg  io_g2_v; // @[Valid.scala 127:22]
  reg [83:0] io_g2_b; // @[Reg.scala 16:16]
  wire [53:0] _GEN_42 = io_g1_b[83:30]; // @[BoxMuller.scala 98:9]
  wire [53:0] _GEN_44 = io_g2_b[83:30]; // @[BoxMuller.scala 102:9]
  wire [32:0] _GEN_46 = {$signed(trigonometric_io_theta_b), 1'h0}; // @[BoxMuller.scala 65:26]
  TauswortheUniform_24 rng1 ( // @[BoxMuller.scala 51:20]
    .clock(rng1_clock),
    .reset(rng1_reset),
    .io_rand_valid(rng1_io_rand_valid),
    .io_rand_bits(rng1_io_rand_bits)
  );
  TauswortheUniform_25 rng2 ( // @[BoxMuller.scala 52:20]
    .clock(rng2_clock),
    .reset(rng2_reset),
    .io_rand_valid(rng2_io_rand_valid),
    .io_rand_bits(rng2_io_rand_bits)
  );
  Trigonometric trigonometric ( // @[BoxMuller.scala 55:29]
    .clock(trigonometric_clock),
    .reset(trigonometric_reset),
    .io_theta_valid(trigonometric_io_theta_valid),
    .io_theta_bits(trigonometric_io_theta_bits),
    .io_result_valid(trigonometric_io_result_valid),
    .io_result_bits_sine(trigonometric_io_result_bits_sine),
    .io_result_bits_cosine(trigonometric_io_result_bits_cosine)
  );
  SquareRootLog sqrt_log ( // @[BoxMuller.scala 84:24]
    .clock(sqrt_log_clock),
    .reset(sqrt_log_reset),
    .io_uniform_valid(sqrt_log_io_uniform_valid),
    .io_uniform_bits(sqrt_log_io_uniform_bits),
    .io_result_valid(sqrt_log_io_result_valid),
    .io_result_bits(sqrt_log_io_result_bits)
  );
  assign io_g1_valid = io_g1_v; // @[Valid.scala 122:21 123:17]
  assign io_g1_bits = _GEN_42[51:0]; // @[BoxMuller.scala 98:9]
  assign io_g2_valid = io_g2_v; // @[Valid.scala 122:21 123:17]
  assign io_g2_bits = _GEN_44[51:0]; // @[BoxMuller.scala 102:9]
  assign rng1_clock = clock;
  assign rng1_reset = reset;
  assign rng2_clock = clock;
  assign rng2_reset = reset;
  assign trigonometric_clock = clock;
  assign trigonometric_reset = reset;
  assign trigonometric_io_theta_valid = trigonometric_io_theta_v; // @[Valid.scala 122:21 123:17]
  assign trigonometric_io_theta_bits = _GEN_46[31:0]; // @[BoxMuller.scala 65:26]
  assign sqrt_log_clock = clock;
  assign sqrt_log_reset = reset;
  assign sqrt_log_io_uniform_valid = sqrt_log_io_uniform_v; // @[Valid.scala 122:21 123:17]
  assign sqrt_log_io_uniform_bits = {{3{sqrt_log_io_uniform_b[28]}},sqrt_log_io_uniform_b}; // @[BoxMuller.scala 87:23]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits <= rng1_io_rand_bits[31:30]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_1 <= quadrantPipe_valid; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_1 <= quadrantPipe_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_2 <= quadrantPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_1) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_2 <= quadrantPipe_bits_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_3 <= quadrantPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_2) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_3 <= quadrantPipe_bits_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_4 <= quadrantPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_3) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_4 <= quadrantPipe_bits_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_5 <= quadrantPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_4) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_5 <= quadrantPipe_bits_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_6 <= quadrantPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_5) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_6 <= quadrantPipe_bits_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_7 <= quadrantPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_6) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_7 <= quadrantPipe_bits_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_8 <= quadrantPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_7) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_8 <= quadrantPipe_bits_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_9 <= quadrantPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_8) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_9 <= quadrantPipe_bits_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_10 <= quadrantPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_9) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_10 <= quadrantPipe_bits_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_11 <= quadrantPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_10) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_11 <= quadrantPipe_bits_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_12 <= quadrantPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_11) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_12 <= quadrantPipe_bits_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_13 <= quadrantPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_12) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_13 <= quadrantPipe_bits_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_14 <= quadrantPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_13) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_14 <= quadrantPipe_bits_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_15 <= quadrantPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_14) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_15 <= quadrantPipe_bits_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_16 <= quadrantPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_15) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_16 <= quadrantPipe_bits_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_17 <= quadrantPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_16) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_17 <= quadrantPipe_bits_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_18 <= quadrantPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_17) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_18 <= quadrantPipe_bits_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_19 <= quadrantPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_18) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_19 <= quadrantPipe_bits_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_20 <= quadrantPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_19) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_20 <= quadrantPipe_bits_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_21 <= quadrantPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_20) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_21 <= quadrantPipe_bits_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_22 <= quadrantPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_21) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_22 <= quadrantPipe_bits_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_23 <= quadrantPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_22) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_23 <= quadrantPipe_bits_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_24 <= quadrantPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_23) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_24 <= quadrantPipe_bits_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_25 <= quadrantPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_24) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_25 <= quadrantPipe_bits_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_26 <= quadrantPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_25) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_26 <= quadrantPipe_bits_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_27 <= quadrantPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_26) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_27 <= quadrantPipe_bits_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_28 <= quadrantPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_27) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_28 <= quadrantPipe_bits_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_29 <= quadrantPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_28) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_29 <= quadrantPipe_bits_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_30 <= quadrantPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_29) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_30 <= quadrantPipe_bits_29; // @[Reg.scala 17:22]
    end
    if (quadrantPipe_valid_30) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_31 <= quadrantPipe_bits_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      trigonometric_io_theta_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      trigonometric_io_theta_v <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      trigonometric_io_theta_b <= theta; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      cosinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      cosinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_cosine_T_2) begin // @[BoxMuller.scala 69:8]
        cosinePipe_bits <= trigonometric_io_result_bits_cosine;
      end else begin
        cosinePipe_bits <= _cosine_T_5;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      sinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_sine_T_2) begin // @[BoxMuller.scala 77:8]
        sinePipe_bits <= trigonometric_io_result_bits_sine;
      end else begin
        sinePipe_bits <= _sine_T_5;
      end
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      signPipe_bits <= rng2_io_rand_bits[31]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sqrt_log_io_uniform_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sqrt_log_io_uniform_v <= rng2_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      sqrt_log_io_uniform_b <= _sqrt_log_io_uniform_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sign_adjustedPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sign_adjustedPipe_valid <= sqrt_log_io_result_valid; // @[Valid.scala 127:22]
    end
    if (sqrt_log_io_result_valid) begin // @[Reg.scala 17:18]
      if (signPipe_bits) begin // @[BoxMuller.scala 91:8]
        sign_adjustedPipe_bits <= _sign_adjusted_T_3;
      end else begin
        sign_adjustedPipe_bits <= sqrt_log_io_result_bits;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g1_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g1_v <= _io_g1_T; // @[Valid.scala 127:22]
    end
    if (_io_g1_T) begin // @[Reg.scala 17:18]
      io_g1_b <= _io_g1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g2_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g2_v <= _io_g2_T; // @[Valid.scala 127:22]
    end
    if (_io_g2_T) begin // @[Reg.scala 17:18]
      io_g2_b <= _io_g2_T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quadrantPipe_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  quadrantPipe_bits = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  quadrantPipe_valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  quadrantPipe_bits_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  quadrantPipe_valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  quadrantPipe_bits_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  quadrantPipe_valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quadrantPipe_bits_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  quadrantPipe_valid_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  quadrantPipe_bits_4 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  quadrantPipe_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  quadrantPipe_bits_5 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  quadrantPipe_valid_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  quadrantPipe_bits_6 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  quadrantPipe_valid_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  quadrantPipe_bits_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  quadrantPipe_valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  quadrantPipe_bits_8 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  quadrantPipe_valid_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  quadrantPipe_bits_9 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  quadrantPipe_valid_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  quadrantPipe_bits_10 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  quadrantPipe_valid_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  quadrantPipe_bits_11 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  quadrantPipe_valid_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  quadrantPipe_bits_12 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  quadrantPipe_valid_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  quadrantPipe_bits_13 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  quadrantPipe_valid_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  quadrantPipe_bits_14 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  quadrantPipe_valid_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  quadrantPipe_bits_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  quadrantPipe_valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  quadrantPipe_bits_16 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  quadrantPipe_valid_17 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  quadrantPipe_bits_17 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  quadrantPipe_valid_18 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  quadrantPipe_bits_18 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  quadrantPipe_valid_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  quadrantPipe_bits_19 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  quadrantPipe_valid_20 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  quadrantPipe_bits_20 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  quadrantPipe_valid_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  quadrantPipe_bits_21 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  quadrantPipe_valid_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  quadrantPipe_bits_22 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  quadrantPipe_valid_23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  quadrantPipe_bits_23 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  quadrantPipe_valid_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  quadrantPipe_bits_24 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  quadrantPipe_valid_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  quadrantPipe_bits_25 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  quadrantPipe_valid_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  quadrantPipe_bits_26 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  quadrantPipe_valid_27 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  quadrantPipe_bits_27 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  quadrantPipe_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  quadrantPipe_bits_28 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  quadrantPipe_valid_29 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  quadrantPipe_bits_29 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  quadrantPipe_valid_30 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  quadrantPipe_bits_30 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  quadrantPipe_bits_31 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  trigonometric_io_theta_v = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  trigonometric_io_theta_b = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cosinePipe_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cosinePipe_bits = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sinePipe_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sinePipe_bits = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  signPipe_bits = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sqrt_log_io_uniform_v = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sqrt_log_io_uniform_b = _RAND_71[28:0];
  _RAND_72 = {1{`RANDOM}};
  sign_adjustedPipe_valid = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  sign_adjustedPipe_bits = _RAND_73[51:0];
  _RAND_74 = {1{`RANDOM}};
  io_g1_v = _RAND_74[0:0];
  _RAND_75 = {3{`RANDOM}};
  io_g1_b = _RAND_75[83:0];
  _RAND_76 = {1{`RANDOM}};
  io_g2_v = _RAND_76[0:0];
  _RAND_77 = {3{`RANDOM}};
  io_g2_b = _RAND_77[83:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MonteCarlo_12(
  input         clock,
  input         reset,
  output        io_request_0_ready,
  input         io_request_0_valid,
  input  [31:0] io_request_0_bits_time_steps,
  input  [31:0] io_request_0_bits_start_value,
  input  [31:0] io_request_0_bits_coefficient1,
  input  [31:0] io_request_0_bits_coefficient2,
  output        io_request_1_ready,
  input         io_request_1_valid,
  input  [31:0] io_request_1_bits_time_steps,
  input  [31:0] io_request_1_bits_start_value,
  input  [31:0] io_request_1_bits_coefficient1,
  input  [31:0] io_request_1_bits_coefficient2,
  input         io_response_0_ready,
  output        io_response_0_valid,
  output [31:0] io_response_0_bits,
  input         io_response_1_ready,
  output        io_response_1_valid,
  output [31:0] io_response_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rng_clock; // @[MonteCarlo.scala 42:19]
  wire  rng_reset; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g1_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g1_bits; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g2_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g2_bits; // @[MonteCarlo.scala 42:19]
  wire  initialized = rng_io_g1_valid & rng_io_g2_valid; // @[MonteCarlo.scala 47:37]
  reg [2:0] state; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_2 = $signed(io_request_0_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_3 = io_request_0_ready & io_request_0_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1; // @[Reg.scala 16:16]
  reg [31:0] c2; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_1 = io_request_0_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step; // @[Reg.scala 16:16]
  reg [31:0] price; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T = $signed(price) * $signed(c1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T = $signed(rng_io_g1_bits) * $signed(c2); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T = $signed(price) * $signed(partial_res2); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_2 = $signed(partial_res3) + $signed(partial_res1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_3 = counter == last_step ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_4 = counter == last_step ? counter : _counter_T_1; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_7 = io_response_0_ready & io_response_0_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_5 = _T_7 ? 3'h1 : state; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_6 = 3'h5 == state ? _GEN_5 : state; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_7 = 3'h4 == state ? $signed(_price_T_2) : $signed(price); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_3 : _GEN_6; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_9 = 3'h4 == state ? _GEN_4 : counter; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_64 = {$signed(partial_res3), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_10 = 3'h3 == state ? $signed(_partial_res3_T) : $signed({{12{_GEN_64[51]}},_GEN_64}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_11 = 3'h3 == state ? 3'h4 : _GEN_8; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_65 = {$signed(partial_res1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_14 = 3'h2 == state ? $signed(_partial_res1_T) : $signed({{12{_GEN_65[51]}},_GEN_65}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_66 = {$signed(partial_res2), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_15 = 3'h2 == state ? $signed(_partial_res2_T) : $signed({{20{_GEN_66[63]}},_GEN_66}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_17 = 3'h2 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_10); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_23 = 3'h1 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_14); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_24 = 3'h1 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_15); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_25 = 3'h1 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_17); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_29 = 3'h0 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_23); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_30 = 3'h0 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_24); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_31 = 3'h0 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_25); // @[MonteCarlo.scala 66:19 60:27]
  reg [2:0] state_1; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_6 = $signed(io_request_1_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_7 = io_request_1_ready & io_request_1_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1_1; // @[Reg.scala 16:16]
  reg [31:0] c2_1; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_4 = io_request_1_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step_1; // @[Reg.scala 16:16]
  reg [31:0] price_1; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1_1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2_1; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3_1; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter_1; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T_1 = $signed(price_1) * $signed(c1_1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T_1 = $signed(rng_io_g2_bits) * $signed(c2_1); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T_1 = $signed(price_1) * $signed(partial_res2_1); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_5 = $signed(partial_res3_1) + $signed(partial_res1_1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_35 = counter_1 == last_step_1 ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_36 = counter_1 == last_step_1 ? counter_1 : _counter_T_3; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_15 = io_response_1_ready & io_response_1_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_37 = _T_15 ? 3'h1 : state_1; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_38 = 3'h5 == state_1 ? _GEN_37 : state_1; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_39 = 3'h4 == state_1 ? $signed(_price_T_5) : $signed(price_1); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_40 = 3'h4 == state_1 ? _GEN_35 : _GEN_38; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_41 = 3'h4 == state_1 ? _GEN_36 : counter_1; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_74 = {$signed(partial_res3_1), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_42 = 3'h3 == state_1 ? $signed(_partial_res3_T_1) : $signed({{12{_GEN_74[51]}},_GEN_74}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_43 = 3'h3 == state_1 ? 3'h4 : _GEN_40; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_75 = {$signed(partial_res1_1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_46 = 3'h2 == state_1 ? $signed(_partial_res1_T_1) : $signed({{12{_GEN_75[51]}},_GEN_75}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_76 = {$signed(partial_res2_1), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_47 = 3'h2 == state_1 ? $signed(_partial_res2_T_1) : $signed({{20{_GEN_76[63]}},_GEN_76}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_49 = 3'h2 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_42); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_55 = 3'h1 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_46); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_56 = 3'h1 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_47); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_57 = 3'h1 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_49); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_61 = 3'h0 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_55); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_62 = 3'h0 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_56); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_63 = 3'h0 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_57); // @[MonteCarlo.scala 66:19 60:27]
  wire [43:0] _GEN_84 = _GEN_29[63:20];
  wire [51:0] _GEN_86 = _GEN_30[83:32];
  wire [43:0] _GEN_88 = _GEN_31[63:20];
  wire [43:0] _GEN_90 = _GEN_61[63:20];
  wire [51:0] _GEN_92 = _GEN_62[83:32];
  wire [43:0] _GEN_94 = _GEN_63[63:20];
  BoxMuller_12 rng ( // @[MonteCarlo.scala 42:19]
    .clock(rng_clock),
    .reset(rng_reset),
    .io_g1_valid(rng_io_g1_valid),
    .io_g1_bits(rng_io_g1_bits),
    .io_g2_valid(rng_io_g2_valid),
    .io_g2_bits(rng_io_g2_bits)
  );
  assign io_request_0_ready = state == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_request_1_ready = state_1 == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_response_0_valid = state == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_0_bits = price; // @[MonteCarlo.scala 65:16]
  assign io_response_1_valid = state_1 == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_1_bits = price_1; // @[MonteCarlo.scala 65:16]
  assign rng_clock = clock;
  assign rng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state <= 3'h1;
      end else begin
        state <= 3'h0;
      end
    end else if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_3) begin // @[MonteCarlo.scala 71:23]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[MonteCarlo.scala 66:19]
      state <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state <= _GEN_11;
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c1 <= _c1_T_2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c2 <= io_request_0_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      last_step <= _last_step_T_1; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        price <= io_request_0_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          price <= _GEN_7;
        end
      end
    end
    partial_res1 <= _GEN_84[31:0];
    partial_res2 <= _GEN_86[31:0];
    partial_res3 <= _GEN_88[31:0];
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        counter <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          counter <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state_1 <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state_1 <= 3'h1;
      end else begin
        state_1 <= 3'h0;
      end
    end else if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_7) begin // @[MonteCarlo.scala 71:23]
        state_1 <= 3'h2;
      end else begin
        state_1 <= 3'h1;
      end
    end else if (3'h2 == state_1) begin // @[MonteCarlo.scala 66:19]
      state_1 <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state_1 <= _GEN_43;
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c1_1 <= _c1_T_6; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c2_1 <= io_request_1_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      last_step_1 <= _last_step_T_4; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        price_1 <= io_request_1_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          price_1 <= _GEN_39;
        end
      end
    end
    partial_res1_1 <= _GEN_90[31:0];
    partial_res2_1 <= _GEN_92[31:0];
    partial_res3_1 <= _GEN_94[31:0];
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        counter_1 <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          counter_1 <= _GEN_41;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  c1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_step = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  price = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  partial_res1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  partial_res2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  partial_res3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  c1_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_step_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  price_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  partial_res1_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  partial_res2_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  partial_res3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  counter_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_26(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h36ffb29b : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h3babeb32 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h3e2dd369 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_27(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h2fa537d6 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h37686166 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h222a80d2 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoxMuller_13(
  input         clock,
  input         reset,
  output        io_g1_valid,
  output [51:0] io_g1_bits,
  output        io_g2_valid,
  output [51:0] io_g2_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [95:0] _RAND_77;
`endif // RANDOMIZE_REG_INIT
  wire  rng1_clock; // @[BoxMuller.scala 51:20]
  wire  rng1_reset; // @[BoxMuller.scala 51:20]
  wire  rng1_io_rand_valid; // @[BoxMuller.scala 51:20]
  wire [31:0] rng1_io_rand_bits; // @[BoxMuller.scala 51:20]
  wire  rng2_clock; // @[BoxMuller.scala 52:20]
  wire  rng2_reset; // @[BoxMuller.scala 52:20]
  wire  rng2_io_rand_valid; // @[BoxMuller.scala 52:20]
  wire [31:0] rng2_io_rand_bits; // @[BoxMuller.scala 52:20]
  wire  trigonometric_clock; // @[BoxMuller.scala 55:29]
  wire  trigonometric_reset; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_theta_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_theta_bits; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_result_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_sine; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_cosine; // @[BoxMuller.scala 55:29]
  wire  sqrt_log_clock; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_reset; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_uniform_valid; // @[BoxMuller.scala 84:24]
  wire [31:0] sqrt_log_io_uniform_bits; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_result_valid; // @[BoxMuller.scala 84:24]
  wire [51:0] sqrt_log_io_result_bits; // @[BoxMuller.scala 84:24]
  wire [30:0] _theta_T_3 = {2'h0,rng1_io_rand_bits[28:0]}; // @[BoxMuller.scala 62:18]
  wire [62:0] _theta_T_4 = $signed(_theta_T_3) * 32'sh6487ed51; // @[BoxMuller.scala 62:26]
  reg  quadrantPipe_valid; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_1; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_1; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_2; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_2; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_3; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_3; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_4; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_4; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_5; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_5; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_6; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_6; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_7; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_7; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_8; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_8; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_9; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_9; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_10; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_10; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_11; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_11; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_12; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_12; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_13; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_13; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_14; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_14; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_15; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_15; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_16; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_16; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_17; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_17; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_18; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_18; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_19; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_19; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_20; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_20; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_21; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_21; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_22; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_22; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_23; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_23; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_24; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_24; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_25; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_25; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_26; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_26; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_27; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_27; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_28; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_28; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_29; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_29; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_30; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_30; // @[Reg.scala 16:16]
  reg [1:0] quadrantPipe_bits_31; // @[Reg.scala 16:16]
  reg  trigonometric_io_theta_v; // @[Valid.scala 127:22]
  reg [31:0] trigonometric_io_theta_b; // @[Reg.scala 16:16]
  wire [33:0] _GEN_40 = _theta_T_4[62:29]; // @[BoxMuller.scala 59:19 61:9]
  wire [31:0] theta = _GEN_40[31:0]; // @[BoxMuller.scala 59:19 61:9]
  wire  _cosine_T = quadrantPipe_bits_31 == 2'h0; // @[BoxMuller.scala 70:21]
  wire  _cosine_T_2 = quadrantPipe_bits_31 == 2'h0 | quadrantPipe_bits_31 == 2'h3; // @[BoxMuller.scala 70:29]
  wire [31:0] _cosine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_cosine); // @[BoxMuller.scala 72:7]
  reg  cosinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] cosinePipe_bits; // @[Reg.scala 16:16]
  wire  _sine_T_2 = _cosine_T | quadrantPipe_bits_31 == 2'h2; // @[BoxMuller.scala 78:29]
  wire [31:0] _sine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_sine); // @[BoxMuller.scala 80:7]
  reg  sinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] sinePipe_bits; // @[Reg.scala 16:16]
  reg  signPipe_bits; // @[Reg.scala 16:16]
  wire [28:0] _sqrt_log_io_uniform_T_1 = rng2_io_rand_bits[28:0]; // @[BoxMuller.scala 87:89]
  reg  sqrt_log_io_uniform_v; // @[Valid.scala 127:22]
  reg [28:0] sqrt_log_io_uniform_b; // @[Reg.scala 16:16]
  wire [51:0] _sign_adjusted_T_3 = 52'sh0 - $signed(sqrt_log_io_result_bits); // @[BoxMuller.scala 93:7]
  reg  sign_adjustedPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] sign_adjustedPipe_bits; // @[Reg.scala 16:16]
  wire  _io_g1_T = sign_adjustedPipe_valid & cosinePipe_valid; // @[BoxMuller.scala 99:25]
  wire [83:0] _io_g1_T_1 = $signed(cosinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 100:17]
  reg  io_g1_v; // @[Valid.scala 127:22]
  reg [83:0] io_g1_b; // @[Reg.scala 16:16]
  wire  _io_g2_T = sign_adjustedPipe_valid & sinePipe_valid; // @[BoxMuller.scala 103:25]
  wire [83:0] _io_g2_T_1 = $signed(sinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 104:15]
  reg  io_g2_v; // @[Valid.scala 127:22]
  reg [83:0] io_g2_b; // @[Reg.scala 16:16]
  wire [53:0] _GEN_42 = io_g1_b[83:30]; // @[BoxMuller.scala 98:9]
  wire [53:0] _GEN_44 = io_g2_b[83:30]; // @[BoxMuller.scala 102:9]
  wire [32:0] _GEN_46 = {$signed(trigonometric_io_theta_b), 1'h0}; // @[BoxMuller.scala 65:26]
  TauswortheUniform_26 rng1 ( // @[BoxMuller.scala 51:20]
    .clock(rng1_clock),
    .reset(rng1_reset),
    .io_rand_valid(rng1_io_rand_valid),
    .io_rand_bits(rng1_io_rand_bits)
  );
  TauswortheUniform_27 rng2 ( // @[BoxMuller.scala 52:20]
    .clock(rng2_clock),
    .reset(rng2_reset),
    .io_rand_valid(rng2_io_rand_valid),
    .io_rand_bits(rng2_io_rand_bits)
  );
  Trigonometric trigonometric ( // @[BoxMuller.scala 55:29]
    .clock(trigonometric_clock),
    .reset(trigonometric_reset),
    .io_theta_valid(trigonometric_io_theta_valid),
    .io_theta_bits(trigonometric_io_theta_bits),
    .io_result_valid(trigonometric_io_result_valid),
    .io_result_bits_sine(trigonometric_io_result_bits_sine),
    .io_result_bits_cosine(trigonometric_io_result_bits_cosine)
  );
  SquareRootLog sqrt_log ( // @[BoxMuller.scala 84:24]
    .clock(sqrt_log_clock),
    .reset(sqrt_log_reset),
    .io_uniform_valid(sqrt_log_io_uniform_valid),
    .io_uniform_bits(sqrt_log_io_uniform_bits),
    .io_result_valid(sqrt_log_io_result_valid),
    .io_result_bits(sqrt_log_io_result_bits)
  );
  assign io_g1_valid = io_g1_v; // @[Valid.scala 122:21 123:17]
  assign io_g1_bits = _GEN_42[51:0]; // @[BoxMuller.scala 98:9]
  assign io_g2_valid = io_g2_v; // @[Valid.scala 122:21 123:17]
  assign io_g2_bits = _GEN_44[51:0]; // @[BoxMuller.scala 102:9]
  assign rng1_clock = clock;
  assign rng1_reset = reset;
  assign rng2_clock = clock;
  assign rng2_reset = reset;
  assign trigonometric_clock = clock;
  assign trigonometric_reset = reset;
  assign trigonometric_io_theta_valid = trigonometric_io_theta_v; // @[Valid.scala 122:21 123:17]
  assign trigonometric_io_theta_bits = _GEN_46[31:0]; // @[BoxMuller.scala 65:26]
  assign sqrt_log_clock = clock;
  assign sqrt_log_reset = reset;
  assign sqrt_log_io_uniform_valid = sqrt_log_io_uniform_v; // @[Valid.scala 122:21 123:17]
  assign sqrt_log_io_uniform_bits = {{3{sqrt_log_io_uniform_b[28]}},sqrt_log_io_uniform_b}; // @[BoxMuller.scala 87:23]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits <= rng1_io_rand_bits[31:30]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_1 <= quadrantPipe_valid; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_1 <= quadrantPipe_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_2 <= quadrantPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_1) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_2 <= quadrantPipe_bits_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_3 <= quadrantPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_2) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_3 <= quadrantPipe_bits_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_4 <= quadrantPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_3) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_4 <= quadrantPipe_bits_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_5 <= quadrantPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_4) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_5 <= quadrantPipe_bits_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_6 <= quadrantPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_5) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_6 <= quadrantPipe_bits_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_7 <= quadrantPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_6) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_7 <= quadrantPipe_bits_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_8 <= quadrantPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_7) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_8 <= quadrantPipe_bits_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_9 <= quadrantPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_8) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_9 <= quadrantPipe_bits_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_10 <= quadrantPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_9) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_10 <= quadrantPipe_bits_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_11 <= quadrantPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_10) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_11 <= quadrantPipe_bits_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_12 <= quadrantPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_11) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_12 <= quadrantPipe_bits_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_13 <= quadrantPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_12) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_13 <= quadrantPipe_bits_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_14 <= quadrantPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_13) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_14 <= quadrantPipe_bits_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_15 <= quadrantPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_14) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_15 <= quadrantPipe_bits_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_16 <= quadrantPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_15) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_16 <= quadrantPipe_bits_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_17 <= quadrantPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_16) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_17 <= quadrantPipe_bits_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_18 <= quadrantPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_17) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_18 <= quadrantPipe_bits_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_19 <= quadrantPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_18) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_19 <= quadrantPipe_bits_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_20 <= quadrantPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_19) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_20 <= quadrantPipe_bits_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_21 <= quadrantPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_20) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_21 <= quadrantPipe_bits_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_22 <= quadrantPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_21) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_22 <= quadrantPipe_bits_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_23 <= quadrantPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_22) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_23 <= quadrantPipe_bits_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_24 <= quadrantPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_23) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_24 <= quadrantPipe_bits_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_25 <= quadrantPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_24) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_25 <= quadrantPipe_bits_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_26 <= quadrantPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_25) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_26 <= quadrantPipe_bits_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_27 <= quadrantPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_26) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_27 <= quadrantPipe_bits_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_28 <= quadrantPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_27) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_28 <= quadrantPipe_bits_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_29 <= quadrantPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_28) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_29 <= quadrantPipe_bits_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_30 <= quadrantPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_29) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_30 <= quadrantPipe_bits_29; // @[Reg.scala 17:22]
    end
    if (quadrantPipe_valid_30) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_31 <= quadrantPipe_bits_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      trigonometric_io_theta_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      trigonometric_io_theta_v <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      trigonometric_io_theta_b <= theta; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      cosinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      cosinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_cosine_T_2) begin // @[BoxMuller.scala 69:8]
        cosinePipe_bits <= trigonometric_io_result_bits_cosine;
      end else begin
        cosinePipe_bits <= _cosine_T_5;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      sinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_sine_T_2) begin // @[BoxMuller.scala 77:8]
        sinePipe_bits <= trigonometric_io_result_bits_sine;
      end else begin
        sinePipe_bits <= _sine_T_5;
      end
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      signPipe_bits <= rng2_io_rand_bits[31]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sqrt_log_io_uniform_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sqrt_log_io_uniform_v <= rng2_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      sqrt_log_io_uniform_b <= _sqrt_log_io_uniform_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sign_adjustedPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sign_adjustedPipe_valid <= sqrt_log_io_result_valid; // @[Valid.scala 127:22]
    end
    if (sqrt_log_io_result_valid) begin // @[Reg.scala 17:18]
      if (signPipe_bits) begin // @[BoxMuller.scala 91:8]
        sign_adjustedPipe_bits <= _sign_adjusted_T_3;
      end else begin
        sign_adjustedPipe_bits <= sqrt_log_io_result_bits;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g1_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g1_v <= _io_g1_T; // @[Valid.scala 127:22]
    end
    if (_io_g1_T) begin // @[Reg.scala 17:18]
      io_g1_b <= _io_g1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g2_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g2_v <= _io_g2_T; // @[Valid.scala 127:22]
    end
    if (_io_g2_T) begin // @[Reg.scala 17:18]
      io_g2_b <= _io_g2_T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quadrantPipe_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  quadrantPipe_bits = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  quadrantPipe_valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  quadrantPipe_bits_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  quadrantPipe_valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  quadrantPipe_bits_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  quadrantPipe_valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quadrantPipe_bits_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  quadrantPipe_valid_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  quadrantPipe_bits_4 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  quadrantPipe_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  quadrantPipe_bits_5 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  quadrantPipe_valid_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  quadrantPipe_bits_6 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  quadrantPipe_valid_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  quadrantPipe_bits_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  quadrantPipe_valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  quadrantPipe_bits_8 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  quadrantPipe_valid_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  quadrantPipe_bits_9 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  quadrantPipe_valid_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  quadrantPipe_bits_10 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  quadrantPipe_valid_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  quadrantPipe_bits_11 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  quadrantPipe_valid_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  quadrantPipe_bits_12 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  quadrantPipe_valid_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  quadrantPipe_bits_13 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  quadrantPipe_valid_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  quadrantPipe_bits_14 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  quadrantPipe_valid_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  quadrantPipe_bits_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  quadrantPipe_valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  quadrantPipe_bits_16 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  quadrantPipe_valid_17 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  quadrantPipe_bits_17 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  quadrantPipe_valid_18 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  quadrantPipe_bits_18 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  quadrantPipe_valid_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  quadrantPipe_bits_19 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  quadrantPipe_valid_20 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  quadrantPipe_bits_20 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  quadrantPipe_valid_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  quadrantPipe_bits_21 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  quadrantPipe_valid_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  quadrantPipe_bits_22 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  quadrantPipe_valid_23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  quadrantPipe_bits_23 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  quadrantPipe_valid_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  quadrantPipe_bits_24 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  quadrantPipe_valid_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  quadrantPipe_bits_25 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  quadrantPipe_valid_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  quadrantPipe_bits_26 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  quadrantPipe_valid_27 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  quadrantPipe_bits_27 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  quadrantPipe_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  quadrantPipe_bits_28 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  quadrantPipe_valid_29 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  quadrantPipe_bits_29 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  quadrantPipe_valid_30 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  quadrantPipe_bits_30 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  quadrantPipe_bits_31 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  trigonometric_io_theta_v = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  trigonometric_io_theta_b = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cosinePipe_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cosinePipe_bits = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sinePipe_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sinePipe_bits = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  signPipe_bits = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sqrt_log_io_uniform_v = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sqrt_log_io_uniform_b = _RAND_71[28:0];
  _RAND_72 = {1{`RANDOM}};
  sign_adjustedPipe_valid = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  sign_adjustedPipe_bits = _RAND_73[51:0];
  _RAND_74 = {1{`RANDOM}};
  io_g1_v = _RAND_74[0:0];
  _RAND_75 = {3{`RANDOM}};
  io_g1_b = _RAND_75[83:0];
  _RAND_76 = {1{`RANDOM}};
  io_g2_v = _RAND_76[0:0];
  _RAND_77 = {3{`RANDOM}};
  io_g2_b = _RAND_77[83:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MonteCarlo_13(
  input         clock,
  input         reset,
  output        io_request_0_ready,
  input         io_request_0_valid,
  input  [31:0] io_request_0_bits_time_steps,
  input  [31:0] io_request_0_bits_start_value,
  input  [31:0] io_request_0_bits_coefficient1,
  input  [31:0] io_request_0_bits_coefficient2,
  output        io_request_1_ready,
  input         io_request_1_valid,
  input  [31:0] io_request_1_bits_time_steps,
  input  [31:0] io_request_1_bits_start_value,
  input  [31:0] io_request_1_bits_coefficient1,
  input  [31:0] io_request_1_bits_coefficient2,
  input         io_response_0_ready,
  output        io_response_0_valid,
  output [31:0] io_response_0_bits,
  input         io_response_1_ready,
  output        io_response_1_valid,
  output [31:0] io_response_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rng_clock; // @[MonteCarlo.scala 42:19]
  wire  rng_reset; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g1_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g1_bits; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g2_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g2_bits; // @[MonteCarlo.scala 42:19]
  wire  initialized = rng_io_g1_valid & rng_io_g2_valid; // @[MonteCarlo.scala 47:37]
  reg [2:0] state; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_2 = $signed(io_request_0_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_3 = io_request_0_ready & io_request_0_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1; // @[Reg.scala 16:16]
  reg [31:0] c2; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_1 = io_request_0_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step; // @[Reg.scala 16:16]
  reg [31:0] price; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T = $signed(price) * $signed(c1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T = $signed(rng_io_g1_bits) * $signed(c2); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T = $signed(price) * $signed(partial_res2); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_2 = $signed(partial_res3) + $signed(partial_res1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_3 = counter == last_step ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_4 = counter == last_step ? counter : _counter_T_1; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_7 = io_response_0_ready & io_response_0_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_5 = _T_7 ? 3'h1 : state; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_6 = 3'h5 == state ? _GEN_5 : state; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_7 = 3'h4 == state ? $signed(_price_T_2) : $signed(price); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_3 : _GEN_6; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_9 = 3'h4 == state ? _GEN_4 : counter; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_64 = {$signed(partial_res3), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_10 = 3'h3 == state ? $signed(_partial_res3_T) : $signed({{12{_GEN_64[51]}},_GEN_64}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_11 = 3'h3 == state ? 3'h4 : _GEN_8; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_65 = {$signed(partial_res1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_14 = 3'h2 == state ? $signed(_partial_res1_T) : $signed({{12{_GEN_65[51]}},_GEN_65}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_66 = {$signed(partial_res2), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_15 = 3'h2 == state ? $signed(_partial_res2_T) : $signed({{20{_GEN_66[63]}},_GEN_66}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_17 = 3'h2 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_10); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_23 = 3'h1 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_14); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_24 = 3'h1 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_15); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_25 = 3'h1 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_17); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_29 = 3'h0 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_23); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_30 = 3'h0 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_24); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_31 = 3'h0 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_25); // @[MonteCarlo.scala 66:19 60:27]
  reg [2:0] state_1; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_6 = $signed(io_request_1_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_7 = io_request_1_ready & io_request_1_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1_1; // @[Reg.scala 16:16]
  reg [31:0] c2_1; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_4 = io_request_1_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step_1; // @[Reg.scala 16:16]
  reg [31:0] price_1; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1_1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2_1; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3_1; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter_1; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T_1 = $signed(price_1) * $signed(c1_1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T_1 = $signed(rng_io_g2_bits) * $signed(c2_1); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T_1 = $signed(price_1) * $signed(partial_res2_1); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_5 = $signed(partial_res3_1) + $signed(partial_res1_1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_35 = counter_1 == last_step_1 ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_36 = counter_1 == last_step_1 ? counter_1 : _counter_T_3; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_15 = io_response_1_ready & io_response_1_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_37 = _T_15 ? 3'h1 : state_1; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_38 = 3'h5 == state_1 ? _GEN_37 : state_1; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_39 = 3'h4 == state_1 ? $signed(_price_T_5) : $signed(price_1); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_40 = 3'h4 == state_1 ? _GEN_35 : _GEN_38; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_41 = 3'h4 == state_1 ? _GEN_36 : counter_1; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_74 = {$signed(partial_res3_1), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_42 = 3'h3 == state_1 ? $signed(_partial_res3_T_1) : $signed({{12{_GEN_74[51]}},_GEN_74}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_43 = 3'h3 == state_1 ? 3'h4 : _GEN_40; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_75 = {$signed(partial_res1_1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_46 = 3'h2 == state_1 ? $signed(_partial_res1_T_1) : $signed({{12{_GEN_75[51]}},_GEN_75}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_76 = {$signed(partial_res2_1), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_47 = 3'h2 == state_1 ? $signed(_partial_res2_T_1) : $signed({{20{_GEN_76[63]}},_GEN_76}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_49 = 3'h2 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_42); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_55 = 3'h1 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_46); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_56 = 3'h1 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_47); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_57 = 3'h1 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_49); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_61 = 3'h0 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_55); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_62 = 3'h0 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_56); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_63 = 3'h0 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_57); // @[MonteCarlo.scala 66:19 60:27]
  wire [43:0] _GEN_84 = _GEN_29[63:20];
  wire [51:0] _GEN_86 = _GEN_30[83:32];
  wire [43:0] _GEN_88 = _GEN_31[63:20];
  wire [43:0] _GEN_90 = _GEN_61[63:20];
  wire [51:0] _GEN_92 = _GEN_62[83:32];
  wire [43:0] _GEN_94 = _GEN_63[63:20];
  BoxMuller_13 rng ( // @[MonteCarlo.scala 42:19]
    .clock(rng_clock),
    .reset(rng_reset),
    .io_g1_valid(rng_io_g1_valid),
    .io_g1_bits(rng_io_g1_bits),
    .io_g2_valid(rng_io_g2_valid),
    .io_g2_bits(rng_io_g2_bits)
  );
  assign io_request_0_ready = state == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_request_1_ready = state_1 == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_response_0_valid = state == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_0_bits = price; // @[MonteCarlo.scala 65:16]
  assign io_response_1_valid = state_1 == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_1_bits = price_1; // @[MonteCarlo.scala 65:16]
  assign rng_clock = clock;
  assign rng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state <= 3'h1;
      end else begin
        state <= 3'h0;
      end
    end else if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_3) begin // @[MonteCarlo.scala 71:23]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[MonteCarlo.scala 66:19]
      state <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state <= _GEN_11;
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c1 <= _c1_T_2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c2 <= io_request_0_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      last_step <= _last_step_T_1; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        price <= io_request_0_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          price <= _GEN_7;
        end
      end
    end
    partial_res1 <= _GEN_84[31:0];
    partial_res2 <= _GEN_86[31:0];
    partial_res3 <= _GEN_88[31:0];
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        counter <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          counter <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state_1 <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state_1 <= 3'h1;
      end else begin
        state_1 <= 3'h0;
      end
    end else if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_7) begin // @[MonteCarlo.scala 71:23]
        state_1 <= 3'h2;
      end else begin
        state_1 <= 3'h1;
      end
    end else if (3'h2 == state_1) begin // @[MonteCarlo.scala 66:19]
      state_1 <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state_1 <= _GEN_43;
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c1_1 <= _c1_T_6; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c2_1 <= io_request_1_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      last_step_1 <= _last_step_T_4; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        price_1 <= io_request_1_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          price_1 <= _GEN_39;
        end
      end
    end
    partial_res1_1 <= _GEN_90[31:0];
    partial_res2_1 <= _GEN_92[31:0];
    partial_res3_1 <= _GEN_94[31:0];
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        counter_1 <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          counter_1 <= _GEN_41;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  c1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_step = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  price = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  partial_res1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  partial_res2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  partial_res3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  c1_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_step_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  price_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  partial_res1_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  partial_res2_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  partial_res3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  counter_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_28(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h27348760 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h2e05e10 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'hb748a0e : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_29(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h13eda019 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'hdecac72 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'hd049130 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoxMuller_14(
  input         clock,
  input         reset,
  output        io_g1_valid,
  output [51:0] io_g1_bits,
  output        io_g2_valid,
  output [51:0] io_g2_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [95:0] _RAND_77;
`endif // RANDOMIZE_REG_INIT
  wire  rng1_clock; // @[BoxMuller.scala 51:20]
  wire  rng1_reset; // @[BoxMuller.scala 51:20]
  wire  rng1_io_rand_valid; // @[BoxMuller.scala 51:20]
  wire [31:0] rng1_io_rand_bits; // @[BoxMuller.scala 51:20]
  wire  rng2_clock; // @[BoxMuller.scala 52:20]
  wire  rng2_reset; // @[BoxMuller.scala 52:20]
  wire  rng2_io_rand_valid; // @[BoxMuller.scala 52:20]
  wire [31:0] rng2_io_rand_bits; // @[BoxMuller.scala 52:20]
  wire  trigonometric_clock; // @[BoxMuller.scala 55:29]
  wire  trigonometric_reset; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_theta_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_theta_bits; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_result_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_sine; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_cosine; // @[BoxMuller.scala 55:29]
  wire  sqrt_log_clock; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_reset; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_uniform_valid; // @[BoxMuller.scala 84:24]
  wire [31:0] sqrt_log_io_uniform_bits; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_result_valid; // @[BoxMuller.scala 84:24]
  wire [51:0] sqrt_log_io_result_bits; // @[BoxMuller.scala 84:24]
  wire [30:0] _theta_T_3 = {2'h0,rng1_io_rand_bits[28:0]}; // @[BoxMuller.scala 62:18]
  wire [62:0] _theta_T_4 = $signed(_theta_T_3) * 32'sh6487ed51; // @[BoxMuller.scala 62:26]
  reg  quadrantPipe_valid; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_1; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_1; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_2; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_2; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_3; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_3; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_4; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_4; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_5; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_5; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_6; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_6; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_7; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_7; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_8; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_8; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_9; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_9; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_10; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_10; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_11; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_11; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_12; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_12; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_13; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_13; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_14; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_14; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_15; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_15; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_16; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_16; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_17; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_17; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_18; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_18; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_19; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_19; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_20; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_20; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_21; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_21; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_22; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_22; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_23; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_23; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_24; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_24; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_25; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_25; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_26; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_26; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_27; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_27; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_28; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_28; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_29; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_29; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_30; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_30; // @[Reg.scala 16:16]
  reg [1:0] quadrantPipe_bits_31; // @[Reg.scala 16:16]
  reg  trigonometric_io_theta_v; // @[Valid.scala 127:22]
  reg [31:0] trigonometric_io_theta_b; // @[Reg.scala 16:16]
  wire [33:0] _GEN_40 = _theta_T_4[62:29]; // @[BoxMuller.scala 59:19 61:9]
  wire [31:0] theta = _GEN_40[31:0]; // @[BoxMuller.scala 59:19 61:9]
  wire  _cosine_T = quadrantPipe_bits_31 == 2'h0; // @[BoxMuller.scala 70:21]
  wire  _cosine_T_2 = quadrantPipe_bits_31 == 2'h0 | quadrantPipe_bits_31 == 2'h3; // @[BoxMuller.scala 70:29]
  wire [31:0] _cosine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_cosine); // @[BoxMuller.scala 72:7]
  reg  cosinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] cosinePipe_bits; // @[Reg.scala 16:16]
  wire  _sine_T_2 = _cosine_T | quadrantPipe_bits_31 == 2'h2; // @[BoxMuller.scala 78:29]
  wire [31:0] _sine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_sine); // @[BoxMuller.scala 80:7]
  reg  sinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] sinePipe_bits; // @[Reg.scala 16:16]
  reg  signPipe_bits; // @[Reg.scala 16:16]
  wire [28:0] _sqrt_log_io_uniform_T_1 = rng2_io_rand_bits[28:0]; // @[BoxMuller.scala 87:89]
  reg  sqrt_log_io_uniform_v; // @[Valid.scala 127:22]
  reg [28:0] sqrt_log_io_uniform_b; // @[Reg.scala 16:16]
  wire [51:0] _sign_adjusted_T_3 = 52'sh0 - $signed(sqrt_log_io_result_bits); // @[BoxMuller.scala 93:7]
  reg  sign_adjustedPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] sign_adjustedPipe_bits; // @[Reg.scala 16:16]
  wire  _io_g1_T = sign_adjustedPipe_valid & cosinePipe_valid; // @[BoxMuller.scala 99:25]
  wire [83:0] _io_g1_T_1 = $signed(cosinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 100:17]
  reg  io_g1_v; // @[Valid.scala 127:22]
  reg [83:0] io_g1_b; // @[Reg.scala 16:16]
  wire  _io_g2_T = sign_adjustedPipe_valid & sinePipe_valid; // @[BoxMuller.scala 103:25]
  wire [83:0] _io_g2_T_1 = $signed(sinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 104:15]
  reg  io_g2_v; // @[Valid.scala 127:22]
  reg [83:0] io_g2_b; // @[Reg.scala 16:16]
  wire [53:0] _GEN_42 = io_g1_b[83:30]; // @[BoxMuller.scala 98:9]
  wire [53:0] _GEN_44 = io_g2_b[83:30]; // @[BoxMuller.scala 102:9]
  wire [32:0] _GEN_46 = {$signed(trigonometric_io_theta_b), 1'h0}; // @[BoxMuller.scala 65:26]
  TauswortheUniform_28 rng1 ( // @[BoxMuller.scala 51:20]
    .clock(rng1_clock),
    .reset(rng1_reset),
    .io_rand_valid(rng1_io_rand_valid),
    .io_rand_bits(rng1_io_rand_bits)
  );
  TauswortheUniform_29 rng2 ( // @[BoxMuller.scala 52:20]
    .clock(rng2_clock),
    .reset(rng2_reset),
    .io_rand_valid(rng2_io_rand_valid),
    .io_rand_bits(rng2_io_rand_bits)
  );
  Trigonometric trigonometric ( // @[BoxMuller.scala 55:29]
    .clock(trigonometric_clock),
    .reset(trigonometric_reset),
    .io_theta_valid(trigonometric_io_theta_valid),
    .io_theta_bits(trigonometric_io_theta_bits),
    .io_result_valid(trigonometric_io_result_valid),
    .io_result_bits_sine(trigonometric_io_result_bits_sine),
    .io_result_bits_cosine(trigonometric_io_result_bits_cosine)
  );
  SquareRootLog sqrt_log ( // @[BoxMuller.scala 84:24]
    .clock(sqrt_log_clock),
    .reset(sqrt_log_reset),
    .io_uniform_valid(sqrt_log_io_uniform_valid),
    .io_uniform_bits(sqrt_log_io_uniform_bits),
    .io_result_valid(sqrt_log_io_result_valid),
    .io_result_bits(sqrt_log_io_result_bits)
  );
  assign io_g1_valid = io_g1_v; // @[Valid.scala 122:21 123:17]
  assign io_g1_bits = _GEN_42[51:0]; // @[BoxMuller.scala 98:9]
  assign io_g2_valid = io_g2_v; // @[Valid.scala 122:21 123:17]
  assign io_g2_bits = _GEN_44[51:0]; // @[BoxMuller.scala 102:9]
  assign rng1_clock = clock;
  assign rng1_reset = reset;
  assign rng2_clock = clock;
  assign rng2_reset = reset;
  assign trigonometric_clock = clock;
  assign trigonometric_reset = reset;
  assign trigonometric_io_theta_valid = trigonometric_io_theta_v; // @[Valid.scala 122:21 123:17]
  assign trigonometric_io_theta_bits = _GEN_46[31:0]; // @[BoxMuller.scala 65:26]
  assign sqrt_log_clock = clock;
  assign sqrt_log_reset = reset;
  assign sqrt_log_io_uniform_valid = sqrt_log_io_uniform_v; // @[Valid.scala 122:21 123:17]
  assign sqrt_log_io_uniform_bits = {{3{sqrt_log_io_uniform_b[28]}},sqrt_log_io_uniform_b}; // @[BoxMuller.scala 87:23]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits <= rng1_io_rand_bits[31:30]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_1 <= quadrantPipe_valid; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_1 <= quadrantPipe_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_2 <= quadrantPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_1) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_2 <= quadrantPipe_bits_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_3 <= quadrantPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_2) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_3 <= quadrantPipe_bits_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_4 <= quadrantPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_3) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_4 <= quadrantPipe_bits_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_5 <= quadrantPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_4) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_5 <= quadrantPipe_bits_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_6 <= quadrantPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_5) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_6 <= quadrantPipe_bits_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_7 <= quadrantPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_6) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_7 <= quadrantPipe_bits_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_8 <= quadrantPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_7) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_8 <= quadrantPipe_bits_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_9 <= quadrantPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_8) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_9 <= quadrantPipe_bits_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_10 <= quadrantPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_9) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_10 <= quadrantPipe_bits_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_11 <= quadrantPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_10) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_11 <= quadrantPipe_bits_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_12 <= quadrantPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_11) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_12 <= quadrantPipe_bits_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_13 <= quadrantPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_12) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_13 <= quadrantPipe_bits_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_14 <= quadrantPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_13) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_14 <= quadrantPipe_bits_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_15 <= quadrantPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_14) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_15 <= quadrantPipe_bits_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_16 <= quadrantPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_15) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_16 <= quadrantPipe_bits_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_17 <= quadrantPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_16) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_17 <= quadrantPipe_bits_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_18 <= quadrantPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_17) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_18 <= quadrantPipe_bits_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_19 <= quadrantPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_18) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_19 <= quadrantPipe_bits_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_20 <= quadrantPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_19) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_20 <= quadrantPipe_bits_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_21 <= quadrantPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_20) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_21 <= quadrantPipe_bits_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_22 <= quadrantPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_21) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_22 <= quadrantPipe_bits_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_23 <= quadrantPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_22) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_23 <= quadrantPipe_bits_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_24 <= quadrantPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_23) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_24 <= quadrantPipe_bits_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_25 <= quadrantPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_24) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_25 <= quadrantPipe_bits_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_26 <= quadrantPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_25) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_26 <= quadrantPipe_bits_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_27 <= quadrantPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_26) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_27 <= quadrantPipe_bits_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_28 <= quadrantPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_27) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_28 <= quadrantPipe_bits_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_29 <= quadrantPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_28) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_29 <= quadrantPipe_bits_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_30 <= quadrantPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_29) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_30 <= quadrantPipe_bits_29; // @[Reg.scala 17:22]
    end
    if (quadrantPipe_valid_30) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_31 <= quadrantPipe_bits_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      trigonometric_io_theta_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      trigonometric_io_theta_v <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      trigonometric_io_theta_b <= theta; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      cosinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      cosinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_cosine_T_2) begin // @[BoxMuller.scala 69:8]
        cosinePipe_bits <= trigonometric_io_result_bits_cosine;
      end else begin
        cosinePipe_bits <= _cosine_T_5;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      sinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_sine_T_2) begin // @[BoxMuller.scala 77:8]
        sinePipe_bits <= trigonometric_io_result_bits_sine;
      end else begin
        sinePipe_bits <= _sine_T_5;
      end
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      signPipe_bits <= rng2_io_rand_bits[31]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sqrt_log_io_uniform_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sqrt_log_io_uniform_v <= rng2_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      sqrt_log_io_uniform_b <= _sqrt_log_io_uniform_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sign_adjustedPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sign_adjustedPipe_valid <= sqrt_log_io_result_valid; // @[Valid.scala 127:22]
    end
    if (sqrt_log_io_result_valid) begin // @[Reg.scala 17:18]
      if (signPipe_bits) begin // @[BoxMuller.scala 91:8]
        sign_adjustedPipe_bits <= _sign_adjusted_T_3;
      end else begin
        sign_adjustedPipe_bits <= sqrt_log_io_result_bits;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g1_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g1_v <= _io_g1_T; // @[Valid.scala 127:22]
    end
    if (_io_g1_T) begin // @[Reg.scala 17:18]
      io_g1_b <= _io_g1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g2_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g2_v <= _io_g2_T; // @[Valid.scala 127:22]
    end
    if (_io_g2_T) begin // @[Reg.scala 17:18]
      io_g2_b <= _io_g2_T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quadrantPipe_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  quadrantPipe_bits = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  quadrantPipe_valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  quadrantPipe_bits_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  quadrantPipe_valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  quadrantPipe_bits_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  quadrantPipe_valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quadrantPipe_bits_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  quadrantPipe_valid_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  quadrantPipe_bits_4 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  quadrantPipe_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  quadrantPipe_bits_5 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  quadrantPipe_valid_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  quadrantPipe_bits_6 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  quadrantPipe_valid_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  quadrantPipe_bits_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  quadrantPipe_valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  quadrantPipe_bits_8 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  quadrantPipe_valid_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  quadrantPipe_bits_9 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  quadrantPipe_valid_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  quadrantPipe_bits_10 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  quadrantPipe_valid_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  quadrantPipe_bits_11 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  quadrantPipe_valid_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  quadrantPipe_bits_12 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  quadrantPipe_valid_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  quadrantPipe_bits_13 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  quadrantPipe_valid_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  quadrantPipe_bits_14 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  quadrantPipe_valid_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  quadrantPipe_bits_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  quadrantPipe_valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  quadrantPipe_bits_16 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  quadrantPipe_valid_17 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  quadrantPipe_bits_17 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  quadrantPipe_valid_18 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  quadrantPipe_bits_18 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  quadrantPipe_valid_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  quadrantPipe_bits_19 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  quadrantPipe_valid_20 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  quadrantPipe_bits_20 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  quadrantPipe_valid_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  quadrantPipe_bits_21 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  quadrantPipe_valid_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  quadrantPipe_bits_22 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  quadrantPipe_valid_23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  quadrantPipe_bits_23 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  quadrantPipe_valid_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  quadrantPipe_bits_24 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  quadrantPipe_valid_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  quadrantPipe_bits_25 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  quadrantPipe_valid_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  quadrantPipe_bits_26 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  quadrantPipe_valid_27 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  quadrantPipe_bits_27 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  quadrantPipe_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  quadrantPipe_bits_28 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  quadrantPipe_valid_29 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  quadrantPipe_bits_29 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  quadrantPipe_valid_30 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  quadrantPipe_bits_30 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  quadrantPipe_bits_31 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  trigonometric_io_theta_v = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  trigonometric_io_theta_b = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cosinePipe_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cosinePipe_bits = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sinePipe_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sinePipe_bits = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  signPipe_bits = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sqrt_log_io_uniform_v = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sqrt_log_io_uniform_b = _RAND_71[28:0];
  _RAND_72 = {1{`RANDOM}};
  sign_adjustedPipe_valid = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  sign_adjustedPipe_bits = _RAND_73[51:0];
  _RAND_74 = {1{`RANDOM}};
  io_g1_v = _RAND_74[0:0];
  _RAND_75 = {3{`RANDOM}};
  io_g1_b = _RAND_75[83:0];
  _RAND_76 = {1{`RANDOM}};
  io_g2_v = _RAND_76[0:0];
  _RAND_77 = {3{`RANDOM}};
  io_g2_b = _RAND_77[83:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MonteCarlo_14(
  input         clock,
  input         reset,
  output        io_request_0_ready,
  input         io_request_0_valid,
  input  [31:0] io_request_0_bits_time_steps,
  input  [31:0] io_request_0_bits_start_value,
  input  [31:0] io_request_0_bits_coefficient1,
  input  [31:0] io_request_0_bits_coefficient2,
  output        io_request_1_ready,
  input         io_request_1_valid,
  input  [31:0] io_request_1_bits_time_steps,
  input  [31:0] io_request_1_bits_start_value,
  input  [31:0] io_request_1_bits_coefficient1,
  input  [31:0] io_request_1_bits_coefficient2,
  input         io_response_0_ready,
  output        io_response_0_valid,
  output [31:0] io_response_0_bits,
  input         io_response_1_ready,
  output        io_response_1_valid,
  output [31:0] io_response_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rng_clock; // @[MonteCarlo.scala 42:19]
  wire  rng_reset; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g1_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g1_bits; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g2_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g2_bits; // @[MonteCarlo.scala 42:19]
  wire  initialized = rng_io_g1_valid & rng_io_g2_valid; // @[MonteCarlo.scala 47:37]
  reg [2:0] state; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_2 = $signed(io_request_0_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_3 = io_request_0_ready & io_request_0_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1; // @[Reg.scala 16:16]
  reg [31:0] c2; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_1 = io_request_0_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step; // @[Reg.scala 16:16]
  reg [31:0] price; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T = $signed(price) * $signed(c1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T = $signed(rng_io_g1_bits) * $signed(c2); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T = $signed(price) * $signed(partial_res2); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_2 = $signed(partial_res3) + $signed(partial_res1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_3 = counter == last_step ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_4 = counter == last_step ? counter : _counter_T_1; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_7 = io_response_0_ready & io_response_0_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_5 = _T_7 ? 3'h1 : state; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_6 = 3'h5 == state ? _GEN_5 : state; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_7 = 3'h4 == state ? $signed(_price_T_2) : $signed(price); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_3 : _GEN_6; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_9 = 3'h4 == state ? _GEN_4 : counter; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_64 = {$signed(partial_res3), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_10 = 3'h3 == state ? $signed(_partial_res3_T) : $signed({{12{_GEN_64[51]}},_GEN_64}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_11 = 3'h3 == state ? 3'h4 : _GEN_8; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_65 = {$signed(partial_res1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_14 = 3'h2 == state ? $signed(_partial_res1_T) : $signed({{12{_GEN_65[51]}},_GEN_65}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_66 = {$signed(partial_res2), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_15 = 3'h2 == state ? $signed(_partial_res2_T) : $signed({{20{_GEN_66[63]}},_GEN_66}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_17 = 3'h2 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_10); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_23 = 3'h1 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_14); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_24 = 3'h1 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_15); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_25 = 3'h1 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_17); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_29 = 3'h0 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_23); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_30 = 3'h0 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_24); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_31 = 3'h0 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_25); // @[MonteCarlo.scala 66:19 60:27]
  reg [2:0] state_1; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_6 = $signed(io_request_1_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_7 = io_request_1_ready & io_request_1_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1_1; // @[Reg.scala 16:16]
  reg [31:0] c2_1; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_4 = io_request_1_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step_1; // @[Reg.scala 16:16]
  reg [31:0] price_1; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1_1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2_1; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3_1; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter_1; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T_1 = $signed(price_1) * $signed(c1_1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T_1 = $signed(rng_io_g2_bits) * $signed(c2_1); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T_1 = $signed(price_1) * $signed(partial_res2_1); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_5 = $signed(partial_res3_1) + $signed(partial_res1_1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_35 = counter_1 == last_step_1 ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_36 = counter_1 == last_step_1 ? counter_1 : _counter_T_3; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_15 = io_response_1_ready & io_response_1_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_37 = _T_15 ? 3'h1 : state_1; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_38 = 3'h5 == state_1 ? _GEN_37 : state_1; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_39 = 3'h4 == state_1 ? $signed(_price_T_5) : $signed(price_1); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_40 = 3'h4 == state_1 ? _GEN_35 : _GEN_38; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_41 = 3'h4 == state_1 ? _GEN_36 : counter_1; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_74 = {$signed(partial_res3_1), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_42 = 3'h3 == state_1 ? $signed(_partial_res3_T_1) : $signed({{12{_GEN_74[51]}},_GEN_74}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_43 = 3'h3 == state_1 ? 3'h4 : _GEN_40; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_75 = {$signed(partial_res1_1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_46 = 3'h2 == state_1 ? $signed(_partial_res1_T_1) : $signed({{12{_GEN_75[51]}},_GEN_75}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_76 = {$signed(partial_res2_1), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_47 = 3'h2 == state_1 ? $signed(_partial_res2_T_1) : $signed({{20{_GEN_76[63]}},_GEN_76}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_49 = 3'h2 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_42); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_55 = 3'h1 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_46); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_56 = 3'h1 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_47); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_57 = 3'h1 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_49); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_61 = 3'h0 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_55); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_62 = 3'h0 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_56); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_63 = 3'h0 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_57); // @[MonteCarlo.scala 66:19 60:27]
  wire [43:0] _GEN_84 = _GEN_29[63:20];
  wire [51:0] _GEN_86 = _GEN_30[83:32];
  wire [43:0] _GEN_88 = _GEN_31[63:20];
  wire [43:0] _GEN_90 = _GEN_61[63:20];
  wire [51:0] _GEN_92 = _GEN_62[83:32];
  wire [43:0] _GEN_94 = _GEN_63[63:20];
  BoxMuller_14 rng ( // @[MonteCarlo.scala 42:19]
    .clock(rng_clock),
    .reset(rng_reset),
    .io_g1_valid(rng_io_g1_valid),
    .io_g1_bits(rng_io_g1_bits),
    .io_g2_valid(rng_io_g2_valid),
    .io_g2_bits(rng_io_g2_bits)
  );
  assign io_request_0_ready = state == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_request_1_ready = state_1 == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_response_0_valid = state == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_0_bits = price; // @[MonteCarlo.scala 65:16]
  assign io_response_1_valid = state_1 == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_1_bits = price_1; // @[MonteCarlo.scala 65:16]
  assign rng_clock = clock;
  assign rng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state <= 3'h1;
      end else begin
        state <= 3'h0;
      end
    end else if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_3) begin // @[MonteCarlo.scala 71:23]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[MonteCarlo.scala 66:19]
      state <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state <= _GEN_11;
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c1 <= _c1_T_2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c2 <= io_request_0_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      last_step <= _last_step_T_1; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        price <= io_request_0_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          price <= _GEN_7;
        end
      end
    end
    partial_res1 <= _GEN_84[31:0];
    partial_res2 <= _GEN_86[31:0];
    partial_res3 <= _GEN_88[31:0];
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        counter <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          counter <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state_1 <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state_1 <= 3'h1;
      end else begin
        state_1 <= 3'h0;
      end
    end else if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_7) begin // @[MonteCarlo.scala 71:23]
        state_1 <= 3'h2;
      end else begin
        state_1 <= 3'h1;
      end
    end else if (3'h2 == state_1) begin // @[MonteCarlo.scala 66:19]
      state_1 <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state_1 <= _GEN_43;
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c1_1 <= _c1_T_6; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c2_1 <= io_request_1_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      last_step_1 <= _last_step_T_4; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        price_1 <= io_request_1_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          price_1 <= _GEN_39;
        end
      end
    end
    partial_res1_1 <= _GEN_90[31:0];
    partial_res2_1 <= _GEN_92[31:0];
    partial_res3_1 <= _GEN_94[31:0];
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        counter_1 <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          counter_1 <= _GEN_41;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  c1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_step = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  price = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  partial_res1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  partial_res2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  partial_res3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  c1_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_step_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  price_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  partial_res1_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  partial_res2_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  partial_res3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  counter_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_30(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h36afeaf3 : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h54c5f36 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h9e7d92 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TauswortheUniform_31(
  input         clock,
  input         reset,
  output        io_rand_valid,
  output [31:0] io_rand_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] s0_reg; // @[BoxMuller.scala 20:23]
  reg [31:0] s1_reg; // @[BoxMuller.scala 21:23]
  reg [31:0] s2_reg; // @[BoxMuller.scala 22:23]
  wire [44:0] _GEN_4 = {s0_reg, 13'h0}; // @[BoxMuller.scala 27:23]
  wire [46:0] _b_T = {{2'd0}, _GEN_4}; // @[BoxMuller.scala 27:23]
  wire [46:0] _GEN_5 = {{15'd0}, s0_reg}; // @[BoxMuller.scala 27:32]
  wire [46:0] _b_T_1 = _b_T ^ _GEN_5; // @[BoxMuller.scala 27:32]
  wire [46:0] b = {{19'd0}, _b_T_1[46:19]}; // @[BoxMuller.scala 27:42]
  wire [31:0] _s0_reg_T = s0_reg & 32'hfffffffe; // @[BoxMuller.scala 28:25]
  wire [43:0] _GEN_7 = {_s0_reg_T, 12'h0}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_1 = {{3'd0}, _GEN_7}; // @[BoxMuller.scala 28:48]
  wire [46:0] _s0_reg_T_2 = _s0_reg_T_1 ^ b; // @[BoxMuller.scala 28:57]
  wire [33:0] _GEN_8 = {s1_reg, 2'h0}; // @[BoxMuller.scala 31:23]
  wire [34:0] _b_T_2 = {{1'd0}, _GEN_8}; // @[BoxMuller.scala 31:23]
  wire [34:0] _GEN_9 = {{3'd0}, s1_reg}; // @[BoxMuller.scala 31:31]
  wire [34:0] _b_T_3 = _b_T_2 ^ _GEN_9; // @[BoxMuller.scala 31:31]
  wire [34:0] b_1 = {{25'd0}, _b_T_3[34:25]}; // @[BoxMuller.scala 31:41]
  wire [31:0] _s1_reg_T = s1_reg & 32'hfffffff8; // @[BoxMuller.scala 32:25]
  wire [35:0] _GEN_11 = {_s1_reg_T, 4'h0}; // @[BoxMuller.scala 32:48]
  wire [38:0] _s1_reg_T_1 = {{3'd0}, _GEN_11}; // @[BoxMuller.scala 32:48]
  wire [38:0] _GEN_12 = {{4'd0}, b_1}; // @[BoxMuller.scala 32:56]
  wire [38:0] _s1_reg_T_2 = _s1_reg_T_1 ^ _GEN_12; // @[BoxMuller.scala 32:56]
  wire [34:0] _b_T_4 = {s2_reg, 3'h0}; // @[BoxMuller.scala 35:23]
  wire [34:0] _GEN_13 = {{3'd0}, s2_reg}; // @[BoxMuller.scala 35:31]
  wire [34:0] _b_T_5 = _b_T_4 ^ _GEN_13; // @[BoxMuller.scala 35:31]
  wire [34:0] b_2 = {{11'd0}, _b_T_5[34:11]}; // @[BoxMuller.scala 35:41]
  wire [31:0] _s2_reg_T = s2_reg & 32'hfffffff0; // @[BoxMuller.scala 36:25]
  wire [48:0] _GEN_15 = {_s2_reg_T, 17'h0}; // @[BoxMuller.scala 36:48]
  wire [62:0] _s2_reg_T_1 = {{14'd0}, _GEN_15}; // @[BoxMuller.scala 36:48]
  wire [62:0] _GEN_16 = {{28'd0}, b_2}; // @[BoxMuller.scala 36:57]
  wire [62:0] _s2_reg_T_2 = _s2_reg_T_1 ^ _GEN_16; // @[BoxMuller.scala 36:57]
  wire [31:0] _io_rand_T = s0_reg ^ s1_reg; // @[BoxMuller.scala 39:35]
  reg  io_rand_v; // @[Valid.scala 127:22]
  reg [31:0] io_rand_b; // @[Reg.scala 16:16]
  wire [46:0] _GEN_17 = reset ? 47'h1a8bae5d : _s0_reg_T_2; // @[BoxMuller.scala 20:{23,23}]
  wire [38:0] _GEN_18 = reset ? 39'h2c4e8756 : _s1_reg_T_2; // @[BoxMuller.scala 21:{23,23}]
  wire [62:0] _GEN_19 = reset ? 63'h101cc2e9 : _s2_reg_T_2; // @[BoxMuller.scala 22:{23,23}]
  assign io_rand_valid = io_rand_v; // @[Valid.scala 122:21 123:17]
  assign io_rand_bits = io_rand_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    s0_reg <= _GEN_17[31:0]; // @[BoxMuller.scala 20:{23,23}]
    s1_reg <= _GEN_18[31:0]; // @[BoxMuller.scala 21:{23,23}]
    s2_reg <= _GEN_19[31:0]; // @[BoxMuller.scala 22:{23,23}]
    if (reset) begin // @[Valid.scala 127:22]
      io_rand_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_rand_v <= 1'h1; // @[Valid.scala 127:22]
    end
    io_rand_b <= _io_rand_T ^ s2_reg; // @[BoxMuller.scala 39:44]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s0_reg = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  s1_reg = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  s2_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  io_rand_v = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_rand_b = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BoxMuller_15(
  input         clock,
  input         reset,
  output        io_g1_valid,
  output [51:0] io_g1_bits,
  output        io_g2_valid,
  output [51:0] io_g2_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [63:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [95:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [95:0] _RAND_77;
`endif // RANDOMIZE_REG_INIT
  wire  rng1_clock; // @[BoxMuller.scala 51:20]
  wire  rng1_reset; // @[BoxMuller.scala 51:20]
  wire  rng1_io_rand_valid; // @[BoxMuller.scala 51:20]
  wire [31:0] rng1_io_rand_bits; // @[BoxMuller.scala 51:20]
  wire  rng2_clock; // @[BoxMuller.scala 52:20]
  wire  rng2_reset; // @[BoxMuller.scala 52:20]
  wire  rng2_io_rand_valid; // @[BoxMuller.scala 52:20]
  wire [31:0] rng2_io_rand_bits; // @[BoxMuller.scala 52:20]
  wire  trigonometric_clock; // @[BoxMuller.scala 55:29]
  wire  trigonometric_reset; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_theta_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_theta_bits; // @[BoxMuller.scala 55:29]
  wire  trigonometric_io_result_valid; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_sine; // @[BoxMuller.scala 55:29]
  wire [31:0] trigonometric_io_result_bits_cosine; // @[BoxMuller.scala 55:29]
  wire  sqrt_log_clock; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_reset; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_uniform_valid; // @[BoxMuller.scala 84:24]
  wire [31:0] sqrt_log_io_uniform_bits; // @[BoxMuller.scala 84:24]
  wire  sqrt_log_io_result_valid; // @[BoxMuller.scala 84:24]
  wire [51:0] sqrt_log_io_result_bits; // @[BoxMuller.scala 84:24]
  wire [30:0] _theta_T_3 = {2'h0,rng1_io_rand_bits[28:0]}; // @[BoxMuller.scala 62:18]
  wire [62:0] _theta_T_4 = $signed(_theta_T_3) * 32'sh6487ed51; // @[BoxMuller.scala 62:26]
  reg  quadrantPipe_valid; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_1; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_1; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_2; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_2; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_3; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_3; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_4; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_4; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_5; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_5; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_6; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_6; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_7; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_7; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_8; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_8; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_9; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_9; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_10; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_10; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_11; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_11; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_12; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_12; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_13; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_13; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_14; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_14; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_15; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_15; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_16; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_16; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_17; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_17; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_18; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_18; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_19; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_19; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_20; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_20; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_21; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_21; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_22; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_22; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_23; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_23; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_24; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_24; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_25; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_25; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_26; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_26; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_27; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_27; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_28; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_28; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_29; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_29; // @[Reg.scala 16:16]
  reg  quadrantPipe_valid_30; // @[Valid.scala 127:22]
  reg [1:0] quadrantPipe_bits_30; // @[Reg.scala 16:16]
  reg [1:0] quadrantPipe_bits_31; // @[Reg.scala 16:16]
  reg  trigonometric_io_theta_v; // @[Valid.scala 127:22]
  reg [31:0] trigonometric_io_theta_b; // @[Reg.scala 16:16]
  wire [33:0] _GEN_40 = _theta_T_4[62:29]; // @[BoxMuller.scala 59:19 61:9]
  wire [31:0] theta = _GEN_40[31:0]; // @[BoxMuller.scala 59:19 61:9]
  wire  _cosine_T = quadrantPipe_bits_31 == 2'h0; // @[BoxMuller.scala 70:21]
  wire  _cosine_T_2 = quadrantPipe_bits_31 == 2'h0 | quadrantPipe_bits_31 == 2'h3; // @[BoxMuller.scala 70:29]
  wire [31:0] _cosine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_cosine); // @[BoxMuller.scala 72:7]
  reg  cosinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] cosinePipe_bits; // @[Reg.scala 16:16]
  wire  _sine_T_2 = _cosine_T | quadrantPipe_bits_31 == 2'h2; // @[BoxMuller.scala 78:29]
  wire [31:0] _sine_T_5 = 32'sh0 - $signed(trigonometric_io_result_bits_sine); // @[BoxMuller.scala 80:7]
  reg  sinePipe_valid; // @[Valid.scala 127:22]
  reg [31:0] sinePipe_bits; // @[Reg.scala 16:16]
  reg  signPipe_bits; // @[Reg.scala 16:16]
  wire [28:0] _sqrt_log_io_uniform_T_1 = rng2_io_rand_bits[28:0]; // @[BoxMuller.scala 87:89]
  reg  sqrt_log_io_uniform_v; // @[Valid.scala 127:22]
  reg [28:0] sqrt_log_io_uniform_b; // @[Reg.scala 16:16]
  wire [51:0] _sign_adjusted_T_3 = 52'sh0 - $signed(sqrt_log_io_result_bits); // @[BoxMuller.scala 93:7]
  reg  sign_adjustedPipe_valid; // @[Valid.scala 127:22]
  reg [51:0] sign_adjustedPipe_bits; // @[Reg.scala 16:16]
  wire  _io_g1_T = sign_adjustedPipe_valid & cosinePipe_valid; // @[BoxMuller.scala 99:25]
  wire [83:0] _io_g1_T_1 = $signed(cosinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 100:17]
  reg  io_g1_v; // @[Valid.scala 127:22]
  reg [83:0] io_g1_b; // @[Reg.scala 16:16]
  wire  _io_g2_T = sign_adjustedPipe_valid & sinePipe_valid; // @[BoxMuller.scala 103:25]
  wire [83:0] _io_g2_T_1 = $signed(sinePipe_bits) * $signed(sign_adjustedPipe_bits); // @[BoxMuller.scala 104:15]
  reg  io_g2_v; // @[Valid.scala 127:22]
  reg [83:0] io_g2_b; // @[Reg.scala 16:16]
  wire [53:0] _GEN_42 = io_g1_b[83:30]; // @[BoxMuller.scala 98:9]
  wire [53:0] _GEN_44 = io_g2_b[83:30]; // @[BoxMuller.scala 102:9]
  wire [32:0] _GEN_46 = {$signed(trigonometric_io_theta_b), 1'h0}; // @[BoxMuller.scala 65:26]
  TauswortheUniform_30 rng1 ( // @[BoxMuller.scala 51:20]
    .clock(rng1_clock),
    .reset(rng1_reset),
    .io_rand_valid(rng1_io_rand_valid),
    .io_rand_bits(rng1_io_rand_bits)
  );
  TauswortheUniform_31 rng2 ( // @[BoxMuller.scala 52:20]
    .clock(rng2_clock),
    .reset(rng2_reset),
    .io_rand_valid(rng2_io_rand_valid),
    .io_rand_bits(rng2_io_rand_bits)
  );
  Trigonometric trigonometric ( // @[BoxMuller.scala 55:29]
    .clock(trigonometric_clock),
    .reset(trigonometric_reset),
    .io_theta_valid(trigonometric_io_theta_valid),
    .io_theta_bits(trigonometric_io_theta_bits),
    .io_result_valid(trigonometric_io_result_valid),
    .io_result_bits_sine(trigonometric_io_result_bits_sine),
    .io_result_bits_cosine(trigonometric_io_result_bits_cosine)
  );
  SquareRootLog sqrt_log ( // @[BoxMuller.scala 84:24]
    .clock(sqrt_log_clock),
    .reset(sqrt_log_reset),
    .io_uniform_valid(sqrt_log_io_uniform_valid),
    .io_uniform_bits(sqrt_log_io_uniform_bits),
    .io_result_valid(sqrt_log_io_result_valid),
    .io_result_bits(sqrt_log_io_result_bits)
  );
  assign io_g1_valid = io_g1_v; // @[Valid.scala 122:21 123:17]
  assign io_g1_bits = _GEN_42[51:0]; // @[BoxMuller.scala 98:9]
  assign io_g2_valid = io_g2_v; // @[Valid.scala 122:21 123:17]
  assign io_g2_bits = _GEN_44[51:0]; // @[BoxMuller.scala 102:9]
  assign rng1_clock = clock;
  assign rng1_reset = reset;
  assign rng2_clock = clock;
  assign rng2_reset = reset;
  assign trigonometric_clock = clock;
  assign trigonometric_reset = reset;
  assign trigonometric_io_theta_valid = trigonometric_io_theta_v; // @[Valid.scala 122:21 123:17]
  assign trigonometric_io_theta_bits = _GEN_46[31:0]; // @[BoxMuller.scala 65:26]
  assign sqrt_log_clock = clock;
  assign sqrt_log_reset = reset;
  assign sqrt_log_io_uniform_valid = sqrt_log_io_uniform_v; // @[Valid.scala 122:21 123:17]
  assign sqrt_log_io_uniform_bits = {{3{sqrt_log_io_uniform_b[28]}},sqrt_log_io_uniform_b}; // @[BoxMuller.scala 87:23]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits <= rng1_io_rand_bits[31:30]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_1 <= quadrantPipe_valid; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_1 <= quadrantPipe_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_2 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_2 <= quadrantPipe_valid_1; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_1) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_2 <= quadrantPipe_bits_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_3 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_3 <= quadrantPipe_valid_2; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_2) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_3 <= quadrantPipe_bits_2; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_4 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_4 <= quadrantPipe_valid_3; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_3) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_4 <= quadrantPipe_bits_3; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_5 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_5 <= quadrantPipe_valid_4; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_4) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_5 <= quadrantPipe_bits_4; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_6 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_6 <= quadrantPipe_valid_5; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_5) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_6 <= quadrantPipe_bits_5; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_7 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_7 <= quadrantPipe_valid_6; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_6) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_7 <= quadrantPipe_bits_6; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_8 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_8 <= quadrantPipe_valid_7; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_7) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_8 <= quadrantPipe_bits_7; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_9 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_9 <= quadrantPipe_valid_8; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_8) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_9 <= quadrantPipe_bits_8; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_10 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_10 <= quadrantPipe_valid_9; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_9) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_10 <= quadrantPipe_bits_9; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_11 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_11 <= quadrantPipe_valid_10; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_10) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_11 <= quadrantPipe_bits_10; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_12 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_12 <= quadrantPipe_valid_11; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_11) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_12 <= quadrantPipe_bits_11; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_13 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_13 <= quadrantPipe_valid_12; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_12) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_13 <= quadrantPipe_bits_12; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_14 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_14 <= quadrantPipe_valid_13; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_13) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_14 <= quadrantPipe_bits_13; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_15 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_15 <= quadrantPipe_valid_14; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_14) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_15 <= quadrantPipe_bits_14; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_16 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_16 <= quadrantPipe_valid_15; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_15) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_16 <= quadrantPipe_bits_15; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_17 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_17 <= quadrantPipe_valid_16; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_16) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_17 <= quadrantPipe_bits_16; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_18 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_18 <= quadrantPipe_valid_17; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_17) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_18 <= quadrantPipe_bits_17; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_19 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_19 <= quadrantPipe_valid_18; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_18) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_19 <= quadrantPipe_bits_18; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_20 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_20 <= quadrantPipe_valid_19; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_19) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_20 <= quadrantPipe_bits_19; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_21 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_21 <= quadrantPipe_valid_20; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_20) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_21 <= quadrantPipe_bits_20; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_22 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_22 <= quadrantPipe_valid_21; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_21) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_22 <= quadrantPipe_bits_21; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_23 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_23 <= quadrantPipe_valid_22; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_22) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_23 <= quadrantPipe_bits_22; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_24 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_24 <= quadrantPipe_valid_23; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_23) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_24 <= quadrantPipe_bits_23; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_25 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_25 <= quadrantPipe_valid_24; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_24) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_25 <= quadrantPipe_bits_24; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_26 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_26 <= quadrantPipe_valid_25; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_25) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_26 <= quadrantPipe_bits_25; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_27 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_27 <= quadrantPipe_valid_26; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_26) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_27 <= quadrantPipe_bits_26; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_28 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_28 <= quadrantPipe_valid_27; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_27) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_28 <= quadrantPipe_bits_27; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_29 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_29 <= quadrantPipe_valid_28; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_28) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_29 <= quadrantPipe_bits_28; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      quadrantPipe_valid_30 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      quadrantPipe_valid_30 <= quadrantPipe_valid_29; // @[Valid.scala 127:22]
    end
    if (quadrantPipe_valid_29) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_30 <= quadrantPipe_bits_29; // @[Reg.scala 17:22]
    end
    if (quadrantPipe_valid_30) begin // @[Reg.scala 17:18]
      quadrantPipe_bits_31 <= quadrantPipe_bits_30; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      trigonometric_io_theta_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      trigonometric_io_theta_v <= rng1_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng1_io_rand_valid) begin // @[Reg.scala 17:18]
      trigonometric_io_theta_b <= theta; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      cosinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      cosinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_cosine_T_2) begin // @[BoxMuller.scala 69:8]
        cosinePipe_bits <= trigonometric_io_result_bits_cosine;
      end else begin
        cosinePipe_bits <= _cosine_T_5;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      sinePipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sinePipe_valid <= trigonometric_io_result_valid; // @[Valid.scala 127:22]
    end
    if (trigonometric_io_result_valid) begin // @[Reg.scala 17:18]
      if (_sine_T_2) begin // @[BoxMuller.scala 77:8]
        sinePipe_bits <= trigonometric_io_result_bits_sine;
      end else begin
        sinePipe_bits <= _sine_T_5;
      end
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      signPipe_bits <= rng2_io_rand_bits[31]; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sqrt_log_io_uniform_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sqrt_log_io_uniform_v <= rng2_io_rand_valid; // @[Valid.scala 127:22]
    end
    if (rng2_io_rand_valid) begin // @[Reg.scala 17:18]
      sqrt_log_io_uniform_b <= _sqrt_log_io_uniform_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      sign_adjustedPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      sign_adjustedPipe_valid <= sqrt_log_io_result_valid; // @[Valid.scala 127:22]
    end
    if (sqrt_log_io_result_valid) begin // @[Reg.scala 17:18]
      if (signPipe_bits) begin // @[BoxMuller.scala 91:8]
        sign_adjustedPipe_bits <= _sign_adjusted_T_3;
      end else begin
        sign_adjustedPipe_bits <= sqrt_log_io_result_bits;
      end
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g1_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g1_v <= _io_g1_T; // @[Valid.scala 127:22]
    end
    if (_io_g1_T) begin // @[Reg.scala 17:18]
      io_g1_b <= _io_g1_T_1; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_g2_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_g2_v <= _io_g2_T; // @[Valid.scala 127:22]
    end
    if (_io_g2_T) begin // @[Reg.scala 17:18]
      io_g2_b <= _io_g2_T_1; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  quadrantPipe_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  quadrantPipe_bits = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  quadrantPipe_valid_1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  quadrantPipe_bits_1 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  quadrantPipe_valid_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  quadrantPipe_bits_2 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  quadrantPipe_valid_3 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  quadrantPipe_bits_3 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  quadrantPipe_valid_4 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  quadrantPipe_bits_4 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  quadrantPipe_valid_5 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  quadrantPipe_bits_5 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  quadrantPipe_valid_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  quadrantPipe_bits_6 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  quadrantPipe_valid_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  quadrantPipe_bits_7 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  quadrantPipe_valid_8 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  quadrantPipe_bits_8 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  quadrantPipe_valid_9 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  quadrantPipe_bits_9 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  quadrantPipe_valid_10 = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  quadrantPipe_bits_10 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  quadrantPipe_valid_11 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  quadrantPipe_bits_11 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  quadrantPipe_valid_12 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  quadrantPipe_bits_12 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  quadrantPipe_valid_13 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  quadrantPipe_bits_13 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  quadrantPipe_valid_14 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  quadrantPipe_bits_14 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  quadrantPipe_valid_15 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  quadrantPipe_bits_15 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  quadrantPipe_valid_16 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  quadrantPipe_bits_16 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  quadrantPipe_valid_17 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  quadrantPipe_bits_17 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  quadrantPipe_valid_18 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  quadrantPipe_bits_18 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  quadrantPipe_valid_19 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  quadrantPipe_bits_19 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  quadrantPipe_valid_20 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  quadrantPipe_bits_20 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  quadrantPipe_valid_21 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  quadrantPipe_bits_21 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  quadrantPipe_valid_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  quadrantPipe_bits_22 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  quadrantPipe_valid_23 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  quadrantPipe_bits_23 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  quadrantPipe_valid_24 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  quadrantPipe_bits_24 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  quadrantPipe_valid_25 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  quadrantPipe_bits_25 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  quadrantPipe_valid_26 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  quadrantPipe_bits_26 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  quadrantPipe_valid_27 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  quadrantPipe_bits_27 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  quadrantPipe_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  quadrantPipe_bits_28 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  quadrantPipe_valid_29 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  quadrantPipe_bits_29 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  quadrantPipe_valid_30 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  quadrantPipe_bits_30 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  quadrantPipe_bits_31 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  trigonometric_io_theta_v = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  trigonometric_io_theta_b = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  cosinePipe_valid = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cosinePipe_bits = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  sinePipe_valid = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  sinePipe_bits = _RAND_68[31:0];
  _RAND_69 = {1{`RANDOM}};
  signPipe_bits = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  sqrt_log_io_uniform_v = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  sqrt_log_io_uniform_b = _RAND_71[28:0];
  _RAND_72 = {1{`RANDOM}};
  sign_adjustedPipe_valid = _RAND_72[0:0];
  _RAND_73 = {2{`RANDOM}};
  sign_adjustedPipe_bits = _RAND_73[51:0];
  _RAND_74 = {1{`RANDOM}};
  io_g1_v = _RAND_74[0:0];
  _RAND_75 = {3{`RANDOM}};
  io_g1_b = _RAND_75[83:0];
  _RAND_76 = {1{`RANDOM}};
  io_g2_v = _RAND_76[0:0];
  _RAND_77 = {3{`RANDOM}};
  io_g2_b = _RAND_77[83:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MonteCarlo_15(
  input         clock,
  input         reset,
  output        io_request_0_ready,
  input         io_request_0_valid,
  input  [31:0] io_request_0_bits_time_steps,
  input  [31:0] io_request_0_bits_start_value,
  input  [31:0] io_request_0_bits_coefficient1,
  input  [31:0] io_request_0_bits_coefficient2,
  output        io_request_1_ready,
  input         io_request_1_valid,
  input  [31:0] io_request_1_bits_time_steps,
  input  [31:0] io_request_1_bits_start_value,
  input  [31:0] io_request_1_bits_coefficient1,
  input  [31:0] io_request_1_bits_coefficient2,
  input         io_response_0_ready,
  output        io_response_0_valid,
  output [31:0] io_response_0_bits,
  input         io_response_1_ready,
  output        io_response_1_valid,
  output [31:0] io_response_1_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire  rng_clock; // @[MonteCarlo.scala 42:19]
  wire  rng_reset; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g1_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g1_bits; // @[MonteCarlo.scala 42:19]
  wire  rng_io_g2_valid; // @[MonteCarlo.scala 42:19]
  wire [51:0] rng_io_g2_bits; // @[MonteCarlo.scala 42:19]
  wire  initialized = rng_io_g1_valid & rng_io_g2_valid; // @[MonteCarlo.scala 47:37]
  reg [2:0] state; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_2 = $signed(io_request_0_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_3 = io_request_0_ready & io_request_0_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1; // @[Reg.scala 16:16]
  reg [31:0] c2; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_1 = io_request_0_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step; // @[Reg.scala 16:16]
  reg [31:0] price; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T = $signed(price) * $signed(c1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T = $signed(rng_io_g1_bits) * $signed(c2); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T = $signed(price) * $signed(partial_res2); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_2 = $signed(partial_res3) + $signed(partial_res1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_1 = counter + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_3 = counter == last_step ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_4 = counter == last_step ? counter : _counter_T_1; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_7 = io_response_0_ready & io_response_0_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_5 = _T_7 ? 3'h1 : state; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_6 = 3'h5 == state ? _GEN_5 : state; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_7 = 3'h4 == state ? $signed(_price_T_2) : $signed(price); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_8 = 3'h4 == state ? _GEN_3 : _GEN_6; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_9 = 3'h4 == state ? _GEN_4 : counter; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_64 = {$signed(partial_res3), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_10 = 3'h3 == state ? $signed(_partial_res3_T) : $signed({{12{_GEN_64[51]}},_GEN_64}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_11 = 3'h3 == state ? 3'h4 : _GEN_8; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_65 = {$signed(partial_res1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_14 = 3'h2 == state ? $signed(_partial_res1_T) : $signed({{12{_GEN_65[51]}},_GEN_65}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_66 = {$signed(partial_res2), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_15 = 3'h2 == state ? $signed(_partial_res2_T) : $signed({{20{_GEN_66[63]}},_GEN_66}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_17 = 3'h2 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_10); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_23 = 3'h1 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_14); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_24 = 3'h1 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_15); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_25 = 3'h1 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_17); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_29 = 3'h0 == state ? $signed({{12{_GEN_65[51]}},_GEN_65}) : $signed(_GEN_23); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_30 = 3'h0 == state ? $signed({{20{_GEN_66[63]}},_GEN_66}) : $signed(_GEN_24); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_31 = 3'h0 == state ? $signed({{12{_GEN_64[51]}},_GEN_64}) : $signed(_GEN_25); // @[MonteCarlo.scala 66:19 60:27]
  reg [2:0] state_1; // @[MonteCarlo.scala 52:24]
  wire [31:0] _c1_T_6 = $signed(io_request_1_bits_coefficient1) + 32'sh100000; // @[MonteCarlo.scala 54:56]
  wire  _c1_T_7 = io_request_1_ready & io_request_1_valid; // @[Decoupled.scala 50:35]
  reg [31:0] c1_1; // @[Reg.scala 16:16]
  reg [31:0] c2_1; // @[Reg.scala 16:16]
  wire [31:0] _last_step_T_4 = io_request_1_bits_time_steps - 32'h1; // @[MonteCarlo.scala 56:54]
  reg [31:0] last_step_1; // @[Reg.scala 16:16]
  reg [31:0] price_1; // @[MonteCarlo.scala 57:27]
  reg [31:0] partial_res1_1; // @[MonteCarlo.scala 58:27]
  reg [31:0] partial_res2_1; // @[MonteCarlo.scala 59:27]
  reg [31:0] partial_res3_1; // @[MonteCarlo.scala 60:27]
  reg [31:0] counter_1; // @[MonteCarlo.scala 62:22]
  wire [63:0] _partial_res1_T_1 = $signed(price_1) * $signed(c1_1); // @[MonteCarlo.scala 77:31]
  wire [83:0] _partial_res2_T_1 = $signed(rng_io_g2_bits) * $signed(c2_1); // @[MonteCarlo.scala 78:32]
  wire [63:0] _partial_res3_T_1 = $signed(price_1) * $signed(partial_res2_1); // @[MonteCarlo.scala 82:31]
  wire [31:0] _price_T_5 = $signed(partial_res3_1) + $signed(partial_res1_1); // @[MonteCarlo.scala 86:31]
  wire [31:0] _counter_T_3 = counter_1 + 32'h1; // @[MonteCarlo.scala 91:30]
  wire [2:0] _GEN_35 = counter_1 == last_step_1 ? 3'h5 : 3'h2; // @[MonteCarlo.scala 87:37 88:17 90:19]
  wire [31:0] _GEN_36 = counter_1 == last_step_1 ? counter_1 : _counter_T_3; // @[MonteCarlo.scala 62:22 87:37 91:19]
  wire  _T_15 = io_response_1_ready & io_response_1_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_37 = _T_15 ? 3'h1 : state_1; // @[MonteCarlo.scala 52:24 95:{25,33}]
  wire [2:0] _GEN_38 = 3'h5 == state_1 ? _GEN_37 : state_1; // @[MonteCarlo.scala 66:19 52:24]
  wire [31:0] _GEN_39 = 3'h4 == state_1 ? $signed(_price_T_5) : $signed(price_1); // @[MonteCarlo.scala 66:19 86:15 57:27]
  wire [2:0] _GEN_40 = 3'h4 == state_1 ? _GEN_35 : _GEN_38; // @[MonteCarlo.scala 66:19]
  wire [31:0] _GEN_41 = 3'h4 == state_1 ? _GEN_36 : counter_1; // @[MonteCarlo.scala 66:19 62:22]
  wire [51:0] _GEN_74 = {$signed(partial_res3_1), 20'h0}; // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [63:0] _GEN_42 = 3'h3 == state_1 ? $signed(_partial_res3_T_1) : $signed({{12{_GEN_74[51]}},_GEN_74}); // @[MonteCarlo.scala 66:19 82:22 60:27]
  wire [2:0] _GEN_43 = 3'h3 == state_1 ? 3'h4 : _GEN_40; // @[MonteCarlo.scala 66:19 83:22]
  wire [51:0] _GEN_75 = {$signed(partial_res1_1), 20'h0}; // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_46 = 3'h2 == state_1 ? $signed(_partial_res1_T_1) : $signed({{12{_GEN_75[51]}},_GEN_75}); // @[MonteCarlo.scala 66:19 77:22 58:27]
  wire [63:0] _GEN_76 = {$signed(partial_res2_1), 32'h0}; // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [83:0] _GEN_47 = 3'h2 == state_1 ? $signed(_partial_res2_T_1) : $signed({{20{_GEN_76[63]}},_GEN_76}); // @[MonteCarlo.scala 66:19 78:22 59:27]
  wire [63:0] _GEN_49 = 3'h2 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_42); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_55 = 3'h1 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_46); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_56 = 3'h1 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_47); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_57 = 3'h1 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_49); // @[MonteCarlo.scala 66:19 60:27]
  wire [63:0] _GEN_61 = 3'h0 == state_1 ? $signed({{12{_GEN_75[51]}},_GEN_75}) : $signed(_GEN_55); // @[MonteCarlo.scala 66:19 58:27]
  wire [83:0] _GEN_62 = 3'h0 == state_1 ? $signed({{20{_GEN_76[63]}},_GEN_76}) : $signed(_GEN_56); // @[MonteCarlo.scala 66:19 59:27]
  wire [63:0] _GEN_63 = 3'h0 == state_1 ? $signed({{12{_GEN_74[51]}},_GEN_74}) : $signed(_GEN_57); // @[MonteCarlo.scala 66:19 60:27]
  wire [43:0] _GEN_84 = _GEN_29[63:20];
  wire [51:0] _GEN_86 = _GEN_30[83:32];
  wire [43:0] _GEN_88 = _GEN_31[63:20];
  wire [43:0] _GEN_90 = _GEN_61[63:20];
  wire [51:0] _GEN_92 = _GEN_62[83:32];
  wire [43:0] _GEN_94 = _GEN_63[63:20];
  BoxMuller_15 rng ( // @[MonteCarlo.scala 42:19]
    .clock(rng_clock),
    .reset(rng_reset),
    .io_g1_valid(rng_io_g1_valid),
    .io_g1_bits(rng_io_g1_bits),
    .io_g2_valid(rng_io_g2_valid),
    .io_g2_bits(rng_io_g2_bits)
  );
  assign io_request_0_ready = state == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_request_1_ready = state_1 == 3'h1; // @[MonteCarlo.scala 63:26]
  assign io_response_0_valid = state == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_0_bits = price; // @[MonteCarlo.scala 65:16]
  assign io_response_1_valid = state_1 == 3'h5; // @[MonteCarlo.scala 64:26]
  assign io_response_1_bits = price_1; // @[MonteCarlo.scala 65:16]
  assign rng_clock = clock;
  assign rng_reset = reset;
  always @(posedge clock) begin
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state <= 3'h1;
      end else begin
        state <= 3'h0;
      end
    end else if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_3) begin // @[MonteCarlo.scala 71:23]
        state <= 3'h2;
      end else begin
        state <= 3'h1;
      end
    end else if (3'h2 == state) begin // @[MonteCarlo.scala 66:19]
      state <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state <= _GEN_11;
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c1 <= _c1_T_2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      c2 <= io_request_0_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_3) begin // @[Reg.scala 17:18]
      last_step <= _last_step_T_1; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        price <= io_request_0_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          price <= _GEN_7;
        end
      end
    end
    partial_res1 <= _GEN_84[31:0];
    partial_res2 <= _GEN_86[31:0];
    partial_res3 <= _GEN_88[31:0];
    if (!(3'h0 == state)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state) begin // @[MonteCarlo.scala 66:19]
        counter <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state)) begin // @[MonteCarlo.scala 66:19]
          counter <= _GEN_9;
        end
      end
    end
    if (reset) begin // @[MonteCarlo.scala 52:24]
      state_1 <= 3'h0; // @[MonteCarlo.scala 52:24]
    end else if (3'h0 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (initialized) begin // @[MonteCarlo.scala 68:21]
        state_1 <= 3'h1;
      end else begin
        state_1 <= 3'h0;
      end
    end else if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
      if (_c1_T_7) begin // @[MonteCarlo.scala 71:23]
        state_1 <= 3'h2;
      end else begin
        state_1 <= 3'h1;
      end
    end else if (3'h2 == state_1) begin // @[MonteCarlo.scala 66:19]
      state_1 <= 3'h3; // @[MonteCarlo.scala 79:22]
    end else begin
      state_1 <= _GEN_43;
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c1_1 <= _c1_T_6; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      c2_1 <= io_request_1_bits_coefficient2; // @[Reg.scala 17:22]
    end
    if (_c1_T_7) begin // @[Reg.scala 17:18]
      last_step_1 <= _last_step_T_4; // @[Reg.scala 17:22]
    end
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        price_1 <= io_request_1_bits_start_value; // @[MonteCarlo.scala 72:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          price_1 <= _GEN_39;
        end
      end
    end
    partial_res1_1 <= _GEN_90[31:0];
    partial_res2_1 <= _GEN_92[31:0];
    partial_res3_1 <= _GEN_94[31:0];
    if (!(3'h0 == state_1)) begin // @[MonteCarlo.scala 66:19]
      if (3'h1 == state_1) begin // @[MonteCarlo.scala 66:19]
        counter_1 <= 32'h0; // @[MonteCarlo.scala 73:17]
      end else if (!(3'h2 == state_1)) begin // @[MonteCarlo.scala 66:19]
        if (!(3'h3 == state_1)) begin // @[MonteCarlo.scala 66:19]
          counter_1 <= _GEN_41;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  c1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  c2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_step = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  price = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  partial_res1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  partial_res2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  partial_res3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  counter = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  state_1 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  c1_1 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  c2_1 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_step_1 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  price_1 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  partial_res1_1 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  partial_res2_1 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  partial_res3_1 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  counter_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SkidBuffer(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_time_steps,
  input  [31:0] io_enq_bits_start_value,
  input  [31:0] io_enq_bits_coefficient1,
  input  [31:0] io_enq_bits_coefficient2,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_time_steps,
  output [31:0] io_deq_bits_start_value,
  output [31:0] io_deq_bits_coefficient1,
  output [31:0] io_deq_bits_coefficient2
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] data_buffer_time_steps; // @[MonteCarlo.scala 116:24]
  reg [31:0] data_buffer_start_value; // @[MonteCarlo.scala 116:24]
  reg [31:0] data_buffer_coefficient1; // @[MonteCarlo.scala 116:24]
  reg [31:0] data_buffer_coefficient2; // @[MonteCarlo.scala 116:24]
  reg [31:0] skid_buffer_time_steps; // @[MonteCarlo.scala 117:24]
  reg [31:0] skid_buffer_start_value; // @[MonteCarlo.scala 117:24]
  reg [31:0] skid_buffer_coefficient1; // @[MonteCarlo.scala 117:24]
  reg [31:0] skid_buffer_coefficient2; // @[MonteCarlo.scala 117:24]
  reg [1:0] state; // @[MonteCarlo.scala 122:27]
  wire  _T_1 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _GEN_0 = _T_1 ? 2'h1 : 2'h0; // @[MonteCarlo.scala 129:25 130:20 132:20]
  wire  _T_3 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _GEN_10 = _T_1 ? 2'h2 : 2'h1; // @[MonteCarlo.scala 147:31 150:21 152:20]
  wire [1:0] _GEN_15 = _T_3 & _T_1 ? _GEN_0 : _GEN_10; // @[MonteCarlo.scala 138:40]
  wire [1:0] _GEN_24 = _T_3 ? 2'h1 : 2'h2; // @[MonteCarlo.scala 156:25 159:21 161:20]
  wire [1:0] _GEN_29 = 2'h2 == state ? _GEN_24 : 2'h0; // @[MonteCarlo.scala 127:17]
  wire [1:0] _GEN_34 = 2'h1 == state ? _GEN_15 : _GEN_29; // @[MonteCarlo.scala 127:17]
  wire [1:0] state_next = 2'h0 == state ? _GEN_0 : _GEN_34; // @[MonteCarlo.scala 127:17]
  reg  io_enq_ready_REG; // @[MonteCarlo.scala 124:26]
  reg  io_deq_valid_REG; // @[MonteCarlo.scala 125:26]
  assign io_enq_ready = io_enq_ready_REG; // @[MonteCarlo.scala 124:16]
  assign io_deq_valid = io_deq_valid_REG; // @[MonteCarlo.scala 125:16]
  assign io_deq_bits_time_steps = skid_buffer_time_steps; // @[MonteCarlo.scala 166:15]
  assign io_deq_bits_start_value = skid_buffer_start_value; // @[MonteCarlo.scala 166:15]
  assign io_deq_bits_coefficient1 = skid_buffer_coefficient1; // @[MonteCarlo.scala 166:15]
  assign io_deq_bits_coefficient2 = skid_buffer_coefficient2; // @[MonteCarlo.scala 166:15]
  always @(posedge clock) begin
    if (!(2'h0 == state)) begin // @[MonteCarlo.scala 127:17]
      if (2'h1 == state) begin // @[MonteCarlo.scala 127:17]
        if (!(_T_3 & _T_1)) begin // @[MonteCarlo.scala 138:40]
          if (_T_1) begin // @[MonteCarlo.scala 147:31]
            data_buffer_time_steps <= io_enq_bits_time_steps; // @[MonteCarlo.scala 149:21]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[MonteCarlo.scala 127:17]
      if (2'h1 == state) begin // @[MonteCarlo.scala 127:17]
        if (!(_T_3 & _T_1)) begin // @[MonteCarlo.scala 138:40]
          if (_T_1) begin // @[MonteCarlo.scala 147:31]
            data_buffer_start_value <= io_enq_bits_start_value; // @[MonteCarlo.scala 149:21]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[MonteCarlo.scala 127:17]
      if (2'h1 == state) begin // @[MonteCarlo.scala 127:17]
        if (!(_T_3 & _T_1)) begin // @[MonteCarlo.scala 138:40]
          if (_T_1) begin // @[MonteCarlo.scala 147:31]
            data_buffer_coefficient1 <= io_enq_bits_coefficient1; // @[MonteCarlo.scala 149:21]
          end
        end
      end
    end
    if (!(2'h0 == state)) begin // @[MonteCarlo.scala 127:17]
      if (2'h1 == state) begin // @[MonteCarlo.scala 127:17]
        if (!(_T_3 & _T_1)) begin // @[MonteCarlo.scala 138:40]
          if (_T_1) begin // @[MonteCarlo.scala 147:31]
            data_buffer_coefficient2 <= io_enq_bits_coefficient2; // @[MonteCarlo.scala 149:21]
          end
        end
      end
    end
    if (2'h0 == state) begin // @[MonteCarlo.scala 127:17]
      skid_buffer_time_steps <= io_enq_bits_time_steps; // @[MonteCarlo.scala 135:19]
    end else if (2'h1 == state) begin // @[MonteCarlo.scala 127:17]
      if (_T_3 & _T_1) begin // @[MonteCarlo.scala 138:40]
        if (_T_1) begin // @[MonteCarlo.scala 139:27]
          skid_buffer_time_steps <= io_enq_bits_time_steps; // @[MonteCarlo.scala 141:23]
        end
      end
    end else if (2'h2 == state) begin // @[MonteCarlo.scala 127:17]
      if (_T_3) begin // @[MonteCarlo.scala 156:25]
        skid_buffer_time_steps <= data_buffer_time_steps; // @[MonteCarlo.scala 158:21]
      end
    end
    if (2'h0 == state) begin // @[MonteCarlo.scala 127:17]
      skid_buffer_start_value <= io_enq_bits_start_value; // @[MonteCarlo.scala 135:19]
    end else if (2'h1 == state) begin // @[MonteCarlo.scala 127:17]
      if (_T_3 & _T_1) begin // @[MonteCarlo.scala 138:40]
        if (_T_1) begin // @[MonteCarlo.scala 139:27]
          skid_buffer_start_value <= io_enq_bits_start_value; // @[MonteCarlo.scala 141:23]
        end
      end
    end else if (2'h2 == state) begin // @[MonteCarlo.scala 127:17]
      if (_T_3) begin // @[MonteCarlo.scala 156:25]
        skid_buffer_start_value <= data_buffer_start_value; // @[MonteCarlo.scala 158:21]
      end
    end
    if (2'h0 == state) begin // @[MonteCarlo.scala 127:17]
      skid_buffer_coefficient1 <= io_enq_bits_coefficient1; // @[MonteCarlo.scala 135:19]
    end else if (2'h1 == state) begin // @[MonteCarlo.scala 127:17]
      if (_T_3 & _T_1) begin // @[MonteCarlo.scala 138:40]
        if (_T_1) begin // @[MonteCarlo.scala 139:27]
          skid_buffer_coefficient1 <= io_enq_bits_coefficient1; // @[MonteCarlo.scala 141:23]
        end
      end
    end else if (2'h2 == state) begin // @[MonteCarlo.scala 127:17]
      if (_T_3) begin // @[MonteCarlo.scala 156:25]
        skid_buffer_coefficient1 <= data_buffer_coefficient1; // @[MonteCarlo.scala 158:21]
      end
    end
    if (2'h0 == state) begin // @[MonteCarlo.scala 127:17]
      skid_buffer_coefficient2 <= io_enq_bits_coefficient2; // @[MonteCarlo.scala 135:19]
    end else if (2'h1 == state) begin // @[MonteCarlo.scala 127:17]
      if (_T_3 & _T_1) begin // @[MonteCarlo.scala 138:40]
        if (_T_1) begin // @[MonteCarlo.scala 139:27]
          skid_buffer_coefficient2 <= io_enq_bits_coefficient2; // @[MonteCarlo.scala 141:23]
        end
      end
    end else if (2'h2 == state) begin // @[MonteCarlo.scala 127:17]
      if (_T_3) begin // @[MonteCarlo.scala 156:25]
        skid_buffer_coefficient2 <= data_buffer_coefficient2; // @[MonteCarlo.scala 158:21]
      end
    end
    if (reset) begin // @[MonteCarlo.scala 122:27]
      state <= 2'h0; // @[MonteCarlo.scala 122:27]
    end else if (2'h0 == state) begin // @[MonteCarlo.scala 127:17]
      state <= _GEN_0;
    end else if (2'h1 == state) begin // @[MonteCarlo.scala 127:17]
      if (_T_3 & _T_1) begin // @[MonteCarlo.scala 138:40]
        state <= _GEN_0;
      end else begin
        state <= _GEN_10;
      end
    end else if (2'h2 == state) begin // @[MonteCarlo.scala 127:17]
      state <= _GEN_24;
    end else begin
      state <= 2'h0;
    end
    io_enq_ready_REG <= reset | state_next != 2'h2; // @[MonteCarlo.scala 124:{26,26,26}]
    if (reset) begin // @[MonteCarlo.scala 125:26]
      io_deq_valid_REG <= 1'h0; // @[MonteCarlo.scala 125:26]
    end else begin
      io_deq_valid_REG <= state_next != 2'h0; // @[MonteCarlo.scala 125:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_buffer_time_steps = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  data_buffer_start_value = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  data_buffer_coefficient1 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  data_buffer_coefficient2 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  skid_buffer_time_steps = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  skid_buffer_start_value = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  skid_buffer_coefficient1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  skid_buffer_coefficient2 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  state = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  io_enq_ready_REG = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  io_deq_valid_REG = _RAND_10[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SkidBuffer_62(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] data_buffer; // @[MonteCarlo.scala 116:24]
  reg [31:0] skid_buffer; // @[MonteCarlo.scala 117:24]
  reg [1:0] state; // @[MonteCarlo.scala 122:27]
  wire  _T_1 = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _GEN_0 = _T_1 ? 2'h1 : 2'h0; // @[MonteCarlo.scala 129:25 130:20 132:20]
  wire  _T_3 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _GEN_4 = _T_1 ? 2'h2 : 2'h1; // @[MonteCarlo.scala 147:31 150:21 152:20]
  wire [1:0] _GEN_6 = _T_3 & _T_1 ? _GEN_0 : _GEN_4; // @[MonteCarlo.scala 138:40]
  wire [1:0] _GEN_9 = _T_3 ? 2'h1 : 2'h2; // @[MonteCarlo.scala 156:25 159:21 161:20]
  wire [1:0] _GEN_11 = 2'h2 == state ? _GEN_9 : 2'h0; // @[MonteCarlo.scala 127:17]
  wire [1:0] _GEN_13 = 2'h1 == state ? _GEN_6 : _GEN_11; // @[MonteCarlo.scala 127:17]
  wire [1:0] state_next = 2'h0 == state ? _GEN_0 : _GEN_13; // @[MonteCarlo.scala 127:17]
  reg  io_enq_ready_REG; // @[MonteCarlo.scala 124:26]
  reg  io_deq_valid_REG; // @[MonteCarlo.scala 125:26]
  assign io_enq_ready = io_enq_ready_REG; // @[MonteCarlo.scala 124:16]
  assign io_deq_valid = io_deq_valid_REG; // @[MonteCarlo.scala 125:16]
  assign io_deq_bits = skid_buffer; // @[MonteCarlo.scala 166:15]
  always @(posedge clock) begin
    if (!(2'h0 == state)) begin // @[MonteCarlo.scala 127:17]
      if (2'h1 == state) begin // @[MonteCarlo.scala 127:17]
        if (!(_T_3 & _T_1)) begin // @[MonteCarlo.scala 138:40]
          if (_T_1) begin // @[MonteCarlo.scala 147:31]
            data_buffer <= io_enq_bits; // @[MonteCarlo.scala 149:21]
          end
        end
      end
    end
    if (2'h0 == state) begin // @[MonteCarlo.scala 127:17]
      skid_buffer <= io_enq_bits; // @[MonteCarlo.scala 135:19]
    end else if (2'h1 == state) begin // @[MonteCarlo.scala 127:17]
      if (_T_3 & _T_1) begin // @[MonteCarlo.scala 138:40]
        if (_T_1) begin // @[MonteCarlo.scala 139:27]
          skid_buffer <= io_enq_bits; // @[MonteCarlo.scala 141:23]
        end
      end
    end else if (2'h2 == state) begin // @[MonteCarlo.scala 127:17]
      if (_T_3) begin // @[MonteCarlo.scala 156:25]
        skid_buffer <= data_buffer; // @[MonteCarlo.scala 158:21]
      end
    end
    if (reset) begin // @[MonteCarlo.scala 122:27]
      state <= 2'h0; // @[MonteCarlo.scala 122:27]
    end else if (2'h0 == state) begin // @[MonteCarlo.scala 127:17]
      state <= _GEN_0;
    end else if (2'h1 == state) begin // @[MonteCarlo.scala 127:17]
      if (_T_3 & _T_1) begin // @[MonteCarlo.scala 138:40]
        state <= _GEN_0;
      end else begin
        state <= _GEN_4;
      end
    end else if (2'h2 == state) begin // @[MonteCarlo.scala 127:17]
      state <= _GEN_9;
    end else begin
      state <= 2'h0;
    end
    io_enq_ready_REG <= reset | state_next != 2'h2; // @[MonteCarlo.scala 124:{26,26,26}]
    if (reset) begin // @[MonteCarlo.scala 125:26]
      io_deq_valid_REG <= 1'h0; // @[MonteCarlo.scala 125:26]
    end else begin
      io_deq_valid_REG <= state_next != 2'h0; // @[MonteCarlo.scala 125:26]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  data_buffer = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  skid_buffer = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  io_enq_ready_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_deq_valid_REG = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PipelinedMean(
  input         clock,
  input         reset,
  output        io_lanes_0_ready,
  input         io_lanes_0_valid,
  input  [31:0] io_lanes_0_bits,
  output        io_lanes_1_ready,
  input         io_lanes_1_valid,
  input  [31:0] io_lanes_1_bits,
  output        io_lanes_2_ready,
  input         io_lanes_2_valid,
  input  [31:0] io_lanes_2_bits,
  output        io_lanes_3_ready,
  input         io_lanes_3_valid,
  input  [31:0] io_lanes_3_bits,
  output        io_lanes_4_ready,
  input         io_lanes_4_valid,
  input  [31:0] io_lanes_4_bits,
  output        io_lanes_5_ready,
  input         io_lanes_5_valid,
  input  [31:0] io_lanes_5_bits,
  output        io_lanes_6_ready,
  input         io_lanes_6_valid,
  input  [31:0] io_lanes_6_bits,
  output        io_lanes_7_ready,
  input         io_lanes_7_valid,
  input  [31:0] io_lanes_7_bits,
  output        io_lanes_8_ready,
  input         io_lanes_8_valid,
  input  [31:0] io_lanes_8_bits,
  output        io_lanes_9_ready,
  input         io_lanes_9_valid,
  input  [31:0] io_lanes_9_bits,
  output        io_lanes_10_ready,
  input         io_lanes_10_valid,
  input  [31:0] io_lanes_10_bits,
  output        io_lanes_11_ready,
  input         io_lanes_11_valid,
  input  [31:0] io_lanes_11_bits,
  output        io_lanes_12_ready,
  input         io_lanes_12_valid,
  input  [31:0] io_lanes_12_bits,
  output        io_lanes_13_ready,
  input         io_lanes_13_valid,
  input  [31:0] io_lanes_13_bits,
  output        io_lanes_14_ready,
  input         io_lanes_14_valid,
  input  [31:0] io_lanes_14_bits,
  output        io_lanes_15_ready,
  input         io_lanes_15_valid,
  input  [31:0] io_lanes_15_bits,
  output        io_lanes_16_ready,
  input         io_lanes_16_valid,
  input  [31:0] io_lanes_16_bits,
  output        io_lanes_17_ready,
  input         io_lanes_17_valid,
  input  [31:0] io_lanes_17_bits,
  output        io_lanes_18_ready,
  input         io_lanes_18_valid,
  input  [31:0] io_lanes_18_bits,
  output        io_lanes_19_ready,
  input         io_lanes_19_valid,
  input  [31:0] io_lanes_19_bits,
  output        io_lanes_20_ready,
  input         io_lanes_20_valid,
  input  [31:0] io_lanes_20_bits,
  output        io_lanes_21_ready,
  input         io_lanes_21_valid,
  input  [31:0] io_lanes_21_bits,
  output        io_lanes_22_ready,
  input         io_lanes_22_valid,
  input  [31:0] io_lanes_22_bits,
  output        io_lanes_23_ready,
  input         io_lanes_23_valid,
  input  [31:0] io_lanes_23_bits,
  output        io_lanes_24_ready,
  input         io_lanes_24_valid,
  input  [31:0] io_lanes_24_bits,
  output        io_lanes_25_ready,
  input         io_lanes_25_valid,
  input  [31:0] io_lanes_25_bits,
  output        io_lanes_26_ready,
  input         io_lanes_26_valid,
  input  [31:0] io_lanes_26_bits,
  output        io_lanes_27_ready,
  input         io_lanes_27_valid,
  input  [31:0] io_lanes_27_bits,
  output        io_lanes_28_ready,
  input         io_lanes_28_valid,
  input  [31:0] io_lanes_28_bits,
  output        io_lanes_29_ready,
  input         io_lanes_29_valid,
  input  [31:0] io_lanes_29_bits,
  output        io_lanes_30_ready,
  input         io_lanes_30_valid,
  input  [31:0] io_lanes_30_bits,
  output        io_lanes_31_ready,
  input         io_lanes_31_valid,
  input  [31:0] io_lanes_31_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
  wire  io_result_next_b_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_1_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_1_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_1_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_1_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_1_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_1_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_1_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_1_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_2_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_2_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_2_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_2_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_2_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_2_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_2_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_2_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_3_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_3_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_3_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_3_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_3_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_3_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_3_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_3_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_4_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_4_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_4_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_4_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_4_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_4_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_4_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_4_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_5_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_5_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_5_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_5_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_5_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_5_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_5_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_5_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_6_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_6_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_6_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_6_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_6_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_6_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_6_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_6_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_7_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_7_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_7_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_7_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_7_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_7_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_7_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_7_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_8_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_8_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_8_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_8_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_8_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_8_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_8_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_8_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_9_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_9_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_9_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_9_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_9_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_9_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_9_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_9_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_10_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_10_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_10_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_10_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_10_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_10_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_10_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_10_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_11_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_11_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_11_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_11_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_11_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_11_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_11_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_11_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_12_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_12_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_12_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_12_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_12_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_12_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_12_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_12_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_13_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_13_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_13_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_13_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_13_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_13_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_13_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_13_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_14_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_14_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_14_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_14_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_14_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_14_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_14_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_14_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_15_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_15_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_15_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_15_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_15_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_15_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_15_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_15_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_16_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_16_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_16_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_16_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_16_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_16_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_16_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_16_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_17_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_17_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_17_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_17_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_17_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_17_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_17_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_17_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_18_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_18_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_18_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_18_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_18_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_18_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_18_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_18_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_19_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_19_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_19_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_19_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_19_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_19_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_19_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_19_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_20_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_20_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_20_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_20_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_20_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_20_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_20_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_20_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_21_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_21_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_21_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_21_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_21_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_21_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_21_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_21_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_22_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_22_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_22_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_22_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_22_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_22_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_22_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_22_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_23_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_23_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_23_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_23_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_23_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_23_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_23_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_23_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_24_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_24_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_24_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_24_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_24_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_24_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_24_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_24_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_25_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_25_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_25_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_25_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_25_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_25_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_25_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_25_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_26_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_26_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_26_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_26_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_26_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_26_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_26_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_26_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_27_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_27_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_27_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_27_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_27_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_27_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_27_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_27_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_28_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_28_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_28_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_28_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_28_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_28_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_28_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_28_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_29_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_29_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_29_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_29_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_29_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_29_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_29_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_29_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_30_clock; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_30_reset; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_30_io_enq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_30_io_enq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_30_io_enq_bits; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_30_io_deq_ready; // @[MonteCarlo.scala 191:25]
  wire  io_result_next_b_30_io_deq_valid; // @[MonteCarlo.scala 191:25]
  wire [31:0] io_result_next_b_30_io_deq_bits; // @[MonteCarlo.scala 191:25]
  wire [31:0] _io_result_next_r_T_2 = $signed(io_lanes_0_bits) + $signed(io_lanes_1_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r = _io_result_next_r_T_2[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T = io_lanes_0_valid & io_lanes_1_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_5 = $signed(io_lanes_2_bits) + $signed(io_lanes_3_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_1 = _io_result_next_r_T_5[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_1 = io_lanes_2_valid & io_lanes_3_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_8 = $signed(io_lanes_4_bits) + $signed(io_lanes_5_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_2 = _io_result_next_r_T_8[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_2 = io_lanes_4_valid & io_lanes_5_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_11 = $signed(io_lanes_6_bits) + $signed(io_lanes_7_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_3 = _io_result_next_r_T_11[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_3 = io_lanes_6_valid & io_lanes_7_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_14 = $signed(io_lanes_8_bits) + $signed(io_lanes_9_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_4 = _io_result_next_r_T_14[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_4 = io_lanes_8_valid & io_lanes_9_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_17 = $signed(io_lanes_10_bits) + $signed(io_lanes_11_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_5 = _io_result_next_r_T_17[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_5 = io_lanes_10_valid & io_lanes_11_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_20 = $signed(io_lanes_12_bits) + $signed(io_lanes_13_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_6 = _io_result_next_r_T_20[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_6 = io_lanes_12_valid & io_lanes_13_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_23 = $signed(io_lanes_14_bits) + $signed(io_lanes_15_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_7 = _io_result_next_r_T_23[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_7 = io_lanes_14_valid & io_lanes_15_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_26 = $signed(io_lanes_16_bits) + $signed(io_lanes_17_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_8 = _io_result_next_r_T_26[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_8 = io_lanes_16_valid & io_lanes_17_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_29 = $signed(io_lanes_18_bits) + $signed(io_lanes_19_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_9 = _io_result_next_r_T_29[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_9 = io_lanes_18_valid & io_lanes_19_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_32 = $signed(io_lanes_20_bits) + $signed(io_lanes_21_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_10 = _io_result_next_r_T_32[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_10 = io_lanes_20_valid & io_lanes_21_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_35 = $signed(io_lanes_22_bits) + $signed(io_lanes_23_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_11 = _io_result_next_r_T_35[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_11 = io_lanes_22_valid & io_lanes_23_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_38 = $signed(io_lanes_24_bits) + $signed(io_lanes_25_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_12 = _io_result_next_r_T_38[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_12 = io_lanes_24_valid & io_lanes_25_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_41 = $signed(io_lanes_26_bits) + $signed(io_lanes_27_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_13 = _io_result_next_r_T_41[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_13 = io_lanes_26_valid & io_lanes_27_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_44 = $signed(io_lanes_28_bits) + $signed(io_lanes_29_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_14 = _io_result_next_r_T_44[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_14 = io_lanes_28_valid & io_lanes_29_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_47 = $signed(io_lanes_30_bits) + $signed(io_lanes_31_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_15 = _io_result_next_r_T_47[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_15 = io_lanes_30_valid & io_lanes_31_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_50 = $signed(io_result_next_b_io_deq_bits) + $signed(io_result_next_b_1_io_deq_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_16 = _io_result_next_r_T_50[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_16 = io_result_next_b_io_deq_valid & io_result_next_b_1_io_deq_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_53 = $signed(io_result_next_b_2_io_deq_bits) + $signed(io_result_next_b_3_io_deq_bits)
    ; // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_17 = _io_result_next_r_T_53[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_17 = io_result_next_b_2_io_deq_valid & io_result_next_b_3_io_deq_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_56 = $signed(io_result_next_b_4_io_deq_bits) + $signed(io_result_next_b_5_io_deq_bits)
    ; // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_18 = _io_result_next_r_T_56[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_18 = io_result_next_b_4_io_deq_valid & io_result_next_b_5_io_deq_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_59 = $signed(io_result_next_b_6_io_deq_bits) + $signed(io_result_next_b_7_io_deq_bits)
    ; // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_19 = _io_result_next_r_T_59[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_19 = io_result_next_b_6_io_deq_valid & io_result_next_b_7_io_deq_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_62 = $signed(io_result_next_b_8_io_deq_bits) + $signed(io_result_next_b_9_io_deq_bits)
    ; // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_20 = _io_result_next_r_T_62[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_20 = io_result_next_b_8_io_deq_valid & io_result_next_b_9_io_deq_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_65 = $signed(io_result_next_b_10_io_deq_bits) + $signed(
    io_result_next_b_11_io_deq_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_21 = _io_result_next_r_T_65[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_21 = io_result_next_b_10_io_deq_valid & io_result_next_b_11_io_deq_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_68 = $signed(io_result_next_b_12_io_deq_bits) + $signed(
    io_result_next_b_13_io_deq_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_22 = _io_result_next_r_T_68[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_22 = io_result_next_b_12_io_deq_valid & io_result_next_b_13_io_deq_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_71 = $signed(io_result_next_b_14_io_deq_bits) + $signed(
    io_result_next_b_15_io_deq_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_23 = _io_result_next_r_T_71[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_23 = io_result_next_b_14_io_deq_valid & io_result_next_b_15_io_deq_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_74 = $signed(io_result_next_b_16_io_deq_bits) + $signed(
    io_result_next_b_17_io_deq_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_24 = _io_result_next_r_T_74[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_24 = io_result_next_b_16_io_deq_valid & io_result_next_b_17_io_deq_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_77 = $signed(io_result_next_b_18_io_deq_bits) + $signed(
    io_result_next_b_19_io_deq_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_25 = _io_result_next_r_T_77[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_25 = io_result_next_b_18_io_deq_valid & io_result_next_b_19_io_deq_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_80 = $signed(io_result_next_b_20_io_deq_bits) + $signed(
    io_result_next_b_21_io_deq_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_26 = _io_result_next_r_T_80[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_26 = io_result_next_b_20_io_deq_valid & io_result_next_b_21_io_deq_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_83 = $signed(io_result_next_b_22_io_deq_bits) + $signed(
    io_result_next_b_23_io_deq_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_27 = _io_result_next_r_T_83[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_27 = io_result_next_b_22_io_deq_valid & io_result_next_b_23_io_deq_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_86 = $signed(io_result_next_b_24_io_deq_bits) + $signed(
    io_result_next_b_25_io_deq_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_28 = _io_result_next_r_T_86[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_28 = io_result_next_b_24_io_deq_valid & io_result_next_b_25_io_deq_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_89 = $signed(io_result_next_b_26_io_deq_bits) + $signed(
    io_result_next_b_27_io_deq_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_29 = _io_result_next_r_T_89[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_29 = io_result_next_b_26_io_deq_valid & io_result_next_b_27_io_deq_valid; // @[MonteCarlo.scala 193:42]
  wire [31:0] _io_result_next_r_T_92 = $signed(io_result_next_b_28_io_deq_bits) + $signed(
    io_result_next_b_29_io_deq_bits); // @[MonteCarlo.scala 190:32]
  wire [30:0] io_result_next_r_30 = _io_result_next_r_T_92[31:1]; // @[MonteCarlo.scala 190:47]
  wire  _io_result_next_b_io_enq_valid_T_30 = io_result_next_b_28_io_deq_valid & io_result_next_b_29_io_deq_valid; // @[MonteCarlo.scala 193:42]
  SkidBuffer_62 io_result_next_b ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_clock),
    .reset(io_result_next_b_reset),
    .io_enq_ready(io_result_next_b_io_enq_ready),
    .io_enq_valid(io_result_next_b_io_enq_valid),
    .io_enq_bits(io_result_next_b_io_enq_bits),
    .io_deq_ready(io_result_next_b_io_deq_ready),
    .io_deq_valid(io_result_next_b_io_deq_valid),
    .io_deq_bits(io_result_next_b_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_1 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_1_clock),
    .reset(io_result_next_b_1_reset),
    .io_enq_ready(io_result_next_b_1_io_enq_ready),
    .io_enq_valid(io_result_next_b_1_io_enq_valid),
    .io_enq_bits(io_result_next_b_1_io_enq_bits),
    .io_deq_ready(io_result_next_b_1_io_deq_ready),
    .io_deq_valid(io_result_next_b_1_io_deq_valid),
    .io_deq_bits(io_result_next_b_1_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_2 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_2_clock),
    .reset(io_result_next_b_2_reset),
    .io_enq_ready(io_result_next_b_2_io_enq_ready),
    .io_enq_valid(io_result_next_b_2_io_enq_valid),
    .io_enq_bits(io_result_next_b_2_io_enq_bits),
    .io_deq_ready(io_result_next_b_2_io_deq_ready),
    .io_deq_valid(io_result_next_b_2_io_deq_valid),
    .io_deq_bits(io_result_next_b_2_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_3 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_3_clock),
    .reset(io_result_next_b_3_reset),
    .io_enq_ready(io_result_next_b_3_io_enq_ready),
    .io_enq_valid(io_result_next_b_3_io_enq_valid),
    .io_enq_bits(io_result_next_b_3_io_enq_bits),
    .io_deq_ready(io_result_next_b_3_io_deq_ready),
    .io_deq_valid(io_result_next_b_3_io_deq_valid),
    .io_deq_bits(io_result_next_b_3_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_4 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_4_clock),
    .reset(io_result_next_b_4_reset),
    .io_enq_ready(io_result_next_b_4_io_enq_ready),
    .io_enq_valid(io_result_next_b_4_io_enq_valid),
    .io_enq_bits(io_result_next_b_4_io_enq_bits),
    .io_deq_ready(io_result_next_b_4_io_deq_ready),
    .io_deq_valid(io_result_next_b_4_io_deq_valid),
    .io_deq_bits(io_result_next_b_4_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_5 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_5_clock),
    .reset(io_result_next_b_5_reset),
    .io_enq_ready(io_result_next_b_5_io_enq_ready),
    .io_enq_valid(io_result_next_b_5_io_enq_valid),
    .io_enq_bits(io_result_next_b_5_io_enq_bits),
    .io_deq_ready(io_result_next_b_5_io_deq_ready),
    .io_deq_valid(io_result_next_b_5_io_deq_valid),
    .io_deq_bits(io_result_next_b_5_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_6 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_6_clock),
    .reset(io_result_next_b_6_reset),
    .io_enq_ready(io_result_next_b_6_io_enq_ready),
    .io_enq_valid(io_result_next_b_6_io_enq_valid),
    .io_enq_bits(io_result_next_b_6_io_enq_bits),
    .io_deq_ready(io_result_next_b_6_io_deq_ready),
    .io_deq_valid(io_result_next_b_6_io_deq_valid),
    .io_deq_bits(io_result_next_b_6_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_7 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_7_clock),
    .reset(io_result_next_b_7_reset),
    .io_enq_ready(io_result_next_b_7_io_enq_ready),
    .io_enq_valid(io_result_next_b_7_io_enq_valid),
    .io_enq_bits(io_result_next_b_7_io_enq_bits),
    .io_deq_ready(io_result_next_b_7_io_deq_ready),
    .io_deq_valid(io_result_next_b_7_io_deq_valid),
    .io_deq_bits(io_result_next_b_7_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_8 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_8_clock),
    .reset(io_result_next_b_8_reset),
    .io_enq_ready(io_result_next_b_8_io_enq_ready),
    .io_enq_valid(io_result_next_b_8_io_enq_valid),
    .io_enq_bits(io_result_next_b_8_io_enq_bits),
    .io_deq_ready(io_result_next_b_8_io_deq_ready),
    .io_deq_valid(io_result_next_b_8_io_deq_valid),
    .io_deq_bits(io_result_next_b_8_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_9 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_9_clock),
    .reset(io_result_next_b_9_reset),
    .io_enq_ready(io_result_next_b_9_io_enq_ready),
    .io_enq_valid(io_result_next_b_9_io_enq_valid),
    .io_enq_bits(io_result_next_b_9_io_enq_bits),
    .io_deq_ready(io_result_next_b_9_io_deq_ready),
    .io_deq_valid(io_result_next_b_9_io_deq_valid),
    .io_deq_bits(io_result_next_b_9_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_10 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_10_clock),
    .reset(io_result_next_b_10_reset),
    .io_enq_ready(io_result_next_b_10_io_enq_ready),
    .io_enq_valid(io_result_next_b_10_io_enq_valid),
    .io_enq_bits(io_result_next_b_10_io_enq_bits),
    .io_deq_ready(io_result_next_b_10_io_deq_ready),
    .io_deq_valid(io_result_next_b_10_io_deq_valid),
    .io_deq_bits(io_result_next_b_10_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_11 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_11_clock),
    .reset(io_result_next_b_11_reset),
    .io_enq_ready(io_result_next_b_11_io_enq_ready),
    .io_enq_valid(io_result_next_b_11_io_enq_valid),
    .io_enq_bits(io_result_next_b_11_io_enq_bits),
    .io_deq_ready(io_result_next_b_11_io_deq_ready),
    .io_deq_valid(io_result_next_b_11_io_deq_valid),
    .io_deq_bits(io_result_next_b_11_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_12 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_12_clock),
    .reset(io_result_next_b_12_reset),
    .io_enq_ready(io_result_next_b_12_io_enq_ready),
    .io_enq_valid(io_result_next_b_12_io_enq_valid),
    .io_enq_bits(io_result_next_b_12_io_enq_bits),
    .io_deq_ready(io_result_next_b_12_io_deq_ready),
    .io_deq_valid(io_result_next_b_12_io_deq_valid),
    .io_deq_bits(io_result_next_b_12_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_13 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_13_clock),
    .reset(io_result_next_b_13_reset),
    .io_enq_ready(io_result_next_b_13_io_enq_ready),
    .io_enq_valid(io_result_next_b_13_io_enq_valid),
    .io_enq_bits(io_result_next_b_13_io_enq_bits),
    .io_deq_ready(io_result_next_b_13_io_deq_ready),
    .io_deq_valid(io_result_next_b_13_io_deq_valid),
    .io_deq_bits(io_result_next_b_13_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_14 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_14_clock),
    .reset(io_result_next_b_14_reset),
    .io_enq_ready(io_result_next_b_14_io_enq_ready),
    .io_enq_valid(io_result_next_b_14_io_enq_valid),
    .io_enq_bits(io_result_next_b_14_io_enq_bits),
    .io_deq_ready(io_result_next_b_14_io_deq_ready),
    .io_deq_valid(io_result_next_b_14_io_deq_valid),
    .io_deq_bits(io_result_next_b_14_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_15 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_15_clock),
    .reset(io_result_next_b_15_reset),
    .io_enq_ready(io_result_next_b_15_io_enq_ready),
    .io_enq_valid(io_result_next_b_15_io_enq_valid),
    .io_enq_bits(io_result_next_b_15_io_enq_bits),
    .io_deq_ready(io_result_next_b_15_io_deq_ready),
    .io_deq_valid(io_result_next_b_15_io_deq_valid),
    .io_deq_bits(io_result_next_b_15_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_16 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_16_clock),
    .reset(io_result_next_b_16_reset),
    .io_enq_ready(io_result_next_b_16_io_enq_ready),
    .io_enq_valid(io_result_next_b_16_io_enq_valid),
    .io_enq_bits(io_result_next_b_16_io_enq_bits),
    .io_deq_ready(io_result_next_b_16_io_deq_ready),
    .io_deq_valid(io_result_next_b_16_io_deq_valid),
    .io_deq_bits(io_result_next_b_16_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_17 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_17_clock),
    .reset(io_result_next_b_17_reset),
    .io_enq_ready(io_result_next_b_17_io_enq_ready),
    .io_enq_valid(io_result_next_b_17_io_enq_valid),
    .io_enq_bits(io_result_next_b_17_io_enq_bits),
    .io_deq_ready(io_result_next_b_17_io_deq_ready),
    .io_deq_valid(io_result_next_b_17_io_deq_valid),
    .io_deq_bits(io_result_next_b_17_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_18 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_18_clock),
    .reset(io_result_next_b_18_reset),
    .io_enq_ready(io_result_next_b_18_io_enq_ready),
    .io_enq_valid(io_result_next_b_18_io_enq_valid),
    .io_enq_bits(io_result_next_b_18_io_enq_bits),
    .io_deq_ready(io_result_next_b_18_io_deq_ready),
    .io_deq_valid(io_result_next_b_18_io_deq_valid),
    .io_deq_bits(io_result_next_b_18_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_19 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_19_clock),
    .reset(io_result_next_b_19_reset),
    .io_enq_ready(io_result_next_b_19_io_enq_ready),
    .io_enq_valid(io_result_next_b_19_io_enq_valid),
    .io_enq_bits(io_result_next_b_19_io_enq_bits),
    .io_deq_ready(io_result_next_b_19_io_deq_ready),
    .io_deq_valid(io_result_next_b_19_io_deq_valid),
    .io_deq_bits(io_result_next_b_19_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_20 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_20_clock),
    .reset(io_result_next_b_20_reset),
    .io_enq_ready(io_result_next_b_20_io_enq_ready),
    .io_enq_valid(io_result_next_b_20_io_enq_valid),
    .io_enq_bits(io_result_next_b_20_io_enq_bits),
    .io_deq_ready(io_result_next_b_20_io_deq_ready),
    .io_deq_valid(io_result_next_b_20_io_deq_valid),
    .io_deq_bits(io_result_next_b_20_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_21 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_21_clock),
    .reset(io_result_next_b_21_reset),
    .io_enq_ready(io_result_next_b_21_io_enq_ready),
    .io_enq_valid(io_result_next_b_21_io_enq_valid),
    .io_enq_bits(io_result_next_b_21_io_enq_bits),
    .io_deq_ready(io_result_next_b_21_io_deq_ready),
    .io_deq_valid(io_result_next_b_21_io_deq_valid),
    .io_deq_bits(io_result_next_b_21_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_22 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_22_clock),
    .reset(io_result_next_b_22_reset),
    .io_enq_ready(io_result_next_b_22_io_enq_ready),
    .io_enq_valid(io_result_next_b_22_io_enq_valid),
    .io_enq_bits(io_result_next_b_22_io_enq_bits),
    .io_deq_ready(io_result_next_b_22_io_deq_ready),
    .io_deq_valid(io_result_next_b_22_io_deq_valid),
    .io_deq_bits(io_result_next_b_22_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_23 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_23_clock),
    .reset(io_result_next_b_23_reset),
    .io_enq_ready(io_result_next_b_23_io_enq_ready),
    .io_enq_valid(io_result_next_b_23_io_enq_valid),
    .io_enq_bits(io_result_next_b_23_io_enq_bits),
    .io_deq_ready(io_result_next_b_23_io_deq_ready),
    .io_deq_valid(io_result_next_b_23_io_deq_valid),
    .io_deq_bits(io_result_next_b_23_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_24 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_24_clock),
    .reset(io_result_next_b_24_reset),
    .io_enq_ready(io_result_next_b_24_io_enq_ready),
    .io_enq_valid(io_result_next_b_24_io_enq_valid),
    .io_enq_bits(io_result_next_b_24_io_enq_bits),
    .io_deq_ready(io_result_next_b_24_io_deq_ready),
    .io_deq_valid(io_result_next_b_24_io_deq_valid),
    .io_deq_bits(io_result_next_b_24_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_25 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_25_clock),
    .reset(io_result_next_b_25_reset),
    .io_enq_ready(io_result_next_b_25_io_enq_ready),
    .io_enq_valid(io_result_next_b_25_io_enq_valid),
    .io_enq_bits(io_result_next_b_25_io_enq_bits),
    .io_deq_ready(io_result_next_b_25_io_deq_ready),
    .io_deq_valid(io_result_next_b_25_io_deq_valid),
    .io_deq_bits(io_result_next_b_25_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_26 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_26_clock),
    .reset(io_result_next_b_26_reset),
    .io_enq_ready(io_result_next_b_26_io_enq_ready),
    .io_enq_valid(io_result_next_b_26_io_enq_valid),
    .io_enq_bits(io_result_next_b_26_io_enq_bits),
    .io_deq_ready(io_result_next_b_26_io_deq_ready),
    .io_deq_valid(io_result_next_b_26_io_deq_valid),
    .io_deq_bits(io_result_next_b_26_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_27 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_27_clock),
    .reset(io_result_next_b_27_reset),
    .io_enq_ready(io_result_next_b_27_io_enq_ready),
    .io_enq_valid(io_result_next_b_27_io_enq_valid),
    .io_enq_bits(io_result_next_b_27_io_enq_bits),
    .io_deq_ready(io_result_next_b_27_io_deq_ready),
    .io_deq_valid(io_result_next_b_27_io_deq_valid),
    .io_deq_bits(io_result_next_b_27_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_28 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_28_clock),
    .reset(io_result_next_b_28_reset),
    .io_enq_ready(io_result_next_b_28_io_enq_ready),
    .io_enq_valid(io_result_next_b_28_io_enq_valid),
    .io_enq_bits(io_result_next_b_28_io_enq_bits),
    .io_deq_ready(io_result_next_b_28_io_deq_ready),
    .io_deq_valid(io_result_next_b_28_io_deq_valid),
    .io_deq_bits(io_result_next_b_28_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_29 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_29_clock),
    .reset(io_result_next_b_29_reset),
    .io_enq_ready(io_result_next_b_29_io_enq_ready),
    .io_enq_valid(io_result_next_b_29_io_enq_valid),
    .io_enq_bits(io_result_next_b_29_io_enq_bits),
    .io_deq_ready(io_result_next_b_29_io_deq_ready),
    .io_deq_valid(io_result_next_b_29_io_deq_valid),
    .io_deq_bits(io_result_next_b_29_io_deq_bits)
  );
  SkidBuffer_62 io_result_next_b_30 ( // @[MonteCarlo.scala 191:25]
    .clock(io_result_next_b_30_clock),
    .reset(io_result_next_b_30_reset),
    .io_enq_ready(io_result_next_b_30_io_enq_ready),
    .io_enq_valid(io_result_next_b_30_io_enq_valid),
    .io_enq_bits(io_result_next_b_30_io_enq_bits),
    .io_deq_ready(io_result_next_b_30_io_deq_ready),
    .io_deq_valid(io_result_next_b_30_io_deq_valid),
    .io_deq_bits(io_result_next_b_30_io_deq_bits)
  );
  assign io_lanes_0_ready = io_result_next_b_io_enq_ready & _io_result_next_b_io_enq_valid_T; // @[MonteCarlo.scala 194:44]
  assign io_lanes_1_ready = io_result_next_b_io_enq_ready & _io_result_next_b_io_enq_valid_T; // @[MonteCarlo.scala 195:44]
  assign io_lanes_2_ready = io_result_next_b_1_io_enq_ready & _io_result_next_b_io_enq_valid_T_1; // @[MonteCarlo.scala 194:44]
  assign io_lanes_3_ready = io_result_next_b_1_io_enq_ready & _io_result_next_b_io_enq_valid_T_1; // @[MonteCarlo.scala 195:44]
  assign io_lanes_4_ready = io_result_next_b_2_io_enq_ready & _io_result_next_b_io_enq_valid_T_2; // @[MonteCarlo.scala 194:44]
  assign io_lanes_5_ready = io_result_next_b_2_io_enq_ready & _io_result_next_b_io_enq_valid_T_2; // @[MonteCarlo.scala 195:44]
  assign io_lanes_6_ready = io_result_next_b_3_io_enq_ready & _io_result_next_b_io_enq_valid_T_3; // @[MonteCarlo.scala 194:44]
  assign io_lanes_7_ready = io_result_next_b_3_io_enq_ready & _io_result_next_b_io_enq_valid_T_3; // @[MonteCarlo.scala 195:44]
  assign io_lanes_8_ready = io_result_next_b_4_io_enq_ready & _io_result_next_b_io_enq_valid_T_4; // @[MonteCarlo.scala 194:44]
  assign io_lanes_9_ready = io_result_next_b_4_io_enq_ready & _io_result_next_b_io_enq_valid_T_4; // @[MonteCarlo.scala 195:44]
  assign io_lanes_10_ready = io_result_next_b_5_io_enq_ready & _io_result_next_b_io_enq_valid_T_5; // @[MonteCarlo.scala 194:44]
  assign io_lanes_11_ready = io_result_next_b_5_io_enq_ready & _io_result_next_b_io_enq_valid_T_5; // @[MonteCarlo.scala 195:44]
  assign io_lanes_12_ready = io_result_next_b_6_io_enq_ready & _io_result_next_b_io_enq_valid_T_6; // @[MonteCarlo.scala 194:44]
  assign io_lanes_13_ready = io_result_next_b_6_io_enq_ready & _io_result_next_b_io_enq_valid_T_6; // @[MonteCarlo.scala 195:44]
  assign io_lanes_14_ready = io_result_next_b_7_io_enq_ready & _io_result_next_b_io_enq_valid_T_7; // @[MonteCarlo.scala 194:44]
  assign io_lanes_15_ready = io_result_next_b_7_io_enq_ready & _io_result_next_b_io_enq_valid_T_7; // @[MonteCarlo.scala 195:44]
  assign io_lanes_16_ready = io_result_next_b_8_io_enq_ready & _io_result_next_b_io_enq_valid_T_8; // @[MonteCarlo.scala 194:44]
  assign io_lanes_17_ready = io_result_next_b_8_io_enq_ready & _io_result_next_b_io_enq_valid_T_8; // @[MonteCarlo.scala 195:44]
  assign io_lanes_18_ready = io_result_next_b_9_io_enq_ready & _io_result_next_b_io_enq_valid_T_9; // @[MonteCarlo.scala 194:44]
  assign io_lanes_19_ready = io_result_next_b_9_io_enq_ready & _io_result_next_b_io_enq_valid_T_9; // @[MonteCarlo.scala 195:44]
  assign io_lanes_20_ready = io_result_next_b_10_io_enq_ready & _io_result_next_b_io_enq_valid_T_10; // @[MonteCarlo.scala 194:44]
  assign io_lanes_21_ready = io_result_next_b_10_io_enq_ready & _io_result_next_b_io_enq_valid_T_10; // @[MonteCarlo.scala 195:44]
  assign io_lanes_22_ready = io_result_next_b_11_io_enq_ready & _io_result_next_b_io_enq_valid_T_11; // @[MonteCarlo.scala 194:44]
  assign io_lanes_23_ready = io_result_next_b_11_io_enq_ready & _io_result_next_b_io_enq_valid_T_11; // @[MonteCarlo.scala 195:44]
  assign io_lanes_24_ready = io_result_next_b_12_io_enq_ready & _io_result_next_b_io_enq_valid_T_12; // @[MonteCarlo.scala 194:44]
  assign io_lanes_25_ready = io_result_next_b_12_io_enq_ready & _io_result_next_b_io_enq_valid_T_12; // @[MonteCarlo.scala 195:44]
  assign io_lanes_26_ready = io_result_next_b_13_io_enq_ready & _io_result_next_b_io_enq_valid_T_13; // @[MonteCarlo.scala 194:44]
  assign io_lanes_27_ready = io_result_next_b_13_io_enq_ready & _io_result_next_b_io_enq_valid_T_13; // @[MonteCarlo.scala 195:44]
  assign io_lanes_28_ready = io_result_next_b_14_io_enq_ready & _io_result_next_b_io_enq_valid_T_14; // @[MonteCarlo.scala 194:44]
  assign io_lanes_29_ready = io_result_next_b_14_io_enq_ready & _io_result_next_b_io_enq_valid_T_14; // @[MonteCarlo.scala 195:44]
  assign io_lanes_30_ready = io_result_next_b_15_io_enq_ready & _io_result_next_b_io_enq_valid_T_15; // @[MonteCarlo.scala 194:44]
  assign io_lanes_31_ready = io_result_next_b_15_io_enq_ready & _io_result_next_b_io_enq_valid_T_15; // @[MonteCarlo.scala 195:44]
  assign io_result_valid = io_result_next_b_30_io_deq_valid; // @[MonteCarlo.scala 208:13]
  assign io_result_bits = io_result_next_b_30_io_deq_bits; // @[MonteCarlo.scala 208:13]
  assign io_result_next_b_clock = clock;
  assign io_result_next_b_reset = reset;
  assign io_result_next_b_io_enq_valid = io_lanes_0_valid & io_lanes_1_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_io_enq_bits = {{1{io_result_next_r[30]}},io_result_next_r}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_io_deq_ready = io_result_next_b_16_io_enq_ready & _io_result_next_b_io_enq_valid_T_16; // @[MonteCarlo.scala 194:44]
  assign io_result_next_b_1_clock = clock;
  assign io_result_next_b_1_reset = reset;
  assign io_result_next_b_1_io_enq_valid = io_lanes_2_valid & io_lanes_3_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_1_io_enq_bits = {{1{io_result_next_r_1[30]}},io_result_next_r_1}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_1_io_deq_ready = io_result_next_b_16_io_enq_ready & _io_result_next_b_io_enq_valid_T_16; // @[MonteCarlo.scala 195:44]
  assign io_result_next_b_2_clock = clock;
  assign io_result_next_b_2_reset = reset;
  assign io_result_next_b_2_io_enq_valid = io_lanes_4_valid & io_lanes_5_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_2_io_enq_bits = {{1{io_result_next_r_2[30]}},io_result_next_r_2}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_2_io_deq_ready = io_result_next_b_17_io_enq_ready & _io_result_next_b_io_enq_valid_T_17; // @[MonteCarlo.scala 194:44]
  assign io_result_next_b_3_clock = clock;
  assign io_result_next_b_3_reset = reset;
  assign io_result_next_b_3_io_enq_valid = io_lanes_6_valid & io_lanes_7_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_3_io_enq_bits = {{1{io_result_next_r_3[30]}},io_result_next_r_3}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_3_io_deq_ready = io_result_next_b_17_io_enq_ready & _io_result_next_b_io_enq_valid_T_17; // @[MonteCarlo.scala 195:44]
  assign io_result_next_b_4_clock = clock;
  assign io_result_next_b_4_reset = reset;
  assign io_result_next_b_4_io_enq_valid = io_lanes_8_valid & io_lanes_9_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_4_io_enq_bits = {{1{io_result_next_r_4[30]}},io_result_next_r_4}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_4_io_deq_ready = io_result_next_b_18_io_enq_ready & _io_result_next_b_io_enq_valid_T_18; // @[MonteCarlo.scala 194:44]
  assign io_result_next_b_5_clock = clock;
  assign io_result_next_b_5_reset = reset;
  assign io_result_next_b_5_io_enq_valid = io_lanes_10_valid & io_lanes_11_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_5_io_enq_bits = {{1{io_result_next_r_5[30]}},io_result_next_r_5}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_5_io_deq_ready = io_result_next_b_18_io_enq_ready & _io_result_next_b_io_enq_valid_T_18; // @[MonteCarlo.scala 195:44]
  assign io_result_next_b_6_clock = clock;
  assign io_result_next_b_6_reset = reset;
  assign io_result_next_b_6_io_enq_valid = io_lanes_12_valid & io_lanes_13_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_6_io_enq_bits = {{1{io_result_next_r_6[30]}},io_result_next_r_6}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_6_io_deq_ready = io_result_next_b_19_io_enq_ready & _io_result_next_b_io_enq_valid_T_19; // @[MonteCarlo.scala 194:44]
  assign io_result_next_b_7_clock = clock;
  assign io_result_next_b_7_reset = reset;
  assign io_result_next_b_7_io_enq_valid = io_lanes_14_valid & io_lanes_15_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_7_io_enq_bits = {{1{io_result_next_r_7[30]}},io_result_next_r_7}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_7_io_deq_ready = io_result_next_b_19_io_enq_ready & _io_result_next_b_io_enq_valid_T_19; // @[MonteCarlo.scala 195:44]
  assign io_result_next_b_8_clock = clock;
  assign io_result_next_b_8_reset = reset;
  assign io_result_next_b_8_io_enq_valid = io_lanes_16_valid & io_lanes_17_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_8_io_enq_bits = {{1{io_result_next_r_8[30]}},io_result_next_r_8}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_8_io_deq_ready = io_result_next_b_20_io_enq_ready & _io_result_next_b_io_enq_valid_T_20; // @[MonteCarlo.scala 194:44]
  assign io_result_next_b_9_clock = clock;
  assign io_result_next_b_9_reset = reset;
  assign io_result_next_b_9_io_enq_valid = io_lanes_18_valid & io_lanes_19_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_9_io_enq_bits = {{1{io_result_next_r_9[30]}},io_result_next_r_9}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_9_io_deq_ready = io_result_next_b_20_io_enq_ready & _io_result_next_b_io_enq_valid_T_20; // @[MonteCarlo.scala 195:44]
  assign io_result_next_b_10_clock = clock;
  assign io_result_next_b_10_reset = reset;
  assign io_result_next_b_10_io_enq_valid = io_lanes_20_valid & io_lanes_21_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_10_io_enq_bits = {{1{io_result_next_r_10[30]}},io_result_next_r_10}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_10_io_deq_ready = io_result_next_b_21_io_enq_ready & _io_result_next_b_io_enq_valid_T_21; // @[MonteCarlo.scala 194:44]
  assign io_result_next_b_11_clock = clock;
  assign io_result_next_b_11_reset = reset;
  assign io_result_next_b_11_io_enq_valid = io_lanes_22_valid & io_lanes_23_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_11_io_enq_bits = {{1{io_result_next_r_11[30]}},io_result_next_r_11}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_11_io_deq_ready = io_result_next_b_21_io_enq_ready & _io_result_next_b_io_enq_valid_T_21; // @[MonteCarlo.scala 195:44]
  assign io_result_next_b_12_clock = clock;
  assign io_result_next_b_12_reset = reset;
  assign io_result_next_b_12_io_enq_valid = io_lanes_24_valid & io_lanes_25_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_12_io_enq_bits = {{1{io_result_next_r_12[30]}},io_result_next_r_12}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_12_io_deq_ready = io_result_next_b_22_io_enq_ready & _io_result_next_b_io_enq_valid_T_22; // @[MonteCarlo.scala 194:44]
  assign io_result_next_b_13_clock = clock;
  assign io_result_next_b_13_reset = reset;
  assign io_result_next_b_13_io_enq_valid = io_lanes_26_valid & io_lanes_27_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_13_io_enq_bits = {{1{io_result_next_r_13[30]}},io_result_next_r_13}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_13_io_deq_ready = io_result_next_b_22_io_enq_ready & _io_result_next_b_io_enq_valid_T_22; // @[MonteCarlo.scala 195:44]
  assign io_result_next_b_14_clock = clock;
  assign io_result_next_b_14_reset = reset;
  assign io_result_next_b_14_io_enq_valid = io_lanes_28_valid & io_lanes_29_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_14_io_enq_bits = {{1{io_result_next_r_14[30]}},io_result_next_r_14}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_14_io_deq_ready = io_result_next_b_23_io_enq_ready & _io_result_next_b_io_enq_valid_T_23; // @[MonteCarlo.scala 194:44]
  assign io_result_next_b_15_clock = clock;
  assign io_result_next_b_15_reset = reset;
  assign io_result_next_b_15_io_enq_valid = io_lanes_30_valid & io_lanes_31_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_15_io_enq_bits = {{1{io_result_next_r_15[30]}},io_result_next_r_15}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_15_io_deq_ready = io_result_next_b_23_io_enq_ready & _io_result_next_b_io_enq_valid_T_23; // @[MonteCarlo.scala 195:44]
  assign io_result_next_b_16_clock = clock;
  assign io_result_next_b_16_reset = reset;
  assign io_result_next_b_16_io_enq_valid = io_result_next_b_io_deq_valid & io_result_next_b_1_io_deq_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_16_io_enq_bits = {{1{io_result_next_r_16[30]}},io_result_next_r_16}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_16_io_deq_ready = io_result_next_b_24_io_enq_ready & _io_result_next_b_io_enq_valid_T_24; // @[MonteCarlo.scala 194:44]
  assign io_result_next_b_17_clock = clock;
  assign io_result_next_b_17_reset = reset;
  assign io_result_next_b_17_io_enq_valid = io_result_next_b_2_io_deq_valid & io_result_next_b_3_io_deq_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_17_io_enq_bits = {{1{io_result_next_r_17[30]}},io_result_next_r_17}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_17_io_deq_ready = io_result_next_b_24_io_enq_ready & _io_result_next_b_io_enq_valid_T_24; // @[MonteCarlo.scala 195:44]
  assign io_result_next_b_18_clock = clock;
  assign io_result_next_b_18_reset = reset;
  assign io_result_next_b_18_io_enq_valid = io_result_next_b_4_io_deq_valid & io_result_next_b_5_io_deq_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_18_io_enq_bits = {{1{io_result_next_r_18[30]}},io_result_next_r_18}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_18_io_deq_ready = io_result_next_b_25_io_enq_ready & _io_result_next_b_io_enq_valid_T_25; // @[MonteCarlo.scala 194:44]
  assign io_result_next_b_19_clock = clock;
  assign io_result_next_b_19_reset = reset;
  assign io_result_next_b_19_io_enq_valid = io_result_next_b_6_io_deq_valid & io_result_next_b_7_io_deq_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_19_io_enq_bits = {{1{io_result_next_r_19[30]}},io_result_next_r_19}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_19_io_deq_ready = io_result_next_b_25_io_enq_ready & _io_result_next_b_io_enq_valid_T_25; // @[MonteCarlo.scala 195:44]
  assign io_result_next_b_20_clock = clock;
  assign io_result_next_b_20_reset = reset;
  assign io_result_next_b_20_io_enq_valid = io_result_next_b_8_io_deq_valid & io_result_next_b_9_io_deq_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_20_io_enq_bits = {{1{io_result_next_r_20[30]}},io_result_next_r_20}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_20_io_deq_ready = io_result_next_b_26_io_enq_ready & _io_result_next_b_io_enq_valid_T_26; // @[MonteCarlo.scala 194:44]
  assign io_result_next_b_21_clock = clock;
  assign io_result_next_b_21_reset = reset;
  assign io_result_next_b_21_io_enq_valid = io_result_next_b_10_io_deq_valid & io_result_next_b_11_io_deq_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_21_io_enq_bits = {{1{io_result_next_r_21[30]}},io_result_next_r_21}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_21_io_deq_ready = io_result_next_b_26_io_enq_ready & _io_result_next_b_io_enq_valid_T_26; // @[MonteCarlo.scala 195:44]
  assign io_result_next_b_22_clock = clock;
  assign io_result_next_b_22_reset = reset;
  assign io_result_next_b_22_io_enq_valid = io_result_next_b_12_io_deq_valid & io_result_next_b_13_io_deq_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_22_io_enq_bits = {{1{io_result_next_r_22[30]}},io_result_next_r_22}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_22_io_deq_ready = io_result_next_b_27_io_enq_ready & _io_result_next_b_io_enq_valid_T_27; // @[MonteCarlo.scala 194:44]
  assign io_result_next_b_23_clock = clock;
  assign io_result_next_b_23_reset = reset;
  assign io_result_next_b_23_io_enq_valid = io_result_next_b_14_io_deq_valid & io_result_next_b_15_io_deq_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_23_io_enq_bits = {{1{io_result_next_r_23[30]}},io_result_next_r_23}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_23_io_deq_ready = io_result_next_b_27_io_enq_ready & _io_result_next_b_io_enq_valid_T_27; // @[MonteCarlo.scala 195:44]
  assign io_result_next_b_24_clock = clock;
  assign io_result_next_b_24_reset = reset;
  assign io_result_next_b_24_io_enq_valid = io_result_next_b_16_io_deq_valid & io_result_next_b_17_io_deq_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_24_io_enq_bits = {{1{io_result_next_r_24[30]}},io_result_next_r_24}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_24_io_deq_ready = io_result_next_b_28_io_enq_ready & _io_result_next_b_io_enq_valid_T_28; // @[MonteCarlo.scala 194:44]
  assign io_result_next_b_25_clock = clock;
  assign io_result_next_b_25_reset = reset;
  assign io_result_next_b_25_io_enq_valid = io_result_next_b_18_io_deq_valid & io_result_next_b_19_io_deq_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_25_io_enq_bits = {{1{io_result_next_r_25[30]}},io_result_next_r_25}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_25_io_deq_ready = io_result_next_b_28_io_enq_ready & _io_result_next_b_io_enq_valid_T_28; // @[MonteCarlo.scala 195:44]
  assign io_result_next_b_26_clock = clock;
  assign io_result_next_b_26_reset = reset;
  assign io_result_next_b_26_io_enq_valid = io_result_next_b_20_io_deq_valid & io_result_next_b_21_io_deq_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_26_io_enq_bits = {{1{io_result_next_r_26[30]}},io_result_next_r_26}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_26_io_deq_ready = io_result_next_b_29_io_enq_ready & _io_result_next_b_io_enq_valid_T_29; // @[MonteCarlo.scala 194:44]
  assign io_result_next_b_27_clock = clock;
  assign io_result_next_b_27_reset = reset;
  assign io_result_next_b_27_io_enq_valid = io_result_next_b_22_io_deq_valid & io_result_next_b_23_io_deq_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_27_io_enq_bits = {{1{io_result_next_r_27[30]}},io_result_next_r_27}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_27_io_deq_ready = io_result_next_b_29_io_enq_ready & _io_result_next_b_io_enq_valid_T_29; // @[MonteCarlo.scala 195:44]
  assign io_result_next_b_28_clock = clock;
  assign io_result_next_b_28_reset = reset;
  assign io_result_next_b_28_io_enq_valid = io_result_next_b_24_io_deq_valid & io_result_next_b_25_io_deq_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_28_io_enq_bits = {{1{io_result_next_r_28[30]}},io_result_next_r_28}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_28_io_deq_ready = io_result_next_b_30_io_enq_ready & _io_result_next_b_io_enq_valid_T_30; // @[MonteCarlo.scala 194:44]
  assign io_result_next_b_29_clock = clock;
  assign io_result_next_b_29_reset = reset;
  assign io_result_next_b_29_io_enq_valid = io_result_next_b_26_io_deq_valid & io_result_next_b_27_io_deq_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_29_io_enq_bits = {{1{io_result_next_r_29[30]}},io_result_next_r_29}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_29_io_deq_ready = io_result_next_b_30_io_enq_ready & _io_result_next_b_io_enq_valid_T_30; // @[MonteCarlo.scala 195:44]
  assign io_result_next_b_30_clock = clock;
  assign io_result_next_b_30_reset = reset;
  assign io_result_next_b_30_io_enq_valid = io_result_next_b_28_io_deq_valid & io_result_next_b_29_io_deq_valid; // @[MonteCarlo.scala 193:42]
  assign io_result_next_b_30_io_enq_bits = {{1{io_result_next_r_30[30]}},io_result_next_r_30}; // @[MonteCarlo.scala 192:26]
  assign io_result_next_b_30_io_deq_ready = io_result_ready; // @[MonteCarlo.scala 208:13]
endmodule
module MonteCarloAccelerator(
  input         clock,
  input         reset,
  output        io_request_ready,
  input         io_request_valid,
  input  [31:0] io_request_bits_time_steps,
  input  [31:0] io_request_bits_start_value,
  input  [31:0] io_request_bits_coefficient1,
  input  [31:0] io_request_bits_coefficient2,
  input         io_response_ready,
  output        io_response_valid,
  output [31:0] io_response_bits
);
  wire  engines_0_clock; // @[MonteCarlo.scala 254:48]
  wire  engines_0_reset; // @[MonteCarlo.scala 254:48]
  wire  engines_0_io_request_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_0_io_request_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_0_io_request_0_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_0_io_request_0_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_0_io_request_0_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_0_io_request_0_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_0_io_request_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_0_io_request_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_0_io_request_1_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_0_io_request_1_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_0_io_request_1_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_0_io_request_1_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_0_io_response_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_0_io_response_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_0_io_response_0_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_0_io_response_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_0_io_response_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_0_io_response_1_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_1_clock; // @[MonteCarlo.scala 254:48]
  wire  engines_1_reset; // @[MonteCarlo.scala 254:48]
  wire  engines_1_io_request_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_1_io_request_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_1_io_request_0_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_1_io_request_0_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_1_io_request_0_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_1_io_request_0_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_1_io_request_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_1_io_request_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_1_io_request_1_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_1_io_request_1_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_1_io_request_1_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_1_io_request_1_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_1_io_response_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_1_io_response_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_1_io_response_0_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_1_io_response_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_1_io_response_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_1_io_response_1_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_2_clock; // @[MonteCarlo.scala 254:48]
  wire  engines_2_reset; // @[MonteCarlo.scala 254:48]
  wire  engines_2_io_request_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_2_io_request_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_2_io_request_0_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_2_io_request_0_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_2_io_request_0_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_2_io_request_0_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_2_io_request_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_2_io_request_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_2_io_request_1_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_2_io_request_1_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_2_io_request_1_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_2_io_request_1_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_2_io_response_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_2_io_response_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_2_io_response_0_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_2_io_response_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_2_io_response_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_2_io_response_1_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_3_clock; // @[MonteCarlo.scala 254:48]
  wire  engines_3_reset; // @[MonteCarlo.scala 254:48]
  wire  engines_3_io_request_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_3_io_request_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_3_io_request_0_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_3_io_request_0_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_3_io_request_0_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_3_io_request_0_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_3_io_request_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_3_io_request_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_3_io_request_1_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_3_io_request_1_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_3_io_request_1_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_3_io_request_1_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_3_io_response_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_3_io_response_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_3_io_response_0_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_3_io_response_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_3_io_response_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_3_io_response_1_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_4_clock; // @[MonteCarlo.scala 254:48]
  wire  engines_4_reset; // @[MonteCarlo.scala 254:48]
  wire  engines_4_io_request_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_4_io_request_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_4_io_request_0_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_4_io_request_0_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_4_io_request_0_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_4_io_request_0_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_4_io_request_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_4_io_request_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_4_io_request_1_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_4_io_request_1_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_4_io_request_1_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_4_io_request_1_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_4_io_response_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_4_io_response_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_4_io_response_0_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_4_io_response_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_4_io_response_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_4_io_response_1_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_5_clock; // @[MonteCarlo.scala 254:48]
  wire  engines_5_reset; // @[MonteCarlo.scala 254:48]
  wire  engines_5_io_request_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_5_io_request_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_5_io_request_0_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_5_io_request_0_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_5_io_request_0_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_5_io_request_0_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_5_io_request_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_5_io_request_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_5_io_request_1_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_5_io_request_1_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_5_io_request_1_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_5_io_request_1_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_5_io_response_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_5_io_response_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_5_io_response_0_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_5_io_response_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_5_io_response_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_5_io_response_1_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_6_clock; // @[MonteCarlo.scala 254:48]
  wire  engines_6_reset; // @[MonteCarlo.scala 254:48]
  wire  engines_6_io_request_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_6_io_request_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_6_io_request_0_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_6_io_request_0_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_6_io_request_0_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_6_io_request_0_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_6_io_request_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_6_io_request_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_6_io_request_1_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_6_io_request_1_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_6_io_request_1_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_6_io_request_1_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_6_io_response_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_6_io_response_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_6_io_response_0_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_6_io_response_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_6_io_response_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_6_io_response_1_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_7_clock; // @[MonteCarlo.scala 254:48]
  wire  engines_7_reset; // @[MonteCarlo.scala 254:48]
  wire  engines_7_io_request_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_7_io_request_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_7_io_request_0_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_7_io_request_0_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_7_io_request_0_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_7_io_request_0_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_7_io_request_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_7_io_request_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_7_io_request_1_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_7_io_request_1_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_7_io_request_1_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_7_io_request_1_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_7_io_response_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_7_io_response_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_7_io_response_0_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_7_io_response_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_7_io_response_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_7_io_response_1_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_8_clock; // @[MonteCarlo.scala 254:48]
  wire  engines_8_reset; // @[MonteCarlo.scala 254:48]
  wire  engines_8_io_request_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_8_io_request_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_8_io_request_0_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_8_io_request_0_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_8_io_request_0_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_8_io_request_0_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_8_io_request_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_8_io_request_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_8_io_request_1_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_8_io_request_1_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_8_io_request_1_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_8_io_request_1_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_8_io_response_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_8_io_response_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_8_io_response_0_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_8_io_response_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_8_io_response_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_8_io_response_1_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_9_clock; // @[MonteCarlo.scala 254:48]
  wire  engines_9_reset; // @[MonteCarlo.scala 254:48]
  wire  engines_9_io_request_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_9_io_request_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_9_io_request_0_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_9_io_request_0_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_9_io_request_0_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_9_io_request_0_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_9_io_request_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_9_io_request_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_9_io_request_1_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_9_io_request_1_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_9_io_request_1_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_9_io_request_1_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_9_io_response_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_9_io_response_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_9_io_response_0_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_9_io_response_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_9_io_response_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_9_io_response_1_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_10_clock; // @[MonteCarlo.scala 254:48]
  wire  engines_10_reset; // @[MonteCarlo.scala 254:48]
  wire  engines_10_io_request_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_10_io_request_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_10_io_request_0_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_10_io_request_0_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_10_io_request_0_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_10_io_request_0_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_10_io_request_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_10_io_request_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_10_io_request_1_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_10_io_request_1_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_10_io_request_1_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_10_io_request_1_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_10_io_response_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_10_io_response_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_10_io_response_0_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_10_io_response_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_10_io_response_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_10_io_response_1_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_11_clock; // @[MonteCarlo.scala 254:48]
  wire  engines_11_reset; // @[MonteCarlo.scala 254:48]
  wire  engines_11_io_request_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_11_io_request_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_11_io_request_0_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_11_io_request_0_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_11_io_request_0_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_11_io_request_0_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_11_io_request_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_11_io_request_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_11_io_request_1_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_11_io_request_1_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_11_io_request_1_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_11_io_request_1_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_11_io_response_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_11_io_response_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_11_io_response_0_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_11_io_response_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_11_io_response_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_11_io_response_1_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_12_clock; // @[MonteCarlo.scala 254:48]
  wire  engines_12_reset; // @[MonteCarlo.scala 254:48]
  wire  engines_12_io_request_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_12_io_request_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_12_io_request_0_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_12_io_request_0_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_12_io_request_0_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_12_io_request_0_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_12_io_request_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_12_io_request_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_12_io_request_1_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_12_io_request_1_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_12_io_request_1_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_12_io_request_1_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_12_io_response_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_12_io_response_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_12_io_response_0_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_12_io_response_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_12_io_response_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_12_io_response_1_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_13_clock; // @[MonteCarlo.scala 254:48]
  wire  engines_13_reset; // @[MonteCarlo.scala 254:48]
  wire  engines_13_io_request_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_13_io_request_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_13_io_request_0_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_13_io_request_0_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_13_io_request_0_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_13_io_request_0_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_13_io_request_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_13_io_request_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_13_io_request_1_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_13_io_request_1_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_13_io_request_1_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_13_io_request_1_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_13_io_response_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_13_io_response_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_13_io_response_0_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_13_io_response_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_13_io_response_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_13_io_response_1_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_14_clock; // @[MonteCarlo.scala 254:48]
  wire  engines_14_reset; // @[MonteCarlo.scala 254:48]
  wire  engines_14_io_request_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_14_io_request_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_14_io_request_0_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_14_io_request_0_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_14_io_request_0_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_14_io_request_0_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_14_io_request_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_14_io_request_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_14_io_request_1_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_14_io_request_1_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_14_io_request_1_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_14_io_request_1_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_14_io_response_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_14_io_response_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_14_io_response_0_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_14_io_response_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_14_io_response_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_14_io_response_1_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_15_clock; // @[MonteCarlo.scala 254:48]
  wire  engines_15_reset; // @[MonteCarlo.scala 254:48]
  wire  engines_15_io_request_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_15_io_request_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_15_io_request_0_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_15_io_request_0_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_15_io_request_0_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_15_io_request_0_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_15_io_request_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_15_io_request_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_15_io_request_1_bits_time_steps; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_15_io_request_1_bits_start_value; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_15_io_request_1_bits_coefficient1; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_15_io_request_1_bits_coefficient2; // @[MonteCarlo.scala 254:48]
  wire  engines_15_io_response_0_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_15_io_response_0_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_15_io_response_0_bits; // @[MonteCarlo.scala 254:48]
  wire  engines_15_io_response_1_ready; // @[MonteCarlo.scala 254:48]
  wire  engines_15_io_response_1_valid; // @[MonteCarlo.scala 254:48]
  wire [31:0] engines_15_io_response_1_bits; // @[MonteCarlo.scala 254:48]
  wire  b1_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_1_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_1_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_1_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_1_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_1_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_1_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_1_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_1_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_1_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_1_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_1_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_1_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_1_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_1_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_1_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_1_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_1_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_1_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_1_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_1_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_1_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_1_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_1_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_1_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_1_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_1_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_1_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_1_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_2_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_2_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_2_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_2_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_2_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_2_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_2_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_2_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_2_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_2_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_2_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_2_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_2_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_2_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_2_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_2_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_2_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_2_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_2_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_2_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_2_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_2_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_2_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_2_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_2_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_2_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_2_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_2_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_3_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_3_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_3_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_3_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_3_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_3_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_3_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_3_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_3_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_3_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_3_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_3_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_3_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_3_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_3_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_3_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_3_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_3_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_3_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_3_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_3_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_3_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_3_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_3_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_3_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_3_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_3_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_3_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_4_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_4_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_4_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_4_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_4_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_4_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_4_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_4_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_4_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_4_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_4_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_4_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_4_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_4_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_4_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_4_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_4_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_4_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_4_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_4_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_4_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_4_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_4_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_4_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_4_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_4_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_4_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_4_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_5_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_5_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_5_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_5_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_5_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_5_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_5_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_5_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_5_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_5_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_5_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_5_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_5_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_5_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_5_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_5_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_5_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_5_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_5_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_5_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_5_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_5_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_5_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_5_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_5_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_5_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_5_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_5_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_6_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_6_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_6_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_6_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_6_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_6_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_6_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_6_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_6_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_6_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_6_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_6_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_6_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_6_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_6_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_6_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_6_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_6_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_6_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_6_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_6_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_6_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_6_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_6_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_6_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_6_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_6_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_6_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_7_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_7_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_7_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_7_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_7_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_7_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_7_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_7_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_7_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_7_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_7_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_7_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_7_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_7_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_7_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_7_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_7_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_7_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_7_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_7_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_7_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_7_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_7_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_7_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_7_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_7_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_7_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_7_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_8_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_8_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_8_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_8_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_8_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_8_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_8_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_8_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_8_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_8_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_8_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_8_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_8_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_8_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_8_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_8_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_8_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_8_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_8_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_8_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_8_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_8_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_8_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_8_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_8_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_8_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_8_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_8_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_9_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_9_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_9_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_9_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_9_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_9_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_9_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_9_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_9_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_9_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_9_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_9_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_9_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_9_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_9_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_9_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_9_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_9_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_9_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_9_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_9_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_9_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_9_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_9_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_9_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_9_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_9_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_9_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_10_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_10_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_10_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_10_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_10_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_10_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_10_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_10_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_10_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_10_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_10_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_10_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_10_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_10_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_10_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_10_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_10_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_10_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_10_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_10_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_10_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_10_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_10_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_10_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_10_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_10_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_10_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_10_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_11_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_11_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_11_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_11_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_11_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_11_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_11_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_11_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_11_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_11_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_11_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_11_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_11_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_11_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_11_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_11_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_11_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_11_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_11_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_11_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_11_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_11_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_11_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_11_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_11_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_11_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_11_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_11_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_12_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_12_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_12_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_12_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_12_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_12_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_12_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_12_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_12_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_12_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_12_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_12_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_12_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_12_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_12_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_12_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_12_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_12_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_12_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_12_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_12_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_12_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_12_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_12_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_12_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_12_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_12_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_12_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_13_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_13_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_13_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_13_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_13_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_13_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_13_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_13_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_13_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_13_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_13_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_13_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_13_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_13_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_13_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_13_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_13_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_13_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_13_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_13_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_13_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_13_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_13_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_13_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_13_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_13_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_13_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_13_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_14_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_14_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_14_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_14_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_14_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_14_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_14_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_14_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_14_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_14_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_14_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_14_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_14_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_14_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_14_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_14_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_14_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_14_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_14_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_14_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_14_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_14_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_14_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_14_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_14_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_14_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_14_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_14_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_15_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_15_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_15_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_15_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_15_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_15_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_15_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_15_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_15_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_15_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_15_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_15_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_15_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_15_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_15_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_15_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_15_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_15_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_15_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_15_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_15_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_15_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_15_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_15_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_15_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_15_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_15_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_15_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_16_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_16_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_16_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_16_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_16_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_16_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_16_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_16_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_16_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_16_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_16_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_16_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_16_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_16_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_16_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_16_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_16_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_16_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_16_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_16_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_16_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_16_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_16_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_16_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_16_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_16_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_16_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_16_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_17_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_17_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_17_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_17_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_17_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_17_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_17_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_17_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_17_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_17_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_17_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_17_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_17_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_17_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_17_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_17_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_17_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_17_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_17_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_17_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_17_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_17_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_17_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_17_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_17_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_17_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_17_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_17_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_18_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_18_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_18_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_18_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_18_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_18_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_18_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_18_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_18_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_18_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_18_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_18_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_18_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_18_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_18_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_18_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_18_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_18_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_18_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_18_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_18_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_18_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_18_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_18_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_18_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_18_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_18_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_18_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_19_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_19_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_19_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_19_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_19_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_19_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_19_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_19_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_19_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_19_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_19_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_19_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_19_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_19_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_19_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_19_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_19_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_19_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_19_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_19_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_19_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_19_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_19_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_19_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_19_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_19_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_19_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_19_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_20_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_20_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_20_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_20_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_20_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_20_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_20_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_20_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_20_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_20_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_20_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_20_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_20_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_20_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_20_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_20_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_20_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_20_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_20_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_20_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_20_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_20_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_20_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_20_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_20_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_20_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_20_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_20_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_21_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_21_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_21_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_21_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_21_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_21_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_21_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_21_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_21_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_21_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_21_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_21_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_21_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_21_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_21_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_21_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_21_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_21_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_21_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_21_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_21_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_21_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_21_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_21_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_21_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_21_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_21_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_21_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_22_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_22_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_22_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_22_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_22_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_22_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_22_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_22_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_22_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_22_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_22_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_22_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_22_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_22_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_22_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_22_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_22_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_22_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_22_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_22_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_22_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_22_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_22_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_22_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_22_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_22_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_22_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_22_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_23_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_23_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_23_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_23_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_23_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_23_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_23_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_23_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_23_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_23_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_23_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_23_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_23_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_23_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_23_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_23_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_23_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_23_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_23_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_23_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_23_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_23_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_23_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_23_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_23_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_23_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_23_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_23_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_24_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_24_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_24_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_24_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_24_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_24_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_24_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_24_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_24_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_24_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_24_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_24_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_24_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_24_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_24_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_24_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_24_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_24_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_24_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_24_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_24_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_24_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_24_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_24_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_24_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_24_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_24_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_24_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_25_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_25_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_25_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_25_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_25_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_25_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_25_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_25_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_25_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_25_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_25_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_25_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_25_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_25_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_25_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_25_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_25_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_25_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_25_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_25_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_25_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_25_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_25_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_25_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_25_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_25_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_25_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_25_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_26_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_26_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_26_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_26_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_26_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_26_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_26_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_26_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_26_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_26_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_26_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_26_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_26_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_26_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_26_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_26_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_26_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_26_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_26_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_26_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_26_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_26_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_26_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_26_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_26_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_26_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_26_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_26_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_27_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_27_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_27_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_27_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_27_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_27_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_27_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_27_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_27_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_27_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_27_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_27_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_27_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_27_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_27_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_27_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_27_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_27_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_27_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_27_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_27_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_27_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_27_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_27_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_27_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_27_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_27_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_27_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_28_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_28_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_28_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_28_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_28_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_28_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_28_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_28_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_28_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_28_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_28_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_28_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_28_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_28_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_28_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_28_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_28_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_28_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_28_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_28_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_28_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_28_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_28_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_28_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_28_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_28_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_28_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_28_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_29_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_29_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_29_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_29_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_29_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_29_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_29_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_29_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_29_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_29_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_29_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_29_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_29_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_29_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_29_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_29_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_29_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_29_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_29_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_29_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_29_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_29_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_29_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_29_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_29_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_29_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_29_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_29_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b1_30_clock; // @[MonteCarlo.scala 239:27]
  wire  b1_30_reset; // @[MonteCarlo.scala 239:27]
  wire  b1_30_io_enq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_30_io_enq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_30_io_enq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_30_io_enq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_30_io_enq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_30_io_enq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b1_30_io_deq_ready; // @[MonteCarlo.scala 239:27]
  wire  b1_30_io_deq_valid; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_30_io_deq_bits_time_steps; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_30_io_deq_bits_start_value; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_30_io_deq_bits_coefficient1; // @[MonteCarlo.scala 239:27]
  wire [31:0] b1_30_io_deq_bits_coefficient2; // @[MonteCarlo.scala 239:27]
  wire  b2_30_clock; // @[MonteCarlo.scala 240:27]
  wire  b2_30_reset; // @[MonteCarlo.scala 240:27]
  wire  b2_30_io_enq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_30_io_enq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_30_io_enq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_30_io_enq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_30_io_enq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_30_io_enq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  b2_30_io_deq_ready; // @[MonteCarlo.scala 240:27]
  wire  b2_30_io_deq_valid; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_30_io_deq_bits_time_steps; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_30_io_deq_bits_start_value; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_30_io_deq_bits_coefficient1; // @[MonteCarlo.scala 240:27]
  wire [31:0] b2_30_io_deq_bits_coefficient2; // @[MonteCarlo.scala 240:27]
  wire  partial_result_impl_clock; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_reset; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_0_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_0_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_0_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_1_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_1_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_1_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_2_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_2_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_2_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_3_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_3_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_3_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_4_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_4_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_4_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_5_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_5_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_5_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_6_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_6_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_6_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_7_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_7_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_7_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_8_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_8_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_8_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_9_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_9_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_9_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_10_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_10_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_10_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_11_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_11_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_11_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_12_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_12_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_12_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_13_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_13_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_13_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_14_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_14_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_14_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_15_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_15_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_15_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_16_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_16_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_16_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_17_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_17_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_17_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_18_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_18_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_18_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_19_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_19_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_19_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_20_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_20_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_20_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_21_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_21_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_21_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_22_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_22_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_22_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_23_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_23_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_23_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_24_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_24_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_24_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_25_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_25_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_25_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_26_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_26_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_26_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_27_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_27_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_27_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_28_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_28_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_28_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_29_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_29_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_29_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_30_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_30_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_30_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_31_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_lanes_31_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_lanes_31_bits; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_result_ready; // @[MonteCarlo.scala 215:22]
  wire  partial_result_impl_io_result_valid; // @[MonteCarlo.scala 215:22]
  wire [31:0] partial_result_impl_io_result_bits; // @[MonteCarlo.scala 215:22]
  MonteCarlo engines_0 ( // @[MonteCarlo.scala 254:48]
    .clock(engines_0_clock),
    .reset(engines_0_reset),
    .io_request_0_ready(engines_0_io_request_0_ready),
    .io_request_0_valid(engines_0_io_request_0_valid),
    .io_request_0_bits_time_steps(engines_0_io_request_0_bits_time_steps),
    .io_request_0_bits_start_value(engines_0_io_request_0_bits_start_value),
    .io_request_0_bits_coefficient1(engines_0_io_request_0_bits_coefficient1),
    .io_request_0_bits_coefficient2(engines_0_io_request_0_bits_coefficient2),
    .io_request_1_ready(engines_0_io_request_1_ready),
    .io_request_1_valid(engines_0_io_request_1_valid),
    .io_request_1_bits_time_steps(engines_0_io_request_1_bits_time_steps),
    .io_request_1_bits_start_value(engines_0_io_request_1_bits_start_value),
    .io_request_1_bits_coefficient1(engines_0_io_request_1_bits_coefficient1),
    .io_request_1_bits_coefficient2(engines_0_io_request_1_bits_coefficient2),
    .io_response_0_ready(engines_0_io_response_0_ready),
    .io_response_0_valid(engines_0_io_response_0_valid),
    .io_response_0_bits(engines_0_io_response_0_bits),
    .io_response_1_ready(engines_0_io_response_1_ready),
    .io_response_1_valid(engines_0_io_response_1_valid),
    .io_response_1_bits(engines_0_io_response_1_bits)
  );
  MonteCarlo_1 engines_1 ( // @[MonteCarlo.scala 254:48]
    .clock(engines_1_clock),
    .reset(engines_1_reset),
    .io_request_0_ready(engines_1_io_request_0_ready),
    .io_request_0_valid(engines_1_io_request_0_valid),
    .io_request_0_bits_time_steps(engines_1_io_request_0_bits_time_steps),
    .io_request_0_bits_start_value(engines_1_io_request_0_bits_start_value),
    .io_request_0_bits_coefficient1(engines_1_io_request_0_bits_coefficient1),
    .io_request_0_bits_coefficient2(engines_1_io_request_0_bits_coefficient2),
    .io_request_1_ready(engines_1_io_request_1_ready),
    .io_request_1_valid(engines_1_io_request_1_valid),
    .io_request_1_bits_time_steps(engines_1_io_request_1_bits_time_steps),
    .io_request_1_bits_start_value(engines_1_io_request_1_bits_start_value),
    .io_request_1_bits_coefficient1(engines_1_io_request_1_bits_coefficient1),
    .io_request_1_bits_coefficient2(engines_1_io_request_1_bits_coefficient2),
    .io_response_0_ready(engines_1_io_response_0_ready),
    .io_response_0_valid(engines_1_io_response_0_valid),
    .io_response_0_bits(engines_1_io_response_0_bits),
    .io_response_1_ready(engines_1_io_response_1_ready),
    .io_response_1_valid(engines_1_io_response_1_valid),
    .io_response_1_bits(engines_1_io_response_1_bits)
  );
  MonteCarlo_2 engines_2 ( // @[MonteCarlo.scala 254:48]
    .clock(engines_2_clock),
    .reset(engines_2_reset),
    .io_request_0_ready(engines_2_io_request_0_ready),
    .io_request_0_valid(engines_2_io_request_0_valid),
    .io_request_0_bits_time_steps(engines_2_io_request_0_bits_time_steps),
    .io_request_0_bits_start_value(engines_2_io_request_0_bits_start_value),
    .io_request_0_bits_coefficient1(engines_2_io_request_0_bits_coefficient1),
    .io_request_0_bits_coefficient2(engines_2_io_request_0_bits_coefficient2),
    .io_request_1_ready(engines_2_io_request_1_ready),
    .io_request_1_valid(engines_2_io_request_1_valid),
    .io_request_1_bits_time_steps(engines_2_io_request_1_bits_time_steps),
    .io_request_1_bits_start_value(engines_2_io_request_1_bits_start_value),
    .io_request_1_bits_coefficient1(engines_2_io_request_1_bits_coefficient1),
    .io_request_1_bits_coefficient2(engines_2_io_request_1_bits_coefficient2),
    .io_response_0_ready(engines_2_io_response_0_ready),
    .io_response_0_valid(engines_2_io_response_0_valid),
    .io_response_0_bits(engines_2_io_response_0_bits),
    .io_response_1_ready(engines_2_io_response_1_ready),
    .io_response_1_valid(engines_2_io_response_1_valid),
    .io_response_1_bits(engines_2_io_response_1_bits)
  );
  MonteCarlo_3 engines_3 ( // @[MonteCarlo.scala 254:48]
    .clock(engines_3_clock),
    .reset(engines_3_reset),
    .io_request_0_ready(engines_3_io_request_0_ready),
    .io_request_0_valid(engines_3_io_request_0_valid),
    .io_request_0_bits_time_steps(engines_3_io_request_0_bits_time_steps),
    .io_request_0_bits_start_value(engines_3_io_request_0_bits_start_value),
    .io_request_0_bits_coefficient1(engines_3_io_request_0_bits_coefficient1),
    .io_request_0_bits_coefficient2(engines_3_io_request_0_bits_coefficient2),
    .io_request_1_ready(engines_3_io_request_1_ready),
    .io_request_1_valid(engines_3_io_request_1_valid),
    .io_request_1_bits_time_steps(engines_3_io_request_1_bits_time_steps),
    .io_request_1_bits_start_value(engines_3_io_request_1_bits_start_value),
    .io_request_1_bits_coefficient1(engines_3_io_request_1_bits_coefficient1),
    .io_request_1_bits_coefficient2(engines_3_io_request_1_bits_coefficient2),
    .io_response_0_ready(engines_3_io_response_0_ready),
    .io_response_0_valid(engines_3_io_response_0_valid),
    .io_response_0_bits(engines_3_io_response_0_bits),
    .io_response_1_ready(engines_3_io_response_1_ready),
    .io_response_1_valid(engines_3_io_response_1_valid),
    .io_response_1_bits(engines_3_io_response_1_bits)
  );
  MonteCarlo_4 engines_4 ( // @[MonteCarlo.scala 254:48]
    .clock(engines_4_clock),
    .reset(engines_4_reset),
    .io_request_0_ready(engines_4_io_request_0_ready),
    .io_request_0_valid(engines_4_io_request_0_valid),
    .io_request_0_bits_time_steps(engines_4_io_request_0_bits_time_steps),
    .io_request_0_bits_start_value(engines_4_io_request_0_bits_start_value),
    .io_request_0_bits_coefficient1(engines_4_io_request_0_bits_coefficient1),
    .io_request_0_bits_coefficient2(engines_4_io_request_0_bits_coefficient2),
    .io_request_1_ready(engines_4_io_request_1_ready),
    .io_request_1_valid(engines_4_io_request_1_valid),
    .io_request_1_bits_time_steps(engines_4_io_request_1_bits_time_steps),
    .io_request_1_bits_start_value(engines_4_io_request_1_bits_start_value),
    .io_request_1_bits_coefficient1(engines_4_io_request_1_bits_coefficient1),
    .io_request_1_bits_coefficient2(engines_4_io_request_1_bits_coefficient2),
    .io_response_0_ready(engines_4_io_response_0_ready),
    .io_response_0_valid(engines_4_io_response_0_valid),
    .io_response_0_bits(engines_4_io_response_0_bits),
    .io_response_1_ready(engines_4_io_response_1_ready),
    .io_response_1_valid(engines_4_io_response_1_valid),
    .io_response_1_bits(engines_4_io_response_1_bits)
  );
  MonteCarlo_5 engines_5 ( // @[MonteCarlo.scala 254:48]
    .clock(engines_5_clock),
    .reset(engines_5_reset),
    .io_request_0_ready(engines_5_io_request_0_ready),
    .io_request_0_valid(engines_5_io_request_0_valid),
    .io_request_0_bits_time_steps(engines_5_io_request_0_bits_time_steps),
    .io_request_0_bits_start_value(engines_5_io_request_0_bits_start_value),
    .io_request_0_bits_coefficient1(engines_5_io_request_0_bits_coefficient1),
    .io_request_0_bits_coefficient2(engines_5_io_request_0_bits_coefficient2),
    .io_request_1_ready(engines_5_io_request_1_ready),
    .io_request_1_valid(engines_5_io_request_1_valid),
    .io_request_1_bits_time_steps(engines_5_io_request_1_bits_time_steps),
    .io_request_1_bits_start_value(engines_5_io_request_1_bits_start_value),
    .io_request_1_bits_coefficient1(engines_5_io_request_1_bits_coefficient1),
    .io_request_1_bits_coefficient2(engines_5_io_request_1_bits_coefficient2),
    .io_response_0_ready(engines_5_io_response_0_ready),
    .io_response_0_valid(engines_5_io_response_0_valid),
    .io_response_0_bits(engines_5_io_response_0_bits),
    .io_response_1_ready(engines_5_io_response_1_ready),
    .io_response_1_valid(engines_5_io_response_1_valid),
    .io_response_1_bits(engines_5_io_response_1_bits)
  );
  MonteCarlo_6 engines_6 ( // @[MonteCarlo.scala 254:48]
    .clock(engines_6_clock),
    .reset(engines_6_reset),
    .io_request_0_ready(engines_6_io_request_0_ready),
    .io_request_0_valid(engines_6_io_request_0_valid),
    .io_request_0_bits_time_steps(engines_6_io_request_0_bits_time_steps),
    .io_request_0_bits_start_value(engines_6_io_request_0_bits_start_value),
    .io_request_0_bits_coefficient1(engines_6_io_request_0_bits_coefficient1),
    .io_request_0_bits_coefficient2(engines_6_io_request_0_bits_coefficient2),
    .io_request_1_ready(engines_6_io_request_1_ready),
    .io_request_1_valid(engines_6_io_request_1_valid),
    .io_request_1_bits_time_steps(engines_6_io_request_1_bits_time_steps),
    .io_request_1_bits_start_value(engines_6_io_request_1_bits_start_value),
    .io_request_1_bits_coefficient1(engines_6_io_request_1_bits_coefficient1),
    .io_request_1_bits_coefficient2(engines_6_io_request_1_bits_coefficient2),
    .io_response_0_ready(engines_6_io_response_0_ready),
    .io_response_0_valid(engines_6_io_response_0_valid),
    .io_response_0_bits(engines_6_io_response_0_bits),
    .io_response_1_ready(engines_6_io_response_1_ready),
    .io_response_1_valid(engines_6_io_response_1_valid),
    .io_response_1_bits(engines_6_io_response_1_bits)
  );
  MonteCarlo_7 engines_7 ( // @[MonteCarlo.scala 254:48]
    .clock(engines_7_clock),
    .reset(engines_7_reset),
    .io_request_0_ready(engines_7_io_request_0_ready),
    .io_request_0_valid(engines_7_io_request_0_valid),
    .io_request_0_bits_time_steps(engines_7_io_request_0_bits_time_steps),
    .io_request_0_bits_start_value(engines_7_io_request_0_bits_start_value),
    .io_request_0_bits_coefficient1(engines_7_io_request_0_bits_coefficient1),
    .io_request_0_bits_coefficient2(engines_7_io_request_0_bits_coefficient2),
    .io_request_1_ready(engines_7_io_request_1_ready),
    .io_request_1_valid(engines_7_io_request_1_valid),
    .io_request_1_bits_time_steps(engines_7_io_request_1_bits_time_steps),
    .io_request_1_bits_start_value(engines_7_io_request_1_bits_start_value),
    .io_request_1_bits_coefficient1(engines_7_io_request_1_bits_coefficient1),
    .io_request_1_bits_coefficient2(engines_7_io_request_1_bits_coefficient2),
    .io_response_0_ready(engines_7_io_response_0_ready),
    .io_response_0_valid(engines_7_io_response_0_valid),
    .io_response_0_bits(engines_7_io_response_0_bits),
    .io_response_1_ready(engines_7_io_response_1_ready),
    .io_response_1_valid(engines_7_io_response_1_valid),
    .io_response_1_bits(engines_7_io_response_1_bits)
  );
  MonteCarlo_8 engines_8 ( // @[MonteCarlo.scala 254:48]
    .clock(engines_8_clock),
    .reset(engines_8_reset),
    .io_request_0_ready(engines_8_io_request_0_ready),
    .io_request_0_valid(engines_8_io_request_0_valid),
    .io_request_0_bits_time_steps(engines_8_io_request_0_bits_time_steps),
    .io_request_0_bits_start_value(engines_8_io_request_0_bits_start_value),
    .io_request_0_bits_coefficient1(engines_8_io_request_0_bits_coefficient1),
    .io_request_0_bits_coefficient2(engines_8_io_request_0_bits_coefficient2),
    .io_request_1_ready(engines_8_io_request_1_ready),
    .io_request_1_valid(engines_8_io_request_1_valid),
    .io_request_1_bits_time_steps(engines_8_io_request_1_bits_time_steps),
    .io_request_1_bits_start_value(engines_8_io_request_1_bits_start_value),
    .io_request_1_bits_coefficient1(engines_8_io_request_1_bits_coefficient1),
    .io_request_1_bits_coefficient2(engines_8_io_request_1_bits_coefficient2),
    .io_response_0_ready(engines_8_io_response_0_ready),
    .io_response_0_valid(engines_8_io_response_0_valid),
    .io_response_0_bits(engines_8_io_response_0_bits),
    .io_response_1_ready(engines_8_io_response_1_ready),
    .io_response_1_valid(engines_8_io_response_1_valid),
    .io_response_1_bits(engines_8_io_response_1_bits)
  );
  MonteCarlo_9 engines_9 ( // @[MonteCarlo.scala 254:48]
    .clock(engines_9_clock),
    .reset(engines_9_reset),
    .io_request_0_ready(engines_9_io_request_0_ready),
    .io_request_0_valid(engines_9_io_request_0_valid),
    .io_request_0_bits_time_steps(engines_9_io_request_0_bits_time_steps),
    .io_request_0_bits_start_value(engines_9_io_request_0_bits_start_value),
    .io_request_0_bits_coefficient1(engines_9_io_request_0_bits_coefficient1),
    .io_request_0_bits_coefficient2(engines_9_io_request_0_bits_coefficient2),
    .io_request_1_ready(engines_9_io_request_1_ready),
    .io_request_1_valid(engines_9_io_request_1_valid),
    .io_request_1_bits_time_steps(engines_9_io_request_1_bits_time_steps),
    .io_request_1_bits_start_value(engines_9_io_request_1_bits_start_value),
    .io_request_1_bits_coefficient1(engines_9_io_request_1_bits_coefficient1),
    .io_request_1_bits_coefficient2(engines_9_io_request_1_bits_coefficient2),
    .io_response_0_ready(engines_9_io_response_0_ready),
    .io_response_0_valid(engines_9_io_response_0_valid),
    .io_response_0_bits(engines_9_io_response_0_bits),
    .io_response_1_ready(engines_9_io_response_1_ready),
    .io_response_1_valid(engines_9_io_response_1_valid),
    .io_response_1_bits(engines_9_io_response_1_bits)
  );
  MonteCarlo_10 engines_10 ( // @[MonteCarlo.scala 254:48]
    .clock(engines_10_clock),
    .reset(engines_10_reset),
    .io_request_0_ready(engines_10_io_request_0_ready),
    .io_request_0_valid(engines_10_io_request_0_valid),
    .io_request_0_bits_time_steps(engines_10_io_request_0_bits_time_steps),
    .io_request_0_bits_start_value(engines_10_io_request_0_bits_start_value),
    .io_request_0_bits_coefficient1(engines_10_io_request_0_bits_coefficient1),
    .io_request_0_bits_coefficient2(engines_10_io_request_0_bits_coefficient2),
    .io_request_1_ready(engines_10_io_request_1_ready),
    .io_request_1_valid(engines_10_io_request_1_valid),
    .io_request_1_bits_time_steps(engines_10_io_request_1_bits_time_steps),
    .io_request_1_bits_start_value(engines_10_io_request_1_bits_start_value),
    .io_request_1_bits_coefficient1(engines_10_io_request_1_bits_coefficient1),
    .io_request_1_bits_coefficient2(engines_10_io_request_1_bits_coefficient2),
    .io_response_0_ready(engines_10_io_response_0_ready),
    .io_response_0_valid(engines_10_io_response_0_valid),
    .io_response_0_bits(engines_10_io_response_0_bits),
    .io_response_1_ready(engines_10_io_response_1_ready),
    .io_response_1_valid(engines_10_io_response_1_valid),
    .io_response_1_bits(engines_10_io_response_1_bits)
  );
  MonteCarlo_11 engines_11 ( // @[MonteCarlo.scala 254:48]
    .clock(engines_11_clock),
    .reset(engines_11_reset),
    .io_request_0_ready(engines_11_io_request_0_ready),
    .io_request_0_valid(engines_11_io_request_0_valid),
    .io_request_0_bits_time_steps(engines_11_io_request_0_bits_time_steps),
    .io_request_0_bits_start_value(engines_11_io_request_0_bits_start_value),
    .io_request_0_bits_coefficient1(engines_11_io_request_0_bits_coefficient1),
    .io_request_0_bits_coefficient2(engines_11_io_request_0_bits_coefficient2),
    .io_request_1_ready(engines_11_io_request_1_ready),
    .io_request_1_valid(engines_11_io_request_1_valid),
    .io_request_1_bits_time_steps(engines_11_io_request_1_bits_time_steps),
    .io_request_1_bits_start_value(engines_11_io_request_1_bits_start_value),
    .io_request_1_bits_coefficient1(engines_11_io_request_1_bits_coefficient1),
    .io_request_1_bits_coefficient2(engines_11_io_request_1_bits_coefficient2),
    .io_response_0_ready(engines_11_io_response_0_ready),
    .io_response_0_valid(engines_11_io_response_0_valid),
    .io_response_0_bits(engines_11_io_response_0_bits),
    .io_response_1_ready(engines_11_io_response_1_ready),
    .io_response_1_valid(engines_11_io_response_1_valid),
    .io_response_1_bits(engines_11_io_response_1_bits)
  );
  MonteCarlo_12 engines_12 ( // @[MonteCarlo.scala 254:48]
    .clock(engines_12_clock),
    .reset(engines_12_reset),
    .io_request_0_ready(engines_12_io_request_0_ready),
    .io_request_0_valid(engines_12_io_request_0_valid),
    .io_request_0_bits_time_steps(engines_12_io_request_0_bits_time_steps),
    .io_request_0_bits_start_value(engines_12_io_request_0_bits_start_value),
    .io_request_0_bits_coefficient1(engines_12_io_request_0_bits_coefficient1),
    .io_request_0_bits_coefficient2(engines_12_io_request_0_bits_coefficient2),
    .io_request_1_ready(engines_12_io_request_1_ready),
    .io_request_1_valid(engines_12_io_request_1_valid),
    .io_request_1_bits_time_steps(engines_12_io_request_1_bits_time_steps),
    .io_request_1_bits_start_value(engines_12_io_request_1_bits_start_value),
    .io_request_1_bits_coefficient1(engines_12_io_request_1_bits_coefficient1),
    .io_request_1_bits_coefficient2(engines_12_io_request_1_bits_coefficient2),
    .io_response_0_ready(engines_12_io_response_0_ready),
    .io_response_0_valid(engines_12_io_response_0_valid),
    .io_response_0_bits(engines_12_io_response_0_bits),
    .io_response_1_ready(engines_12_io_response_1_ready),
    .io_response_1_valid(engines_12_io_response_1_valid),
    .io_response_1_bits(engines_12_io_response_1_bits)
  );
  MonteCarlo_13 engines_13 ( // @[MonteCarlo.scala 254:48]
    .clock(engines_13_clock),
    .reset(engines_13_reset),
    .io_request_0_ready(engines_13_io_request_0_ready),
    .io_request_0_valid(engines_13_io_request_0_valid),
    .io_request_0_bits_time_steps(engines_13_io_request_0_bits_time_steps),
    .io_request_0_bits_start_value(engines_13_io_request_0_bits_start_value),
    .io_request_0_bits_coefficient1(engines_13_io_request_0_bits_coefficient1),
    .io_request_0_bits_coefficient2(engines_13_io_request_0_bits_coefficient2),
    .io_request_1_ready(engines_13_io_request_1_ready),
    .io_request_1_valid(engines_13_io_request_1_valid),
    .io_request_1_bits_time_steps(engines_13_io_request_1_bits_time_steps),
    .io_request_1_bits_start_value(engines_13_io_request_1_bits_start_value),
    .io_request_1_bits_coefficient1(engines_13_io_request_1_bits_coefficient1),
    .io_request_1_bits_coefficient2(engines_13_io_request_1_bits_coefficient2),
    .io_response_0_ready(engines_13_io_response_0_ready),
    .io_response_0_valid(engines_13_io_response_0_valid),
    .io_response_0_bits(engines_13_io_response_0_bits),
    .io_response_1_ready(engines_13_io_response_1_ready),
    .io_response_1_valid(engines_13_io_response_1_valid),
    .io_response_1_bits(engines_13_io_response_1_bits)
  );
  MonteCarlo_14 engines_14 ( // @[MonteCarlo.scala 254:48]
    .clock(engines_14_clock),
    .reset(engines_14_reset),
    .io_request_0_ready(engines_14_io_request_0_ready),
    .io_request_0_valid(engines_14_io_request_0_valid),
    .io_request_0_bits_time_steps(engines_14_io_request_0_bits_time_steps),
    .io_request_0_bits_start_value(engines_14_io_request_0_bits_start_value),
    .io_request_0_bits_coefficient1(engines_14_io_request_0_bits_coefficient1),
    .io_request_0_bits_coefficient2(engines_14_io_request_0_bits_coefficient2),
    .io_request_1_ready(engines_14_io_request_1_ready),
    .io_request_1_valid(engines_14_io_request_1_valid),
    .io_request_1_bits_time_steps(engines_14_io_request_1_bits_time_steps),
    .io_request_1_bits_start_value(engines_14_io_request_1_bits_start_value),
    .io_request_1_bits_coefficient1(engines_14_io_request_1_bits_coefficient1),
    .io_request_1_bits_coefficient2(engines_14_io_request_1_bits_coefficient2),
    .io_response_0_ready(engines_14_io_response_0_ready),
    .io_response_0_valid(engines_14_io_response_0_valid),
    .io_response_0_bits(engines_14_io_response_0_bits),
    .io_response_1_ready(engines_14_io_response_1_ready),
    .io_response_1_valid(engines_14_io_response_1_valid),
    .io_response_1_bits(engines_14_io_response_1_bits)
  );
  MonteCarlo_15 engines_15 ( // @[MonteCarlo.scala 254:48]
    .clock(engines_15_clock),
    .reset(engines_15_reset),
    .io_request_0_ready(engines_15_io_request_0_ready),
    .io_request_0_valid(engines_15_io_request_0_valid),
    .io_request_0_bits_time_steps(engines_15_io_request_0_bits_time_steps),
    .io_request_0_bits_start_value(engines_15_io_request_0_bits_start_value),
    .io_request_0_bits_coefficient1(engines_15_io_request_0_bits_coefficient1),
    .io_request_0_bits_coefficient2(engines_15_io_request_0_bits_coefficient2),
    .io_request_1_ready(engines_15_io_request_1_ready),
    .io_request_1_valid(engines_15_io_request_1_valid),
    .io_request_1_bits_time_steps(engines_15_io_request_1_bits_time_steps),
    .io_request_1_bits_start_value(engines_15_io_request_1_bits_start_value),
    .io_request_1_bits_coefficient1(engines_15_io_request_1_bits_coefficient1),
    .io_request_1_bits_coefficient2(engines_15_io_request_1_bits_coefficient2),
    .io_response_0_ready(engines_15_io_response_0_ready),
    .io_response_0_valid(engines_15_io_response_0_valid),
    .io_response_0_bits(engines_15_io_response_0_bits),
    .io_response_1_ready(engines_15_io_response_1_ready),
    .io_response_1_valid(engines_15_io_response_1_valid),
    .io_response_1_bits(engines_15_io_response_1_bits)
  );
  SkidBuffer b1 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_clock),
    .reset(b1_reset),
    .io_enq_ready(b1_io_enq_ready),
    .io_enq_valid(b1_io_enq_valid),
    .io_enq_bits_time_steps(b1_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_io_enq_bits_coefficient2),
    .io_deq_ready(b1_io_deq_ready),
    .io_deq_valid(b1_io_deq_valid),
    .io_deq_bits_time_steps(b1_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_io_deq_bits_coefficient2)
  );
  SkidBuffer b2 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_clock),
    .reset(b2_reset),
    .io_enq_ready(b2_io_enq_ready),
    .io_enq_valid(b2_io_enq_valid),
    .io_enq_bits_time_steps(b2_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_io_enq_bits_coefficient2),
    .io_deq_ready(b2_io_deq_ready),
    .io_deq_valid(b2_io_deq_valid),
    .io_deq_bits_time_steps(b2_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_1 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_1_clock),
    .reset(b1_1_reset),
    .io_enq_ready(b1_1_io_enq_ready),
    .io_enq_valid(b1_1_io_enq_valid),
    .io_enq_bits_time_steps(b1_1_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_1_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_1_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_1_io_enq_bits_coefficient2),
    .io_deq_ready(b1_1_io_deq_ready),
    .io_deq_valid(b1_1_io_deq_valid),
    .io_deq_bits_time_steps(b1_1_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_1_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_1_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_1_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_1 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_1_clock),
    .reset(b2_1_reset),
    .io_enq_ready(b2_1_io_enq_ready),
    .io_enq_valid(b2_1_io_enq_valid),
    .io_enq_bits_time_steps(b2_1_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_1_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_1_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_1_io_enq_bits_coefficient2),
    .io_deq_ready(b2_1_io_deq_ready),
    .io_deq_valid(b2_1_io_deq_valid),
    .io_deq_bits_time_steps(b2_1_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_1_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_1_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_1_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_2 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_2_clock),
    .reset(b1_2_reset),
    .io_enq_ready(b1_2_io_enq_ready),
    .io_enq_valid(b1_2_io_enq_valid),
    .io_enq_bits_time_steps(b1_2_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_2_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_2_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_2_io_enq_bits_coefficient2),
    .io_deq_ready(b1_2_io_deq_ready),
    .io_deq_valid(b1_2_io_deq_valid),
    .io_deq_bits_time_steps(b1_2_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_2_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_2_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_2_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_2 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_2_clock),
    .reset(b2_2_reset),
    .io_enq_ready(b2_2_io_enq_ready),
    .io_enq_valid(b2_2_io_enq_valid),
    .io_enq_bits_time_steps(b2_2_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_2_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_2_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_2_io_enq_bits_coefficient2),
    .io_deq_ready(b2_2_io_deq_ready),
    .io_deq_valid(b2_2_io_deq_valid),
    .io_deq_bits_time_steps(b2_2_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_2_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_2_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_2_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_3 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_3_clock),
    .reset(b1_3_reset),
    .io_enq_ready(b1_3_io_enq_ready),
    .io_enq_valid(b1_3_io_enq_valid),
    .io_enq_bits_time_steps(b1_3_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_3_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_3_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_3_io_enq_bits_coefficient2),
    .io_deq_ready(b1_3_io_deq_ready),
    .io_deq_valid(b1_3_io_deq_valid),
    .io_deq_bits_time_steps(b1_3_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_3_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_3_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_3_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_3 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_3_clock),
    .reset(b2_3_reset),
    .io_enq_ready(b2_3_io_enq_ready),
    .io_enq_valid(b2_3_io_enq_valid),
    .io_enq_bits_time_steps(b2_3_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_3_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_3_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_3_io_enq_bits_coefficient2),
    .io_deq_ready(b2_3_io_deq_ready),
    .io_deq_valid(b2_3_io_deq_valid),
    .io_deq_bits_time_steps(b2_3_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_3_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_3_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_3_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_4 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_4_clock),
    .reset(b1_4_reset),
    .io_enq_ready(b1_4_io_enq_ready),
    .io_enq_valid(b1_4_io_enq_valid),
    .io_enq_bits_time_steps(b1_4_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_4_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_4_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_4_io_enq_bits_coefficient2),
    .io_deq_ready(b1_4_io_deq_ready),
    .io_deq_valid(b1_4_io_deq_valid),
    .io_deq_bits_time_steps(b1_4_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_4_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_4_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_4_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_4 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_4_clock),
    .reset(b2_4_reset),
    .io_enq_ready(b2_4_io_enq_ready),
    .io_enq_valid(b2_4_io_enq_valid),
    .io_enq_bits_time_steps(b2_4_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_4_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_4_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_4_io_enq_bits_coefficient2),
    .io_deq_ready(b2_4_io_deq_ready),
    .io_deq_valid(b2_4_io_deq_valid),
    .io_deq_bits_time_steps(b2_4_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_4_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_4_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_4_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_5 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_5_clock),
    .reset(b1_5_reset),
    .io_enq_ready(b1_5_io_enq_ready),
    .io_enq_valid(b1_5_io_enq_valid),
    .io_enq_bits_time_steps(b1_5_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_5_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_5_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_5_io_enq_bits_coefficient2),
    .io_deq_ready(b1_5_io_deq_ready),
    .io_deq_valid(b1_5_io_deq_valid),
    .io_deq_bits_time_steps(b1_5_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_5_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_5_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_5_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_5 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_5_clock),
    .reset(b2_5_reset),
    .io_enq_ready(b2_5_io_enq_ready),
    .io_enq_valid(b2_5_io_enq_valid),
    .io_enq_bits_time_steps(b2_5_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_5_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_5_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_5_io_enq_bits_coefficient2),
    .io_deq_ready(b2_5_io_deq_ready),
    .io_deq_valid(b2_5_io_deq_valid),
    .io_deq_bits_time_steps(b2_5_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_5_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_5_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_5_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_6 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_6_clock),
    .reset(b1_6_reset),
    .io_enq_ready(b1_6_io_enq_ready),
    .io_enq_valid(b1_6_io_enq_valid),
    .io_enq_bits_time_steps(b1_6_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_6_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_6_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_6_io_enq_bits_coefficient2),
    .io_deq_ready(b1_6_io_deq_ready),
    .io_deq_valid(b1_6_io_deq_valid),
    .io_deq_bits_time_steps(b1_6_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_6_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_6_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_6_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_6 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_6_clock),
    .reset(b2_6_reset),
    .io_enq_ready(b2_6_io_enq_ready),
    .io_enq_valid(b2_6_io_enq_valid),
    .io_enq_bits_time_steps(b2_6_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_6_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_6_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_6_io_enq_bits_coefficient2),
    .io_deq_ready(b2_6_io_deq_ready),
    .io_deq_valid(b2_6_io_deq_valid),
    .io_deq_bits_time_steps(b2_6_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_6_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_6_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_6_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_7 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_7_clock),
    .reset(b1_7_reset),
    .io_enq_ready(b1_7_io_enq_ready),
    .io_enq_valid(b1_7_io_enq_valid),
    .io_enq_bits_time_steps(b1_7_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_7_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_7_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_7_io_enq_bits_coefficient2),
    .io_deq_ready(b1_7_io_deq_ready),
    .io_deq_valid(b1_7_io_deq_valid),
    .io_deq_bits_time_steps(b1_7_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_7_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_7_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_7_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_7 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_7_clock),
    .reset(b2_7_reset),
    .io_enq_ready(b2_7_io_enq_ready),
    .io_enq_valid(b2_7_io_enq_valid),
    .io_enq_bits_time_steps(b2_7_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_7_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_7_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_7_io_enq_bits_coefficient2),
    .io_deq_ready(b2_7_io_deq_ready),
    .io_deq_valid(b2_7_io_deq_valid),
    .io_deq_bits_time_steps(b2_7_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_7_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_7_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_7_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_8 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_8_clock),
    .reset(b1_8_reset),
    .io_enq_ready(b1_8_io_enq_ready),
    .io_enq_valid(b1_8_io_enq_valid),
    .io_enq_bits_time_steps(b1_8_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_8_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_8_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_8_io_enq_bits_coefficient2),
    .io_deq_ready(b1_8_io_deq_ready),
    .io_deq_valid(b1_8_io_deq_valid),
    .io_deq_bits_time_steps(b1_8_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_8_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_8_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_8_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_8 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_8_clock),
    .reset(b2_8_reset),
    .io_enq_ready(b2_8_io_enq_ready),
    .io_enq_valid(b2_8_io_enq_valid),
    .io_enq_bits_time_steps(b2_8_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_8_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_8_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_8_io_enq_bits_coefficient2),
    .io_deq_ready(b2_8_io_deq_ready),
    .io_deq_valid(b2_8_io_deq_valid),
    .io_deq_bits_time_steps(b2_8_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_8_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_8_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_8_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_9 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_9_clock),
    .reset(b1_9_reset),
    .io_enq_ready(b1_9_io_enq_ready),
    .io_enq_valid(b1_9_io_enq_valid),
    .io_enq_bits_time_steps(b1_9_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_9_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_9_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_9_io_enq_bits_coefficient2),
    .io_deq_ready(b1_9_io_deq_ready),
    .io_deq_valid(b1_9_io_deq_valid),
    .io_deq_bits_time_steps(b1_9_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_9_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_9_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_9_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_9 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_9_clock),
    .reset(b2_9_reset),
    .io_enq_ready(b2_9_io_enq_ready),
    .io_enq_valid(b2_9_io_enq_valid),
    .io_enq_bits_time_steps(b2_9_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_9_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_9_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_9_io_enq_bits_coefficient2),
    .io_deq_ready(b2_9_io_deq_ready),
    .io_deq_valid(b2_9_io_deq_valid),
    .io_deq_bits_time_steps(b2_9_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_9_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_9_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_9_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_10 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_10_clock),
    .reset(b1_10_reset),
    .io_enq_ready(b1_10_io_enq_ready),
    .io_enq_valid(b1_10_io_enq_valid),
    .io_enq_bits_time_steps(b1_10_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_10_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_10_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_10_io_enq_bits_coefficient2),
    .io_deq_ready(b1_10_io_deq_ready),
    .io_deq_valid(b1_10_io_deq_valid),
    .io_deq_bits_time_steps(b1_10_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_10_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_10_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_10_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_10 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_10_clock),
    .reset(b2_10_reset),
    .io_enq_ready(b2_10_io_enq_ready),
    .io_enq_valid(b2_10_io_enq_valid),
    .io_enq_bits_time_steps(b2_10_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_10_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_10_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_10_io_enq_bits_coefficient2),
    .io_deq_ready(b2_10_io_deq_ready),
    .io_deq_valid(b2_10_io_deq_valid),
    .io_deq_bits_time_steps(b2_10_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_10_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_10_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_10_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_11 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_11_clock),
    .reset(b1_11_reset),
    .io_enq_ready(b1_11_io_enq_ready),
    .io_enq_valid(b1_11_io_enq_valid),
    .io_enq_bits_time_steps(b1_11_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_11_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_11_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_11_io_enq_bits_coefficient2),
    .io_deq_ready(b1_11_io_deq_ready),
    .io_deq_valid(b1_11_io_deq_valid),
    .io_deq_bits_time_steps(b1_11_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_11_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_11_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_11_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_11 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_11_clock),
    .reset(b2_11_reset),
    .io_enq_ready(b2_11_io_enq_ready),
    .io_enq_valid(b2_11_io_enq_valid),
    .io_enq_bits_time_steps(b2_11_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_11_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_11_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_11_io_enq_bits_coefficient2),
    .io_deq_ready(b2_11_io_deq_ready),
    .io_deq_valid(b2_11_io_deq_valid),
    .io_deq_bits_time_steps(b2_11_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_11_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_11_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_11_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_12 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_12_clock),
    .reset(b1_12_reset),
    .io_enq_ready(b1_12_io_enq_ready),
    .io_enq_valid(b1_12_io_enq_valid),
    .io_enq_bits_time_steps(b1_12_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_12_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_12_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_12_io_enq_bits_coefficient2),
    .io_deq_ready(b1_12_io_deq_ready),
    .io_deq_valid(b1_12_io_deq_valid),
    .io_deq_bits_time_steps(b1_12_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_12_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_12_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_12_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_12 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_12_clock),
    .reset(b2_12_reset),
    .io_enq_ready(b2_12_io_enq_ready),
    .io_enq_valid(b2_12_io_enq_valid),
    .io_enq_bits_time_steps(b2_12_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_12_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_12_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_12_io_enq_bits_coefficient2),
    .io_deq_ready(b2_12_io_deq_ready),
    .io_deq_valid(b2_12_io_deq_valid),
    .io_deq_bits_time_steps(b2_12_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_12_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_12_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_12_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_13 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_13_clock),
    .reset(b1_13_reset),
    .io_enq_ready(b1_13_io_enq_ready),
    .io_enq_valid(b1_13_io_enq_valid),
    .io_enq_bits_time_steps(b1_13_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_13_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_13_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_13_io_enq_bits_coefficient2),
    .io_deq_ready(b1_13_io_deq_ready),
    .io_deq_valid(b1_13_io_deq_valid),
    .io_deq_bits_time_steps(b1_13_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_13_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_13_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_13_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_13 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_13_clock),
    .reset(b2_13_reset),
    .io_enq_ready(b2_13_io_enq_ready),
    .io_enq_valid(b2_13_io_enq_valid),
    .io_enq_bits_time_steps(b2_13_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_13_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_13_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_13_io_enq_bits_coefficient2),
    .io_deq_ready(b2_13_io_deq_ready),
    .io_deq_valid(b2_13_io_deq_valid),
    .io_deq_bits_time_steps(b2_13_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_13_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_13_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_13_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_14 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_14_clock),
    .reset(b1_14_reset),
    .io_enq_ready(b1_14_io_enq_ready),
    .io_enq_valid(b1_14_io_enq_valid),
    .io_enq_bits_time_steps(b1_14_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_14_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_14_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_14_io_enq_bits_coefficient2),
    .io_deq_ready(b1_14_io_deq_ready),
    .io_deq_valid(b1_14_io_deq_valid),
    .io_deq_bits_time_steps(b1_14_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_14_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_14_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_14_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_14 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_14_clock),
    .reset(b2_14_reset),
    .io_enq_ready(b2_14_io_enq_ready),
    .io_enq_valid(b2_14_io_enq_valid),
    .io_enq_bits_time_steps(b2_14_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_14_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_14_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_14_io_enq_bits_coefficient2),
    .io_deq_ready(b2_14_io_deq_ready),
    .io_deq_valid(b2_14_io_deq_valid),
    .io_deq_bits_time_steps(b2_14_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_14_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_14_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_14_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_15 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_15_clock),
    .reset(b1_15_reset),
    .io_enq_ready(b1_15_io_enq_ready),
    .io_enq_valid(b1_15_io_enq_valid),
    .io_enq_bits_time_steps(b1_15_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_15_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_15_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_15_io_enq_bits_coefficient2),
    .io_deq_ready(b1_15_io_deq_ready),
    .io_deq_valid(b1_15_io_deq_valid),
    .io_deq_bits_time_steps(b1_15_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_15_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_15_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_15_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_15 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_15_clock),
    .reset(b2_15_reset),
    .io_enq_ready(b2_15_io_enq_ready),
    .io_enq_valid(b2_15_io_enq_valid),
    .io_enq_bits_time_steps(b2_15_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_15_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_15_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_15_io_enq_bits_coefficient2),
    .io_deq_ready(b2_15_io_deq_ready),
    .io_deq_valid(b2_15_io_deq_valid),
    .io_deq_bits_time_steps(b2_15_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_15_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_15_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_15_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_16 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_16_clock),
    .reset(b1_16_reset),
    .io_enq_ready(b1_16_io_enq_ready),
    .io_enq_valid(b1_16_io_enq_valid),
    .io_enq_bits_time_steps(b1_16_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_16_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_16_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_16_io_enq_bits_coefficient2),
    .io_deq_ready(b1_16_io_deq_ready),
    .io_deq_valid(b1_16_io_deq_valid),
    .io_deq_bits_time_steps(b1_16_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_16_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_16_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_16_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_16 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_16_clock),
    .reset(b2_16_reset),
    .io_enq_ready(b2_16_io_enq_ready),
    .io_enq_valid(b2_16_io_enq_valid),
    .io_enq_bits_time_steps(b2_16_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_16_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_16_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_16_io_enq_bits_coefficient2),
    .io_deq_ready(b2_16_io_deq_ready),
    .io_deq_valid(b2_16_io_deq_valid),
    .io_deq_bits_time_steps(b2_16_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_16_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_16_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_16_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_17 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_17_clock),
    .reset(b1_17_reset),
    .io_enq_ready(b1_17_io_enq_ready),
    .io_enq_valid(b1_17_io_enq_valid),
    .io_enq_bits_time_steps(b1_17_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_17_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_17_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_17_io_enq_bits_coefficient2),
    .io_deq_ready(b1_17_io_deq_ready),
    .io_deq_valid(b1_17_io_deq_valid),
    .io_deq_bits_time_steps(b1_17_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_17_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_17_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_17_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_17 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_17_clock),
    .reset(b2_17_reset),
    .io_enq_ready(b2_17_io_enq_ready),
    .io_enq_valid(b2_17_io_enq_valid),
    .io_enq_bits_time_steps(b2_17_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_17_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_17_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_17_io_enq_bits_coefficient2),
    .io_deq_ready(b2_17_io_deq_ready),
    .io_deq_valid(b2_17_io_deq_valid),
    .io_deq_bits_time_steps(b2_17_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_17_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_17_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_17_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_18 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_18_clock),
    .reset(b1_18_reset),
    .io_enq_ready(b1_18_io_enq_ready),
    .io_enq_valid(b1_18_io_enq_valid),
    .io_enq_bits_time_steps(b1_18_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_18_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_18_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_18_io_enq_bits_coefficient2),
    .io_deq_ready(b1_18_io_deq_ready),
    .io_deq_valid(b1_18_io_deq_valid),
    .io_deq_bits_time_steps(b1_18_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_18_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_18_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_18_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_18 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_18_clock),
    .reset(b2_18_reset),
    .io_enq_ready(b2_18_io_enq_ready),
    .io_enq_valid(b2_18_io_enq_valid),
    .io_enq_bits_time_steps(b2_18_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_18_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_18_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_18_io_enq_bits_coefficient2),
    .io_deq_ready(b2_18_io_deq_ready),
    .io_deq_valid(b2_18_io_deq_valid),
    .io_deq_bits_time_steps(b2_18_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_18_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_18_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_18_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_19 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_19_clock),
    .reset(b1_19_reset),
    .io_enq_ready(b1_19_io_enq_ready),
    .io_enq_valid(b1_19_io_enq_valid),
    .io_enq_bits_time_steps(b1_19_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_19_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_19_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_19_io_enq_bits_coefficient2),
    .io_deq_ready(b1_19_io_deq_ready),
    .io_deq_valid(b1_19_io_deq_valid),
    .io_deq_bits_time_steps(b1_19_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_19_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_19_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_19_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_19 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_19_clock),
    .reset(b2_19_reset),
    .io_enq_ready(b2_19_io_enq_ready),
    .io_enq_valid(b2_19_io_enq_valid),
    .io_enq_bits_time_steps(b2_19_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_19_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_19_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_19_io_enq_bits_coefficient2),
    .io_deq_ready(b2_19_io_deq_ready),
    .io_deq_valid(b2_19_io_deq_valid),
    .io_deq_bits_time_steps(b2_19_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_19_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_19_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_19_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_20 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_20_clock),
    .reset(b1_20_reset),
    .io_enq_ready(b1_20_io_enq_ready),
    .io_enq_valid(b1_20_io_enq_valid),
    .io_enq_bits_time_steps(b1_20_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_20_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_20_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_20_io_enq_bits_coefficient2),
    .io_deq_ready(b1_20_io_deq_ready),
    .io_deq_valid(b1_20_io_deq_valid),
    .io_deq_bits_time_steps(b1_20_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_20_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_20_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_20_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_20 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_20_clock),
    .reset(b2_20_reset),
    .io_enq_ready(b2_20_io_enq_ready),
    .io_enq_valid(b2_20_io_enq_valid),
    .io_enq_bits_time_steps(b2_20_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_20_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_20_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_20_io_enq_bits_coefficient2),
    .io_deq_ready(b2_20_io_deq_ready),
    .io_deq_valid(b2_20_io_deq_valid),
    .io_deq_bits_time_steps(b2_20_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_20_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_20_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_20_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_21 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_21_clock),
    .reset(b1_21_reset),
    .io_enq_ready(b1_21_io_enq_ready),
    .io_enq_valid(b1_21_io_enq_valid),
    .io_enq_bits_time_steps(b1_21_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_21_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_21_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_21_io_enq_bits_coefficient2),
    .io_deq_ready(b1_21_io_deq_ready),
    .io_deq_valid(b1_21_io_deq_valid),
    .io_deq_bits_time_steps(b1_21_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_21_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_21_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_21_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_21 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_21_clock),
    .reset(b2_21_reset),
    .io_enq_ready(b2_21_io_enq_ready),
    .io_enq_valid(b2_21_io_enq_valid),
    .io_enq_bits_time_steps(b2_21_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_21_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_21_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_21_io_enq_bits_coefficient2),
    .io_deq_ready(b2_21_io_deq_ready),
    .io_deq_valid(b2_21_io_deq_valid),
    .io_deq_bits_time_steps(b2_21_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_21_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_21_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_21_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_22 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_22_clock),
    .reset(b1_22_reset),
    .io_enq_ready(b1_22_io_enq_ready),
    .io_enq_valid(b1_22_io_enq_valid),
    .io_enq_bits_time_steps(b1_22_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_22_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_22_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_22_io_enq_bits_coefficient2),
    .io_deq_ready(b1_22_io_deq_ready),
    .io_deq_valid(b1_22_io_deq_valid),
    .io_deq_bits_time_steps(b1_22_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_22_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_22_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_22_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_22 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_22_clock),
    .reset(b2_22_reset),
    .io_enq_ready(b2_22_io_enq_ready),
    .io_enq_valid(b2_22_io_enq_valid),
    .io_enq_bits_time_steps(b2_22_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_22_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_22_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_22_io_enq_bits_coefficient2),
    .io_deq_ready(b2_22_io_deq_ready),
    .io_deq_valid(b2_22_io_deq_valid),
    .io_deq_bits_time_steps(b2_22_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_22_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_22_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_22_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_23 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_23_clock),
    .reset(b1_23_reset),
    .io_enq_ready(b1_23_io_enq_ready),
    .io_enq_valid(b1_23_io_enq_valid),
    .io_enq_bits_time_steps(b1_23_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_23_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_23_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_23_io_enq_bits_coefficient2),
    .io_deq_ready(b1_23_io_deq_ready),
    .io_deq_valid(b1_23_io_deq_valid),
    .io_deq_bits_time_steps(b1_23_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_23_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_23_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_23_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_23 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_23_clock),
    .reset(b2_23_reset),
    .io_enq_ready(b2_23_io_enq_ready),
    .io_enq_valid(b2_23_io_enq_valid),
    .io_enq_bits_time_steps(b2_23_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_23_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_23_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_23_io_enq_bits_coefficient2),
    .io_deq_ready(b2_23_io_deq_ready),
    .io_deq_valid(b2_23_io_deq_valid),
    .io_deq_bits_time_steps(b2_23_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_23_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_23_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_23_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_24 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_24_clock),
    .reset(b1_24_reset),
    .io_enq_ready(b1_24_io_enq_ready),
    .io_enq_valid(b1_24_io_enq_valid),
    .io_enq_bits_time_steps(b1_24_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_24_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_24_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_24_io_enq_bits_coefficient2),
    .io_deq_ready(b1_24_io_deq_ready),
    .io_deq_valid(b1_24_io_deq_valid),
    .io_deq_bits_time_steps(b1_24_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_24_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_24_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_24_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_24 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_24_clock),
    .reset(b2_24_reset),
    .io_enq_ready(b2_24_io_enq_ready),
    .io_enq_valid(b2_24_io_enq_valid),
    .io_enq_bits_time_steps(b2_24_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_24_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_24_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_24_io_enq_bits_coefficient2),
    .io_deq_ready(b2_24_io_deq_ready),
    .io_deq_valid(b2_24_io_deq_valid),
    .io_deq_bits_time_steps(b2_24_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_24_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_24_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_24_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_25 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_25_clock),
    .reset(b1_25_reset),
    .io_enq_ready(b1_25_io_enq_ready),
    .io_enq_valid(b1_25_io_enq_valid),
    .io_enq_bits_time_steps(b1_25_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_25_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_25_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_25_io_enq_bits_coefficient2),
    .io_deq_ready(b1_25_io_deq_ready),
    .io_deq_valid(b1_25_io_deq_valid),
    .io_deq_bits_time_steps(b1_25_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_25_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_25_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_25_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_25 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_25_clock),
    .reset(b2_25_reset),
    .io_enq_ready(b2_25_io_enq_ready),
    .io_enq_valid(b2_25_io_enq_valid),
    .io_enq_bits_time_steps(b2_25_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_25_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_25_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_25_io_enq_bits_coefficient2),
    .io_deq_ready(b2_25_io_deq_ready),
    .io_deq_valid(b2_25_io_deq_valid),
    .io_deq_bits_time_steps(b2_25_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_25_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_25_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_25_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_26 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_26_clock),
    .reset(b1_26_reset),
    .io_enq_ready(b1_26_io_enq_ready),
    .io_enq_valid(b1_26_io_enq_valid),
    .io_enq_bits_time_steps(b1_26_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_26_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_26_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_26_io_enq_bits_coefficient2),
    .io_deq_ready(b1_26_io_deq_ready),
    .io_deq_valid(b1_26_io_deq_valid),
    .io_deq_bits_time_steps(b1_26_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_26_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_26_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_26_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_26 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_26_clock),
    .reset(b2_26_reset),
    .io_enq_ready(b2_26_io_enq_ready),
    .io_enq_valid(b2_26_io_enq_valid),
    .io_enq_bits_time_steps(b2_26_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_26_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_26_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_26_io_enq_bits_coefficient2),
    .io_deq_ready(b2_26_io_deq_ready),
    .io_deq_valid(b2_26_io_deq_valid),
    .io_deq_bits_time_steps(b2_26_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_26_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_26_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_26_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_27 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_27_clock),
    .reset(b1_27_reset),
    .io_enq_ready(b1_27_io_enq_ready),
    .io_enq_valid(b1_27_io_enq_valid),
    .io_enq_bits_time_steps(b1_27_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_27_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_27_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_27_io_enq_bits_coefficient2),
    .io_deq_ready(b1_27_io_deq_ready),
    .io_deq_valid(b1_27_io_deq_valid),
    .io_deq_bits_time_steps(b1_27_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_27_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_27_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_27_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_27 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_27_clock),
    .reset(b2_27_reset),
    .io_enq_ready(b2_27_io_enq_ready),
    .io_enq_valid(b2_27_io_enq_valid),
    .io_enq_bits_time_steps(b2_27_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_27_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_27_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_27_io_enq_bits_coefficient2),
    .io_deq_ready(b2_27_io_deq_ready),
    .io_deq_valid(b2_27_io_deq_valid),
    .io_deq_bits_time_steps(b2_27_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_27_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_27_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_27_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_28 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_28_clock),
    .reset(b1_28_reset),
    .io_enq_ready(b1_28_io_enq_ready),
    .io_enq_valid(b1_28_io_enq_valid),
    .io_enq_bits_time_steps(b1_28_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_28_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_28_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_28_io_enq_bits_coefficient2),
    .io_deq_ready(b1_28_io_deq_ready),
    .io_deq_valid(b1_28_io_deq_valid),
    .io_deq_bits_time_steps(b1_28_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_28_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_28_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_28_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_28 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_28_clock),
    .reset(b2_28_reset),
    .io_enq_ready(b2_28_io_enq_ready),
    .io_enq_valid(b2_28_io_enq_valid),
    .io_enq_bits_time_steps(b2_28_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_28_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_28_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_28_io_enq_bits_coefficient2),
    .io_deq_ready(b2_28_io_deq_ready),
    .io_deq_valid(b2_28_io_deq_valid),
    .io_deq_bits_time_steps(b2_28_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_28_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_28_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_28_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_29 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_29_clock),
    .reset(b1_29_reset),
    .io_enq_ready(b1_29_io_enq_ready),
    .io_enq_valid(b1_29_io_enq_valid),
    .io_enq_bits_time_steps(b1_29_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_29_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_29_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_29_io_enq_bits_coefficient2),
    .io_deq_ready(b1_29_io_deq_ready),
    .io_deq_valid(b1_29_io_deq_valid),
    .io_deq_bits_time_steps(b1_29_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_29_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_29_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_29_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_29 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_29_clock),
    .reset(b2_29_reset),
    .io_enq_ready(b2_29_io_enq_ready),
    .io_enq_valid(b2_29_io_enq_valid),
    .io_enq_bits_time_steps(b2_29_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_29_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_29_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_29_io_enq_bits_coefficient2),
    .io_deq_ready(b2_29_io_deq_ready),
    .io_deq_valid(b2_29_io_deq_valid),
    .io_deq_bits_time_steps(b2_29_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_29_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_29_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_29_io_deq_bits_coefficient2)
  );
  SkidBuffer b1_30 ( // @[MonteCarlo.scala 239:27]
    .clock(b1_30_clock),
    .reset(b1_30_reset),
    .io_enq_ready(b1_30_io_enq_ready),
    .io_enq_valid(b1_30_io_enq_valid),
    .io_enq_bits_time_steps(b1_30_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b1_30_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b1_30_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b1_30_io_enq_bits_coefficient2),
    .io_deq_ready(b1_30_io_deq_ready),
    .io_deq_valid(b1_30_io_deq_valid),
    .io_deq_bits_time_steps(b1_30_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b1_30_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b1_30_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b1_30_io_deq_bits_coefficient2)
  );
  SkidBuffer b2_30 ( // @[MonteCarlo.scala 240:27]
    .clock(b2_30_clock),
    .reset(b2_30_reset),
    .io_enq_ready(b2_30_io_enq_ready),
    .io_enq_valid(b2_30_io_enq_valid),
    .io_enq_bits_time_steps(b2_30_io_enq_bits_time_steps),
    .io_enq_bits_start_value(b2_30_io_enq_bits_start_value),
    .io_enq_bits_coefficient1(b2_30_io_enq_bits_coefficient1),
    .io_enq_bits_coefficient2(b2_30_io_enq_bits_coefficient2),
    .io_deq_ready(b2_30_io_deq_ready),
    .io_deq_valid(b2_30_io_deq_valid),
    .io_deq_bits_time_steps(b2_30_io_deq_bits_time_steps),
    .io_deq_bits_start_value(b2_30_io_deq_bits_start_value),
    .io_deq_bits_coefficient1(b2_30_io_deq_bits_coefficient1),
    .io_deq_bits_coefficient2(b2_30_io_deq_bits_coefficient2)
  );
  PipelinedMean partial_result_impl ( // @[MonteCarlo.scala 215:22]
    .clock(partial_result_impl_clock),
    .reset(partial_result_impl_reset),
    .io_lanes_0_ready(partial_result_impl_io_lanes_0_ready),
    .io_lanes_0_valid(partial_result_impl_io_lanes_0_valid),
    .io_lanes_0_bits(partial_result_impl_io_lanes_0_bits),
    .io_lanes_1_ready(partial_result_impl_io_lanes_1_ready),
    .io_lanes_1_valid(partial_result_impl_io_lanes_1_valid),
    .io_lanes_1_bits(partial_result_impl_io_lanes_1_bits),
    .io_lanes_2_ready(partial_result_impl_io_lanes_2_ready),
    .io_lanes_2_valid(partial_result_impl_io_lanes_2_valid),
    .io_lanes_2_bits(partial_result_impl_io_lanes_2_bits),
    .io_lanes_3_ready(partial_result_impl_io_lanes_3_ready),
    .io_lanes_3_valid(partial_result_impl_io_lanes_3_valid),
    .io_lanes_3_bits(partial_result_impl_io_lanes_3_bits),
    .io_lanes_4_ready(partial_result_impl_io_lanes_4_ready),
    .io_lanes_4_valid(partial_result_impl_io_lanes_4_valid),
    .io_lanes_4_bits(partial_result_impl_io_lanes_4_bits),
    .io_lanes_5_ready(partial_result_impl_io_lanes_5_ready),
    .io_lanes_5_valid(partial_result_impl_io_lanes_5_valid),
    .io_lanes_5_bits(partial_result_impl_io_lanes_5_bits),
    .io_lanes_6_ready(partial_result_impl_io_lanes_6_ready),
    .io_lanes_6_valid(partial_result_impl_io_lanes_6_valid),
    .io_lanes_6_bits(partial_result_impl_io_lanes_6_bits),
    .io_lanes_7_ready(partial_result_impl_io_lanes_7_ready),
    .io_lanes_7_valid(partial_result_impl_io_lanes_7_valid),
    .io_lanes_7_bits(partial_result_impl_io_lanes_7_bits),
    .io_lanes_8_ready(partial_result_impl_io_lanes_8_ready),
    .io_lanes_8_valid(partial_result_impl_io_lanes_8_valid),
    .io_lanes_8_bits(partial_result_impl_io_lanes_8_bits),
    .io_lanes_9_ready(partial_result_impl_io_lanes_9_ready),
    .io_lanes_9_valid(partial_result_impl_io_lanes_9_valid),
    .io_lanes_9_bits(partial_result_impl_io_lanes_9_bits),
    .io_lanes_10_ready(partial_result_impl_io_lanes_10_ready),
    .io_lanes_10_valid(partial_result_impl_io_lanes_10_valid),
    .io_lanes_10_bits(partial_result_impl_io_lanes_10_bits),
    .io_lanes_11_ready(partial_result_impl_io_lanes_11_ready),
    .io_lanes_11_valid(partial_result_impl_io_lanes_11_valid),
    .io_lanes_11_bits(partial_result_impl_io_lanes_11_bits),
    .io_lanes_12_ready(partial_result_impl_io_lanes_12_ready),
    .io_lanes_12_valid(partial_result_impl_io_lanes_12_valid),
    .io_lanes_12_bits(partial_result_impl_io_lanes_12_bits),
    .io_lanes_13_ready(partial_result_impl_io_lanes_13_ready),
    .io_lanes_13_valid(partial_result_impl_io_lanes_13_valid),
    .io_lanes_13_bits(partial_result_impl_io_lanes_13_bits),
    .io_lanes_14_ready(partial_result_impl_io_lanes_14_ready),
    .io_lanes_14_valid(partial_result_impl_io_lanes_14_valid),
    .io_lanes_14_bits(partial_result_impl_io_lanes_14_bits),
    .io_lanes_15_ready(partial_result_impl_io_lanes_15_ready),
    .io_lanes_15_valid(partial_result_impl_io_lanes_15_valid),
    .io_lanes_15_bits(partial_result_impl_io_lanes_15_bits),
    .io_lanes_16_ready(partial_result_impl_io_lanes_16_ready),
    .io_lanes_16_valid(partial_result_impl_io_lanes_16_valid),
    .io_lanes_16_bits(partial_result_impl_io_lanes_16_bits),
    .io_lanes_17_ready(partial_result_impl_io_lanes_17_ready),
    .io_lanes_17_valid(partial_result_impl_io_lanes_17_valid),
    .io_lanes_17_bits(partial_result_impl_io_lanes_17_bits),
    .io_lanes_18_ready(partial_result_impl_io_lanes_18_ready),
    .io_lanes_18_valid(partial_result_impl_io_lanes_18_valid),
    .io_lanes_18_bits(partial_result_impl_io_lanes_18_bits),
    .io_lanes_19_ready(partial_result_impl_io_lanes_19_ready),
    .io_lanes_19_valid(partial_result_impl_io_lanes_19_valid),
    .io_lanes_19_bits(partial_result_impl_io_lanes_19_bits),
    .io_lanes_20_ready(partial_result_impl_io_lanes_20_ready),
    .io_lanes_20_valid(partial_result_impl_io_lanes_20_valid),
    .io_lanes_20_bits(partial_result_impl_io_lanes_20_bits),
    .io_lanes_21_ready(partial_result_impl_io_lanes_21_ready),
    .io_lanes_21_valid(partial_result_impl_io_lanes_21_valid),
    .io_lanes_21_bits(partial_result_impl_io_lanes_21_bits),
    .io_lanes_22_ready(partial_result_impl_io_lanes_22_ready),
    .io_lanes_22_valid(partial_result_impl_io_lanes_22_valid),
    .io_lanes_22_bits(partial_result_impl_io_lanes_22_bits),
    .io_lanes_23_ready(partial_result_impl_io_lanes_23_ready),
    .io_lanes_23_valid(partial_result_impl_io_lanes_23_valid),
    .io_lanes_23_bits(partial_result_impl_io_lanes_23_bits),
    .io_lanes_24_ready(partial_result_impl_io_lanes_24_ready),
    .io_lanes_24_valid(partial_result_impl_io_lanes_24_valid),
    .io_lanes_24_bits(partial_result_impl_io_lanes_24_bits),
    .io_lanes_25_ready(partial_result_impl_io_lanes_25_ready),
    .io_lanes_25_valid(partial_result_impl_io_lanes_25_valid),
    .io_lanes_25_bits(partial_result_impl_io_lanes_25_bits),
    .io_lanes_26_ready(partial_result_impl_io_lanes_26_ready),
    .io_lanes_26_valid(partial_result_impl_io_lanes_26_valid),
    .io_lanes_26_bits(partial_result_impl_io_lanes_26_bits),
    .io_lanes_27_ready(partial_result_impl_io_lanes_27_ready),
    .io_lanes_27_valid(partial_result_impl_io_lanes_27_valid),
    .io_lanes_27_bits(partial_result_impl_io_lanes_27_bits),
    .io_lanes_28_ready(partial_result_impl_io_lanes_28_ready),
    .io_lanes_28_valid(partial_result_impl_io_lanes_28_valid),
    .io_lanes_28_bits(partial_result_impl_io_lanes_28_bits),
    .io_lanes_29_ready(partial_result_impl_io_lanes_29_ready),
    .io_lanes_29_valid(partial_result_impl_io_lanes_29_valid),
    .io_lanes_29_bits(partial_result_impl_io_lanes_29_bits),
    .io_lanes_30_ready(partial_result_impl_io_lanes_30_ready),
    .io_lanes_30_valid(partial_result_impl_io_lanes_30_valid),
    .io_lanes_30_bits(partial_result_impl_io_lanes_30_bits),
    .io_lanes_31_ready(partial_result_impl_io_lanes_31_ready),
    .io_lanes_31_valid(partial_result_impl_io_lanes_31_valid),
    .io_lanes_31_bits(partial_result_impl_io_lanes_31_bits),
    .io_result_ready(partial_result_impl_io_result_ready),
    .io_result_valid(partial_result_impl_io_result_valid),
    .io_result_bits(partial_result_impl_io_result_bits)
  );
  assign io_request_ready = b1_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign io_response_valid = partial_result_impl_io_result_valid; // @[MonteCarlo.scala 259:15]
  assign io_response_bits = partial_result_impl_io_result_bits; // @[MonteCarlo.scala 259:15]
  assign engines_0_clock = clock;
  assign engines_0_reset = reset;
  assign engines_0_io_request_0_valid = b1_15_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_0_io_request_0_bits_time_steps = b1_15_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_0_io_request_0_bits_start_value = b1_15_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_0_io_request_0_bits_coefficient1 = b1_15_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_0_io_request_0_bits_coefficient2 = b1_15_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_0_io_request_1_valid = b2_15_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_0_io_request_1_bits_time_steps = b2_15_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_0_io_request_1_bits_start_value = b2_15_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_0_io_request_1_bits_coefficient1 = b2_15_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_0_io_request_1_bits_coefficient2 = b2_15_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_0_io_response_0_ready = partial_result_impl_io_lanes_0_ready; // @[MonteCarlo.scala 216:19]
  assign engines_0_io_response_1_ready = partial_result_impl_io_lanes_1_ready; // @[MonteCarlo.scala 216:19]
  assign engines_1_clock = clock;
  assign engines_1_reset = reset;
  assign engines_1_io_request_0_valid = b1_16_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_1_io_request_0_bits_time_steps = b1_16_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_1_io_request_0_bits_start_value = b1_16_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_1_io_request_0_bits_coefficient1 = b1_16_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_1_io_request_0_bits_coefficient2 = b1_16_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_1_io_request_1_valid = b2_16_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_1_io_request_1_bits_time_steps = b2_16_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_1_io_request_1_bits_start_value = b2_16_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_1_io_request_1_bits_coefficient1 = b2_16_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_1_io_request_1_bits_coefficient2 = b2_16_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_1_io_response_0_ready = partial_result_impl_io_lanes_2_ready; // @[MonteCarlo.scala 216:19]
  assign engines_1_io_response_1_ready = partial_result_impl_io_lanes_3_ready; // @[MonteCarlo.scala 216:19]
  assign engines_2_clock = clock;
  assign engines_2_reset = reset;
  assign engines_2_io_request_0_valid = b1_17_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_2_io_request_0_bits_time_steps = b1_17_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_2_io_request_0_bits_start_value = b1_17_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_2_io_request_0_bits_coefficient1 = b1_17_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_2_io_request_0_bits_coefficient2 = b1_17_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_2_io_request_1_valid = b2_17_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_2_io_request_1_bits_time_steps = b2_17_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_2_io_request_1_bits_start_value = b2_17_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_2_io_request_1_bits_coefficient1 = b2_17_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_2_io_request_1_bits_coefficient2 = b2_17_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_2_io_response_0_ready = partial_result_impl_io_lanes_4_ready; // @[MonteCarlo.scala 216:19]
  assign engines_2_io_response_1_ready = partial_result_impl_io_lanes_5_ready; // @[MonteCarlo.scala 216:19]
  assign engines_3_clock = clock;
  assign engines_3_reset = reset;
  assign engines_3_io_request_0_valid = b1_18_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_3_io_request_0_bits_time_steps = b1_18_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_3_io_request_0_bits_start_value = b1_18_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_3_io_request_0_bits_coefficient1 = b1_18_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_3_io_request_0_bits_coefficient2 = b1_18_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_3_io_request_1_valid = b2_18_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_3_io_request_1_bits_time_steps = b2_18_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_3_io_request_1_bits_start_value = b2_18_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_3_io_request_1_bits_coefficient1 = b2_18_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_3_io_request_1_bits_coefficient2 = b2_18_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_3_io_response_0_ready = partial_result_impl_io_lanes_6_ready; // @[MonteCarlo.scala 216:19]
  assign engines_3_io_response_1_ready = partial_result_impl_io_lanes_7_ready; // @[MonteCarlo.scala 216:19]
  assign engines_4_clock = clock;
  assign engines_4_reset = reset;
  assign engines_4_io_request_0_valid = b1_19_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_4_io_request_0_bits_time_steps = b1_19_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_4_io_request_0_bits_start_value = b1_19_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_4_io_request_0_bits_coefficient1 = b1_19_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_4_io_request_0_bits_coefficient2 = b1_19_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_4_io_request_1_valid = b2_19_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_4_io_request_1_bits_time_steps = b2_19_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_4_io_request_1_bits_start_value = b2_19_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_4_io_request_1_bits_coefficient1 = b2_19_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_4_io_request_1_bits_coefficient2 = b2_19_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_4_io_response_0_ready = partial_result_impl_io_lanes_8_ready; // @[MonteCarlo.scala 216:19]
  assign engines_4_io_response_1_ready = partial_result_impl_io_lanes_9_ready; // @[MonteCarlo.scala 216:19]
  assign engines_5_clock = clock;
  assign engines_5_reset = reset;
  assign engines_5_io_request_0_valid = b1_20_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_5_io_request_0_bits_time_steps = b1_20_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_5_io_request_0_bits_start_value = b1_20_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_5_io_request_0_bits_coefficient1 = b1_20_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_5_io_request_0_bits_coefficient2 = b1_20_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_5_io_request_1_valid = b2_20_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_5_io_request_1_bits_time_steps = b2_20_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_5_io_request_1_bits_start_value = b2_20_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_5_io_request_1_bits_coefficient1 = b2_20_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_5_io_request_1_bits_coefficient2 = b2_20_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_5_io_response_0_ready = partial_result_impl_io_lanes_10_ready; // @[MonteCarlo.scala 216:19]
  assign engines_5_io_response_1_ready = partial_result_impl_io_lanes_11_ready; // @[MonteCarlo.scala 216:19]
  assign engines_6_clock = clock;
  assign engines_6_reset = reset;
  assign engines_6_io_request_0_valid = b1_21_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_6_io_request_0_bits_time_steps = b1_21_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_6_io_request_0_bits_start_value = b1_21_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_6_io_request_0_bits_coefficient1 = b1_21_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_6_io_request_0_bits_coefficient2 = b1_21_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_6_io_request_1_valid = b2_21_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_6_io_request_1_bits_time_steps = b2_21_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_6_io_request_1_bits_start_value = b2_21_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_6_io_request_1_bits_coefficient1 = b2_21_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_6_io_request_1_bits_coefficient2 = b2_21_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_6_io_response_0_ready = partial_result_impl_io_lanes_12_ready; // @[MonteCarlo.scala 216:19]
  assign engines_6_io_response_1_ready = partial_result_impl_io_lanes_13_ready; // @[MonteCarlo.scala 216:19]
  assign engines_7_clock = clock;
  assign engines_7_reset = reset;
  assign engines_7_io_request_0_valid = b1_22_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_7_io_request_0_bits_time_steps = b1_22_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_7_io_request_0_bits_start_value = b1_22_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_7_io_request_0_bits_coefficient1 = b1_22_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_7_io_request_0_bits_coefficient2 = b1_22_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_7_io_request_1_valid = b2_22_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_7_io_request_1_bits_time_steps = b2_22_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_7_io_request_1_bits_start_value = b2_22_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_7_io_request_1_bits_coefficient1 = b2_22_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_7_io_request_1_bits_coefficient2 = b2_22_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_7_io_response_0_ready = partial_result_impl_io_lanes_14_ready; // @[MonteCarlo.scala 216:19]
  assign engines_7_io_response_1_ready = partial_result_impl_io_lanes_15_ready; // @[MonteCarlo.scala 216:19]
  assign engines_8_clock = clock;
  assign engines_8_reset = reset;
  assign engines_8_io_request_0_valid = b1_23_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_8_io_request_0_bits_time_steps = b1_23_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_8_io_request_0_bits_start_value = b1_23_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_8_io_request_0_bits_coefficient1 = b1_23_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_8_io_request_0_bits_coefficient2 = b1_23_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_8_io_request_1_valid = b2_23_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_8_io_request_1_bits_time_steps = b2_23_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_8_io_request_1_bits_start_value = b2_23_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_8_io_request_1_bits_coefficient1 = b2_23_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_8_io_request_1_bits_coefficient2 = b2_23_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_8_io_response_0_ready = partial_result_impl_io_lanes_16_ready; // @[MonteCarlo.scala 216:19]
  assign engines_8_io_response_1_ready = partial_result_impl_io_lanes_17_ready; // @[MonteCarlo.scala 216:19]
  assign engines_9_clock = clock;
  assign engines_9_reset = reset;
  assign engines_9_io_request_0_valid = b1_24_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_9_io_request_0_bits_time_steps = b1_24_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_9_io_request_0_bits_start_value = b1_24_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_9_io_request_0_bits_coefficient1 = b1_24_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_9_io_request_0_bits_coefficient2 = b1_24_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_9_io_request_1_valid = b2_24_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_9_io_request_1_bits_time_steps = b2_24_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_9_io_request_1_bits_start_value = b2_24_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_9_io_request_1_bits_coefficient1 = b2_24_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_9_io_request_1_bits_coefficient2 = b2_24_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_9_io_response_0_ready = partial_result_impl_io_lanes_18_ready; // @[MonteCarlo.scala 216:19]
  assign engines_9_io_response_1_ready = partial_result_impl_io_lanes_19_ready; // @[MonteCarlo.scala 216:19]
  assign engines_10_clock = clock;
  assign engines_10_reset = reset;
  assign engines_10_io_request_0_valid = b1_25_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_10_io_request_0_bits_time_steps = b1_25_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_10_io_request_0_bits_start_value = b1_25_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_10_io_request_0_bits_coefficient1 = b1_25_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_10_io_request_0_bits_coefficient2 = b1_25_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_10_io_request_1_valid = b2_25_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_10_io_request_1_bits_time_steps = b2_25_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_10_io_request_1_bits_start_value = b2_25_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_10_io_request_1_bits_coefficient1 = b2_25_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_10_io_request_1_bits_coefficient2 = b2_25_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_10_io_response_0_ready = partial_result_impl_io_lanes_20_ready; // @[MonteCarlo.scala 216:19]
  assign engines_10_io_response_1_ready = partial_result_impl_io_lanes_21_ready; // @[MonteCarlo.scala 216:19]
  assign engines_11_clock = clock;
  assign engines_11_reset = reset;
  assign engines_11_io_request_0_valid = b1_26_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_11_io_request_0_bits_time_steps = b1_26_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_11_io_request_0_bits_start_value = b1_26_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_11_io_request_0_bits_coefficient1 = b1_26_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_11_io_request_0_bits_coefficient2 = b1_26_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_11_io_request_1_valid = b2_26_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_11_io_request_1_bits_time_steps = b2_26_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_11_io_request_1_bits_start_value = b2_26_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_11_io_request_1_bits_coefficient1 = b2_26_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_11_io_request_1_bits_coefficient2 = b2_26_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_11_io_response_0_ready = partial_result_impl_io_lanes_22_ready; // @[MonteCarlo.scala 216:19]
  assign engines_11_io_response_1_ready = partial_result_impl_io_lanes_23_ready; // @[MonteCarlo.scala 216:19]
  assign engines_12_clock = clock;
  assign engines_12_reset = reset;
  assign engines_12_io_request_0_valid = b1_27_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_12_io_request_0_bits_time_steps = b1_27_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_12_io_request_0_bits_start_value = b1_27_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_12_io_request_0_bits_coefficient1 = b1_27_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_12_io_request_0_bits_coefficient2 = b1_27_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_12_io_request_1_valid = b2_27_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_12_io_request_1_bits_time_steps = b2_27_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_12_io_request_1_bits_start_value = b2_27_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_12_io_request_1_bits_coefficient1 = b2_27_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_12_io_request_1_bits_coefficient2 = b2_27_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_12_io_response_0_ready = partial_result_impl_io_lanes_24_ready; // @[MonteCarlo.scala 216:19]
  assign engines_12_io_response_1_ready = partial_result_impl_io_lanes_25_ready; // @[MonteCarlo.scala 216:19]
  assign engines_13_clock = clock;
  assign engines_13_reset = reset;
  assign engines_13_io_request_0_valid = b1_28_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_13_io_request_0_bits_time_steps = b1_28_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_13_io_request_0_bits_start_value = b1_28_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_13_io_request_0_bits_coefficient1 = b1_28_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_13_io_request_0_bits_coefficient2 = b1_28_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_13_io_request_1_valid = b2_28_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_13_io_request_1_bits_time_steps = b2_28_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_13_io_request_1_bits_start_value = b2_28_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_13_io_request_1_bits_coefficient1 = b2_28_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_13_io_request_1_bits_coefficient2 = b2_28_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_13_io_response_0_ready = partial_result_impl_io_lanes_26_ready; // @[MonteCarlo.scala 216:19]
  assign engines_13_io_response_1_ready = partial_result_impl_io_lanes_27_ready; // @[MonteCarlo.scala 216:19]
  assign engines_14_clock = clock;
  assign engines_14_reset = reset;
  assign engines_14_io_request_0_valid = b1_29_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_14_io_request_0_bits_time_steps = b1_29_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_14_io_request_0_bits_start_value = b1_29_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_14_io_request_0_bits_coefficient1 = b1_29_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_14_io_request_0_bits_coefficient2 = b1_29_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_14_io_request_1_valid = b2_29_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_14_io_request_1_bits_time_steps = b2_29_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_14_io_request_1_bits_start_value = b2_29_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_14_io_request_1_bits_coefficient1 = b2_29_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_14_io_request_1_bits_coefficient2 = b2_29_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_14_io_response_0_ready = partial_result_impl_io_lanes_28_ready; // @[MonteCarlo.scala 216:19]
  assign engines_14_io_response_1_ready = partial_result_impl_io_lanes_29_ready; // @[MonteCarlo.scala 216:19]
  assign engines_15_clock = clock;
  assign engines_15_reset = reset;
  assign engines_15_io_request_0_valid = b1_30_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_15_io_request_0_bits_time_steps = b1_30_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_15_io_request_0_bits_start_value = b1_30_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_15_io_request_0_bits_coefficient1 = b1_30_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_15_io_request_0_bits_coefficient2 = b1_30_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_15_io_request_1_valid = b2_30_io_deq_valid; // @[MonteCarlo.scala 255:97]
  assign engines_15_io_request_1_bits_time_steps = b2_30_io_deq_bits_time_steps; // @[MonteCarlo.scala 255:97]
  assign engines_15_io_request_1_bits_start_value = b2_30_io_deq_bits_start_value; // @[MonteCarlo.scala 255:97]
  assign engines_15_io_request_1_bits_coefficient1 = b2_30_io_deq_bits_coefficient1; // @[MonteCarlo.scala 255:97]
  assign engines_15_io_request_1_bits_coefficient2 = b2_30_io_deq_bits_coefficient2; // @[MonteCarlo.scala 255:97]
  assign engines_15_io_response_0_ready = partial_result_impl_io_lanes_30_ready; // @[MonteCarlo.scala 216:19]
  assign engines_15_io_response_1_ready = partial_result_impl_io_lanes_31_ready; // @[MonteCarlo.scala 216:19]
  assign b1_clock = clock;
  assign b1_reset = reset;
  assign b1_io_enq_valid = b1_io_enq_ready & io_request_valid; // @[MonteCarlo.scala 241:56]
  assign b1_io_enq_bits_time_steps = io_request_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_io_enq_bits_start_value = io_request_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_io_enq_bits_coefficient1 = io_request_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_io_enq_bits_coefficient2 = io_request_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_io_deq_ready = b1_1_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b2_clock = clock;
  assign b2_reset = reset;
  assign b2_io_enq_valid = b1_io_enq_ready & io_request_valid; // @[MonteCarlo.scala 241:56]
  assign b2_io_enq_bits_time_steps = io_request_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_io_enq_bits_start_value = io_request_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_io_enq_bits_coefficient1 = io_request_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_io_enq_bits_coefficient2 = io_request_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_io_deq_ready = b1_2_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b1_1_clock = clock;
  assign b1_1_reset = reset;
  assign b1_1_io_enq_valid = b1_1_io_enq_ready & b1_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_1_io_enq_bits_time_steps = b1_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_1_io_enq_bits_start_value = b1_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_1_io_enq_bits_coefficient1 = b1_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_1_io_enq_bits_coefficient2 = b1_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_1_io_deq_ready = b1_3_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b2_1_clock = clock;
  assign b2_1_reset = reset;
  assign b2_1_io_enq_valid = b1_1_io_enq_ready & b1_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_1_io_enq_bits_time_steps = b1_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_1_io_enq_bits_start_value = b1_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_1_io_enq_bits_coefficient1 = b1_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_1_io_enq_bits_coefficient2 = b1_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_1_io_deq_ready = b1_4_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b1_2_clock = clock;
  assign b1_2_reset = reset;
  assign b1_2_io_enq_valid = b1_2_io_enq_ready & b2_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_2_io_enq_bits_time_steps = b2_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_2_io_enq_bits_start_value = b2_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_2_io_enq_bits_coefficient1 = b2_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_2_io_enq_bits_coefficient2 = b2_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_2_io_deq_ready = b1_5_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b2_2_clock = clock;
  assign b2_2_reset = reset;
  assign b2_2_io_enq_valid = b1_2_io_enq_ready & b2_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_2_io_enq_bits_time_steps = b2_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_2_io_enq_bits_start_value = b2_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_2_io_enq_bits_coefficient1 = b2_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_2_io_enq_bits_coefficient2 = b2_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_2_io_deq_ready = b1_6_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b1_3_clock = clock;
  assign b1_3_reset = reset;
  assign b1_3_io_enq_valid = b1_3_io_enq_ready & b1_1_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_3_io_enq_bits_time_steps = b1_1_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_3_io_enq_bits_start_value = b1_1_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_3_io_enq_bits_coefficient1 = b1_1_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_3_io_enq_bits_coefficient2 = b1_1_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_3_io_deq_ready = b1_7_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b2_3_clock = clock;
  assign b2_3_reset = reset;
  assign b2_3_io_enq_valid = b1_3_io_enq_ready & b1_1_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_3_io_enq_bits_time_steps = b1_1_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_3_io_enq_bits_start_value = b1_1_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_3_io_enq_bits_coefficient1 = b1_1_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_3_io_enq_bits_coefficient2 = b1_1_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_3_io_deq_ready = b1_8_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b1_4_clock = clock;
  assign b1_4_reset = reset;
  assign b1_4_io_enq_valid = b1_4_io_enq_ready & b2_1_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_4_io_enq_bits_time_steps = b2_1_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_4_io_enq_bits_start_value = b2_1_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_4_io_enq_bits_coefficient1 = b2_1_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_4_io_enq_bits_coefficient2 = b2_1_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_4_io_deq_ready = b1_9_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b2_4_clock = clock;
  assign b2_4_reset = reset;
  assign b2_4_io_enq_valid = b1_4_io_enq_ready & b2_1_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_4_io_enq_bits_time_steps = b2_1_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_4_io_enq_bits_start_value = b2_1_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_4_io_enq_bits_coefficient1 = b2_1_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_4_io_enq_bits_coefficient2 = b2_1_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_4_io_deq_ready = b1_10_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b1_5_clock = clock;
  assign b1_5_reset = reset;
  assign b1_5_io_enq_valid = b1_5_io_enq_ready & b1_2_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_5_io_enq_bits_time_steps = b1_2_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_5_io_enq_bits_start_value = b1_2_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_5_io_enq_bits_coefficient1 = b1_2_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_5_io_enq_bits_coefficient2 = b1_2_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_5_io_deq_ready = b1_11_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b2_5_clock = clock;
  assign b2_5_reset = reset;
  assign b2_5_io_enq_valid = b1_5_io_enq_ready & b1_2_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_5_io_enq_bits_time_steps = b1_2_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_5_io_enq_bits_start_value = b1_2_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_5_io_enq_bits_coefficient1 = b1_2_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_5_io_enq_bits_coefficient2 = b1_2_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_5_io_deq_ready = b1_12_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b1_6_clock = clock;
  assign b1_6_reset = reset;
  assign b1_6_io_enq_valid = b1_6_io_enq_ready & b2_2_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_6_io_enq_bits_time_steps = b2_2_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_6_io_enq_bits_start_value = b2_2_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_6_io_enq_bits_coefficient1 = b2_2_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_6_io_enq_bits_coefficient2 = b2_2_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_6_io_deq_ready = b1_13_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b2_6_clock = clock;
  assign b2_6_reset = reset;
  assign b2_6_io_enq_valid = b1_6_io_enq_ready & b2_2_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_6_io_enq_bits_time_steps = b2_2_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_6_io_enq_bits_start_value = b2_2_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_6_io_enq_bits_coefficient1 = b2_2_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_6_io_enq_bits_coefficient2 = b2_2_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_6_io_deq_ready = b1_14_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b1_7_clock = clock;
  assign b1_7_reset = reset;
  assign b1_7_io_enq_valid = b1_7_io_enq_ready & b1_3_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_7_io_enq_bits_time_steps = b1_3_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_7_io_enq_bits_start_value = b1_3_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_7_io_enq_bits_coefficient1 = b1_3_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_7_io_enq_bits_coefficient2 = b1_3_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_7_io_deq_ready = b1_15_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b2_7_clock = clock;
  assign b2_7_reset = reset;
  assign b2_7_io_enq_valid = b1_7_io_enq_ready & b1_3_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_7_io_enq_bits_time_steps = b1_3_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_7_io_enq_bits_start_value = b1_3_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_7_io_enq_bits_coefficient1 = b1_3_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_7_io_enq_bits_coefficient2 = b1_3_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_7_io_deq_ready = b1_16_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b1_8_clock = clock;
  assign b1_8_reset = reset;
  assign b1_8_io_enq_valid = b1_8_io_enq_ready & b2_3_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_8_io_enq_bits_time_steps = b2_3_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_8_io_enq_bits_start_value = b2_3_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_8_io_enq_bits_coefficient1 = b2_3_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_8_io_enq_bits_coefficient2 = b2_3_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_8_io_deq_ready = b1_17_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b2_8_clock = clock;
  assign b2_8_reset = reset;
  assign b2_8_io_enq_valid = b1_8_io_enq_ready & b2_3_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_8_io_enq_bits_time_steps = b2_3_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_8_io_enq_bits_start_value = b2_3_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_8_io_enq_bits_coefficient1 = b2_3_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_8_io_enq_bits_coefficient2 = b2_3_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_8_io_deq_ready = b1_18_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b1_9_clock = clock;
  assign b1_9_reset = reset;
  assign b1_9_io_enq_valid = b1_9_io_enq_ready & b1_4_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_9_io_enq_bits_time_steps = b1_4_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_9_io_enq_bits_start_value = b1_4_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_9_io_enq_bits_coefficient1 = b1_4_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_9_io_enq_bits_coefficient2 = b1_4_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_9_io_deq_ready = b1_19_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b2_9_clock = clock;
  assign b2_9_reset = reset;
  assign b2_9_io_enq_valid = b1_9_io_enq_ready & b1_4_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_9_io_enq_bits_time_steps = b1_4_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_9_io_enq_bits_start_value = b1_4_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_9_io_enq_bits_coefficient1 = b1_4_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_9_io_enq_bits_coefficient2 = b1_4_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_9_io_deq_ready = b1_20_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b1_10_clock = clock;
  assign b1_10_reset = reset;
  assign b1_10_io_enq_valid = b1_10_io_enq_ready & b2_4_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_10_io_enq_bits_time_steps = b2_4_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_10_io_enq_bits_start_value = b2_4_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_10_io_enq_bits_coefficient1 = b2_4_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_10_io_enq_bits_coefficient2 = b2_4_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_10_io_deq_ready = b1_21_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b2_10_clock = clock;
  assign b2_10_reset = reset;
  assign b2_10_io_enq_valid = b1_10_io_enq_ready & b2_4_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_10_io_enq_bits_time_steps = b2_4_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_10_io_enq_bits_start_value = b2_4_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_10_io_enq_bits_coefficient1 = b2_4_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_10_io_enq_bits_coefficient2 = b2_4_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_10_io_deq_ready = b1_22_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b1_11_clock = clock;
  assign b1_11_reset = reset;
  assign b1_11_io_enq_valid = b1_11_io_enq_ready & b1_5_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_11_io_enq_bits_time_steps = b1_5_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_11_io_enq_bits_start_value = b1_5_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_11_io_enq_bits_coefficient1 = b1_5_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_11_io_enq_bits_coefficient2 = b1_5_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_11_io_deq_ready = b1_23_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b2_11_clock = clock;
  assign b2_11_reset = reset;
  assign b2_11_io_enq_valid = b1_11_io_enq_ready & b1_5_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_11_io_enq_bits_time_steps = b1_5_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_11_io_enq_bits_start_value = b1_5_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_11_io_enq_bits_coefficient1 = b1_5_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_11_io_enq_bits_coefficient2 = b1_5_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_11_io_deq_ready = b1_24_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b1_12_clock = clock;
  assign b1_12_reset = reset;
  assign b1_12_io_enq_valid = b1_12_io_enq_ready & b2_5_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_12_io_enq_bits_time_steps = b2_5_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_12_io_enq_bits_start_value = b2_5_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_12_io_enq_bits_coefficient1 = b2_5_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_12_io_enq_bits_coefficient2 = b2_5_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_12_io_deq_ready = b1_25_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b2_12_clock = clock;
  assign b2_12_reset = reset;
  assign b2_12_io_enq_valid = b1_12_io_enq_ready & b2_5_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_12_io_enq_bits_time_steps = b2_5_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_12_io_enq_bits_start_value = b2_5_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_12_io_enq_bits_coefficient1 = b2_5_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_12_io_enq_bits_coefficient2 = b2_5_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_12_io_deq_ready = b1_26_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b1_13_clock = clock;
  assign b1_13_reset = reset;
  assign b1_13_io_enq_valid = b1_13_io_enq_ready & b1_6_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_13_io_enq_bits_time_steps = b1_6_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_13_io_enq_bits_start_value = b1_6_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_13_io_enq_bits_coefficient1 = b1_6_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_13_io_enq_bits_coefficient2 = b1_6_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_13_io_deq_ready = b1_27_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b2_13_clock = clock;
  assign b2_13_reset = reset;
  assign b2_13_io_enq_valid = b1_13_io_enq_ready & b1_6_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_13_io_enq_bits_time_steps = b1_6_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_13_io_enq_bits_start_value = b1_6_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_13_io_enq_bits_coefficient1 = b1_6_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_13_io_enq_bits_coefficient2 = b1_6_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_13_io_deq_ready = b1_28_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b1_14_clock = clock;
  assign b1_14_reset = reset;
  assign b1_14_io_enq_valid = b1_14_io_enq_ready & b2_6_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_14_io_enq_bits_time_steps = b2_6_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_14_io_enq_bits_start_value = b2_6_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_14_io_enq_bits_coefficient1 = b2_6_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_14_io_enq_bits_coefficient2 = b2_6_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_14_io_deq_ready = b1_29_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b2_14_clock = clock;
  assign b2_14_reset = reset;
  assign b2_14_io_enq_valid = b1_14_io_enq_ready & b2_6_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_14_io_enq_bits_time_steps = b2_6_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_14_io_enq_bits_start_value = b2_6_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_14_io_enq_bits_coefficient1 = b2_6_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_14_io_enq_bits_coefficient2 = b2_6_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_14_io_deq_ready = b1_30_io_enq_ready; // @[MonteCarlo.scala 242:46]
  assign b1_15_clock = clock;
  assign b1_15_reset = reset;
  assign b1_15_io_enq_valid = b1_15_io_enq_ready & b1_7_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_15_io_enq_bits_time_steps = b1_7_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_15_io_enq_bits_start_value = b1_7_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_15_io_enq_bits_coefficient1 = b1_7_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_15_io_enq_bits_coefficient2 = b1_7_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_15_io_deq_ready = engines_0_io_request_0_ready; // @[MonteCarlo.scala 255:97]
  assign b2_15_clock = clock;
  assign b2_15_reset = reset;
  assign b2_15_io_enq_valid = b1_15_io_enq_ready & b1_7_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_15_io_enq_bits_time_steps = b1_7_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_15_io_enq_bits_start_value = b1_7_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_15_io_enq_bits_coefficient1 = b1_7_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_15_io_enq_bits_coefficient2 = b1_7_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_15_io_deq_ready = engines_0_io_request_1_ready; // @[MonteCarlo.scala 255:97]
  assign b1_16_clock = clock;
  assign b1_16_reset = reset;
  assign b1_16_io_enq_valid = b1_16_io_enq_ready & b2_7_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_16_io_enq_bits_time_steps = b2_7_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_16_io_enq_bits_start_value = b2_7_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_16_io_enq_bits_coefficient1 = b2_7_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_16_io_enq_bits_coefficient2 = b2_7_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_16_io_deq_ready = engines_1_io_request_0_ready; // @[MonteCarlo.scala 255:97]
  assign b2_16_clock = clock;
  assign b2_16_reset = reset;
  assign b2_16_io_enq_valid = b1_16_io_enq_ready & b2_7_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_16_io_enq_bits_time_steps = b2_7_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_16_io_enq_bits_start_value = b2_7_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_16_io_enq_bits_coefficient1 = b2_7_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_16_io_enq_bits_coefficient2 = b2_7_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_16_io_deq_ready = engines_1_io_request_1_ready; // @[MonteCarlo.scala 255:97]
  assign b1_17_clock = clock;
  assign b1_17_reset = reset;
  assign b1_17_io_enq_valid = b1_17_io_enq_ready & b1_8_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_17_io_enq_bits_time_steps = b1_8_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_17_io_enq_bits_start_value = b1_8_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_17_io_enq_bits_coefficient1 = b1_8_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_17_io_enq_bits_coefficient2 = b1_8_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_17_io_deq_ready = engines_2_io_request_0_ready; // @[MonteCarlo.scala 255:97]
  assign b2_17_clock = clock;
  assign b2_17_reset = reset;
  assign b2_17_io_enq_valid = b1_17_io_enq_ready & b1_8_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_17_io_enq_bits_time_steps = b1_8_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_17_io_enq_bits_start_value = b1_8_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_17_io_enq_bits_coefficient1 = b1_8_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_17_io_enq_bits_coefficient2 = b1_8_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_17_io_deq_ready = engines_2_io_request_1_ready; // @[MonteCarlo.scala 255:97]
  assign b1_18_clock = clock;
  assign b1_18_reset = reset;
  assign b1_18_io_enq_valid = b1_18_io_enq_ready & b2_8_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_18_io_enq_bits_time_steps = b2_8_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_18_io_enq_bits_start_value = b2_8_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_18_io_enq_bits_coefficient1 = b2_8_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_18_io_enq_bits_coefficient2 = b2_8_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_18_io_deq_ready = engines_3_io_request_0_ready; // @[MonteCarlo.scala 255:97]
  assign b2_18_clock = clock;
  assign b2_18_reset = reset;
  assign b2_18_io_enq_valid = b1_18_io_enq_ready & b2_8_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_18_io_enq_bits_time_steps = b2_8_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_18_io_enq_bits_start_value = b2_8_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_18_io_enq_bits_coefficient1 = b2_8_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_18_io_enq_bits_coefficient2 = b2_8_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_18_io_deq_ready = engines_3_io_request_1_ready; // @[MonteCarlo.scala 255:97]
  assign b1_19_clock = clock;
  assign b1_19_reset = reset;
  assign b1_19_io_enq_valid = b1_19_io_enq_ready & b1_9_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_19_io_enq_bits_time_steps = b1_9_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_19_io_enq_bits_start_value = b1_9_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_19_io_enq_bits_coefficient1 = b1_9_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_19_io_enq_bits_coefficient2 = b1_9_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_19_io_deq_ready = engines_4_io_request_0_ready; // @[MonteCarlo.scala 255:97]
  assign b2_19_clock = clock;
  assign b2_19_reset = reset;
  assign b2_19_io_enq_valid = b1_19_io_enq_ready & b1_9_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_19_io_enq_bits_time_steps = b1_9_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_19_io_enq_bits_start_value = b1_9_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_19_io_enq_bits_coefficient1 = b1_9_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_19_io_enq_bits_coefficient2 = b1_9_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_19_io_deq_ready = engines_4_io_request_1_ready; // @[MonteCarlo.scala 255:97]
  assign b1_20_clock = clock;
  assign b1_20_reset = reset;
  assign b1_20_io_enq_valid = b1_20_io_enq_ready & b2_9_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_20_io_enq_bits_time_steps = b2_9_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_20_io_enq_bits_start_value = b2_9_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_20_io_enq_bits_coefficient1 = b2_9_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_20_io_enq_bits_coefficient2 = b2_9_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_20_io_deq_ready = engines_5_io_request_0_ready; // @[MonteCarlo.scala 255:97]
  assign b2_20_clock = clock;
  assign b2_20_reset = reset;
  assign b2_20_io_enq_valid = b1_20_io_enq_ready & b2_9_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_20_io_enq_bits_time_steps = b2_9_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_20_io_enq_bits_start_value = b2_9_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_20_io_enq_bits_coefficient1 = b2_9_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_20_io_enq_bits_coefficient2 = b2_9_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_20_io_deq_ready = engines_5_io_request_1_ready; // @[MonteCarlo.scala 255:97]
  assign b1_21_clock = clock;
  assign b1_21_reset = reset;
  assign b1_21_io_enq_valid = b1_21_io_enq_ready & b1_10_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_21_io_enq_bits_time_steps = b1_10_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_21_io_enq_bits_start_value = b1_10_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_21_io_enq_bits_coefficient1 = b1_10_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_21_io_enq_bits_coefficient2 = b1_10_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_21_io_deq_ready = engines_6_io_request_0_ready; // @[MonteCarlo.scala 255:97]
  assign b2_21_clock = clock;
  assign b2_21_reset = reset;
  assign b2_21_io_enq_valid = b1_21_io_enq_ready & b1_10_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_21_io_enq_bits_time_steps = b1_10_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_21_io_enq_bits_start_value = b1_10_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_21_io_enq_bits_coefficient1 = b1_10_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_21_io_enq_bits_coefficient2 = b1_10_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_21_io_deq_ready = engines_6_io_request_1_ready; // @[MonteCarlo.scala 255:97]
  assign b1_22_clock = clock;
  assign b1_22_reset = reset;
  assign b1_22_io_enq_valid = b1_22_io_enq_ready & b2_10_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_22_io_enq_bits_time_steps = b2_10_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_22_io_enq_bits_start_value = b2_10_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_22_io_enq_bits_coefficient1 = b2_10_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_22_io_enq_bits_coefficient2 = b2_10_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_22_io_deq_ready = engines_7_io_request_0_ready; // @[MonteCarlo.scala 255:97]
  assign b2_22_clock = clock;
  assign b2_22_reset = reset;
  assign b2_22_io_enq_valid = b1_22_io_enq_ready & b2_10_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_22_io_enq_bits_time_steps = b2_10_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_22_io_enq_bits_start_value = b2_10_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_22_io_enq_bits_coefficient1 = b2_10_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_22_io_enq_bits_coefficient2 = b2_10_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_22_io_deq_ready = engines_7_io_request_1_ready; // @[MonteCarlo.scala 255:97]
  assign b1_23_clock = clock;
  assign b1_23_reset = reset;
  assign b1_23_io_enq_valid = b1_23_io_enq_ready & b1_11_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_23_io_enq_bits_time_steps = b1_11_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_23_io_enq_bits_start_value = b1_11_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_23_io_enq_bits_coefficient1 = b1_11_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_23_io_enq_bits_coefficient2 = b1_11_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_23_io_deq_ready = engines_8_io_request_0_ready; // @[MonteCarlo.scala 255:97]
  assign b2_23_clock = clock;
  assign b2_23_reset = reset;
  assign b2_23_io_enq_valid = b1_23_io_enq_ready & b1_11_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_23_io_enq_bits_time_steps = b1_11_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_23_io_enq_bits_start_value = b1_11_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_23_io_enq_bits_coefficient1 = b1_11_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_23_io_enq_bits_coefficient2 = b1_11_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_23_io_deq_ready = engines_8_io_request_1_ready; // @[MonteCarlo.scala 255:97]
  assign b1_24_clock = clock;
  assign b1_24_reset = reset;
  assign b1_24_io_enq_valid = b1_24_io_enq_ready & b2_11_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_24_io_enq_bits_time_steps = b2_11_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_24_io_enq_bits_start_value = b2_11_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_24_io_enq_bits_coefficient1 = b2_11_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_24_io_enq_bits_coefficient2 = b2_11_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_24_io_deq_ready = engines_9_io_request_0_ready; // @[MonteCarlo.scala 255:97]
  assign b2_24_clock = clock;
  assign b2_24_reset = reset;
  assign b2_24_io_enq_valid = b1_24_io_enq_ready & b2_11_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_24_io_enq_bits_time_steps = b2_11_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_24_io_enq_bits_start_value = b2_11_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_24_io_enq_bits_coefficient1 = b2_11_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_24_io_enq_bits_coefficient2 = b2_11_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_24_io_deq_ready = engines_9_io_request_1_ready; // @[MonteCarlo.scala 255:97]
  assign b1_25_clock = clock;
  assign b1_25_reset = reset;
  assign b1_25_io_enq_valid = b1_25_io_enq_ready & b1_12_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_25_io_enq_bits_time_steps = b1_12_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_25_io_enq_bits_start_value = b1_12_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_25_io_enq_bits_coefficient1 = b1_12_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_25_io_enq_bits_coefficient2 = b1_12_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_25_io_deq_ready = engines_10_io_request_0_ready; // @[MonteCarlo.scala 255:97]
  assign b2_25_clock = clock;
  assign b2_25_reset = reset;
  assign b2_25_io_enq_valid = b1_25_io_enq_ready & b1_12_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_25_io_enq_bits_time_steps = b1_12_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_25_io_enq_bits_start_value = b1_12_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_25_io_enq_bits_coefficient1 = b1_12_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_25_io_enq_bits_coefficient2 = b1_12_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_25_io_deq_ready = engines_10_io_request_1_ready; // @[MonteCarlo.scala 255:97]
  assign b1_26_clock = clock;
  assign b1_26_reset = reset;
  assign b1_26_io_enq_valid = b1_26_io_enq_ready & b2_12_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_26_io_enq_bits_time_steps = b2_12_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_26_io_enq_bits_start_value = b2_12_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_26_io_enq_bits_coefficient1 = b2_12_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_26_io_enq_bits_coefficient2 = b2_12_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_26_io_deq_ready = engines_11_io_request_0_ready; // @[MonteCarlo.scala 255:97]
  assign b2_26_clock = clock;
  assign b2_26_reset = reset;
  assign b2_26_io_enq_valid = b1_26_io_enq_ready & b2_12_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_26_io_enq_bits_time_steps = b2_12_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_26_io_enq_bits_start_value = b2_12_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_26_io_enq_bits_coefficient1 = b2_12_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_26_io_enq_bits_coefficient2 = b2_12_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_26_io_deq_ready = engines_11_io_request_1_ready; // @[MonteCarlo.scala 255:97]
  assign b1_27_clock = clock;
  assign b1_27_reset = reset;
  assign b1_27_io_enq_valid = b1_27_io_enq_ready & b1_13_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_27_io_enq_bits_time_steps = b1_13_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_27_io_enq_bits_start_value = b1_13_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_27_io_enq_bits_coefficient1 = b1_13_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_27_io_enq_bits_coefficient2 = b1_13_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_27_io_deq_ready = engines_12_io_request_0_ready; // @[MonteCarlo.scala 255:97]
  assign b2_27_clock = clock;
  assign b2_27_reset = reset;
  assign b2_27_io_enq_valid = b1_27_io_enq_ready & b1_13_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_27_io_enq_bits_time_steps = b1_13_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_27_io_enq_bits_start_value = b1_13_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_27_io_enq_bits_coefficient1 = b1_13_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_27_io_enq_bits_coefficient2 = b1_13_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_27_io_deq_ready = engines_12_io_request_1_ready; // @[MonteCarlo.scala 255:97]
  assign b1_28_clock = clock;
  assign b1_28_reset = reset;
  assign b1_28_io_enq_valid = b1_28_io_enq_ready & b2_13_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_28_io_enq_bits_time_steps = b2_13_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_28_io_enq_bits_start_value = b2_13_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_28_io_enq_bits_coefficient1 = b2_13_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_28_io_enq_bits_coefficient2 = b2_13_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_28_io_deq_ready = engines_13_io_request_0_ready; // @[MonteCarlo.scala 255:97]
  assign b2_28_clock = clock;
  assign b2_28_reset = reset;
  assign b2_28_io_enq_valid = b1_28_io_enq_ready & b2_13_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_28_io_enq_bits_time_steps = b2_13_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_28_io_enq_bits_start_value = b2_13_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_28_io_enq_bits_coefficient1 = b2_13_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_28_io_enq_bits_coefficient2 = b2_13_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_28_io_deq_ready = engines_13_io_request_1_ready; // @[MonteCarlo.scala 255:97]
  assign b1_29_clock = clock;
  assign b1_29_reset = reset;
  assign b1_29_io_enq_valid = b1_29_io_enq_ready & b1_14_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_29_io_enq_bits_time_steps = b1_14_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_29_io_enq_bits_start_value = b1_14_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_29_io_enq_bits_coefficient1 = b1_14_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_29_io_enq_bits_coefficient2 = b1_14_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_29_io_deq_ready = engines_14_io_request_0_ready; // @[MonteCarlo.scala 255:97]
  assign b2_29_clock = clock;
  assign b2_29_reset = reset;
  assign b2_29_io_enq_valid = b1_29_io_enq_ready & b1_14_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_29_io_enq_bits_time_steps = b1_14_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_29_io_enq_bits_start_value = b1_14_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_29_io_enq_bits_coefficient1 = b1_14_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_29_io_enq_bits_coefficient2 = b1_14_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_29_io_deq_ready = engines_14_io_request_1_ready; // @[MonteCarlo.scala 255:97]
  assign b1_30_clock = clock;
  assign b1_30_reset = reset;
  assign b1_30_io_enq_valid = b1_30_io_enq_ready & b2_14_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b1_30_io_enq_bits_time_steps = b2_14_io_deq_bits_time_steps; // @[MonteCarlo.scala 243:27]
  assign b1_30_io_enq_bits_start_value = b2_14_io_deq_bits_start_value; // @[MonteCarlo.scala 243:27]
  assign b1_30_io_enq_bits_coefficient1 = b2_14_io_deq_bits_coefficient1; // @[MonteCarlo.scala 243:27]
  assign b1_30_io_enq_bits_coefficient2 = b2_14_io_deq_bits_coefficient2; // @[MonteCarlo.scala 243:27]
  assign b1_30_io_deq_ready = engines_15_io_request_0_ready; // @[MonteCarlo.scala 255:97]
  assign b2_30_clock = clock;
  assign b2_30_reset = reset;
  assign b2_30_io_enq_valid = b1_30_io_enq_ready & b2_14_io_deq_valid; // @[MonteCarlo.scala 241:56]
  assign b2_30_io_enq_bits_time_steps = b2_14_io_deq_bits_time_steps; // @[MonteCarlo.scala 244:27]
  assign b2_30_io_enq_bits_start_value = b2_14_io_deq_bits_start_value; // @[MonteCarlo.scala 244:27]
  assign b2_30_io_enq_bits_coefficient1 = b2_14_io_deq_bits_coefficient1; // @[MonteCarlo.scala 244:27]
  assign b2_30_io_enq_bits_coefficient2 = b2_14_io_deq_bits_coefficient2; // @[MonteCarlo.scala 244:27]
  assign b2_30_io_deq_ready = engines_15_io_request_1_ready; // @[MonteCarlo.scala 255:97]
  assign partial_result_impl_clock = clock;
  assign partial_result_impl_reset = reset;
  assign partial_result_impl_io_lanes_0_valid = engines_0_io_response_0_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_0_bits = engines_0_io_response_0_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_1_valid = engines_0_io_response_1_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_1_bits = engines_0_io_response_1_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_2_valid = engines_1_io_response_0_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_2_bits = engines_1_io_response_0_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_3_valid = engines_1_io_response_1_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_3_bits = engines_1_io_response_1_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_4_valid = engines_2_io_response_0_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_4_bits = engines_2_io_response_0_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_5_valid = engines_2_io_response_1_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_5_bits = engines_2_io_response_1_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_6_valid = engines_3_io_response_0_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_6_bits = engines_3_io_response_0_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_7_valid = engines_3_io_response_1_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_7_bits = engines_3_io_response_1_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_8_valid = engines_4_io_response_0_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_8_bits = engines_4_io_response_0_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_9_valid = engines_4_io_response_1_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_9_bits = engines_4_io_response_1_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_10_valid = engines_5_io_response_0_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_10_bits = engines_5_io_response_0_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_11_valid = engines_5_io_response_1_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_11_bits = engines_5_io_response_1_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_12_valid = engines_6_io_response_0_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_12_bits = engines_6_io_response_0_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_13_valid = engines_6_io_response_1_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_13_bits = engines_6_io_response_1_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_14_valid = engines_7_io_response_0_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_14_bits = engines_7_io_response_0_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_15_valid = engines_7_io_response_1_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_15_bits = engines_7_io_response_1_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_16_valid = engines_8_io_response_0_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_16_bits = engines_8_io_response_0_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_17_valid = engines_8_io_response_1_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_17_bits = engines_8_io_response_1_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_18_valid = engines_9_io_response_0_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_18_bits = engines_9_io_response_0_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_19_valid = engines_9_io_response_1_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_19_bits = engines_9_io_response_1_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_20_valid = engines_10_io_response_0_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_20_bits = engines_10_io_response_0_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_21_valid = engines_10_io_response_1_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_21_bits = engines_10_io_response_1_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_22_valid = engines_11_io_response_0_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_22_bits = engines_11_io_response_0_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_23_valid = engines_11_io_response_1_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_23_bits = engines_11_io_response_1_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_24_valid = engines_12_io_response_0_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_24_bits = engines_12_io_response_0_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_25_valid = engines_12_io_response_1_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_25_bits = engines_12_io_response_1_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_26_valid = engines_13_io_response_0_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_26_bits = engines_13_io_response_0_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_27_valid = engines_13_io_response_1_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_27_bits = engines_13_io_response_1_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_28_valid = engines_14_io_response_0_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_28_bits = engines_14_io_response_0_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_29_valid = engines_14_io_response_1_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_29_bits = engines_14_io_response_1_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_30_valid = engines_15_io_response_0_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_30_bits = engines_15_io_response_0_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_31_valid = engines_15_io_response_1_valid; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_lanes_31_bits = engines_15_io_response_1_bits; // @[MonteCarlo.scala 216:19]
  assign partial_result_impl_io_result_ready = io_response_ready; // @[MonteCarlo.scala 259:15]
endmodule
