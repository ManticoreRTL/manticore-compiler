module VCR(
  input         clock,
  input         reset,
  output        io_host_aw_ready,
  input         io_host_aw_valid,
  input  [15:0] io_host_aw_bits_addr,
  output        io_host_w_ready,
  input         io_host_w_valid,
  input  [31:0] io_host_w_bits_data,
  input         io_host_b_ready,
  output        io_host_b_valid,
  output        io_host_ar_ready,
  input         io_host_ar_valid,
  input  [15:0] io_host_ar_bits_addr,
  input         io_host_r_ready,
  output        io_host_r_valid,
  output [31:0] io_host_r_bits_data,
  output        io_vcr_launch,
  input         io_vcr_finish,
  input         io_vcr_ecnt_0_valid,
  input  [31:0] io_vcr_ecnt_0_bits,
  output [31:0] io_vcr_vals_0,
  output [31:0] io_vcr_ptrs_0,
  output [31:0] io_vcr_ptrs_1,
  output [31:0] io_vcr_ptrs_2,
  output [31:0] io_vcr_ptrs_3,
  output [31:0] io_vcr_ptrs_4,
  output [31:0] io_vcr_ptrs_5,
  input         io_vcr_ucnt_0_valid,
  input  [31:0] io_vcr_ucnt_0_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] waddr; // @[VCR.scala 94:22]
  reg [1:0] wstate; // @[VCR.scala 97:23]
  reg  rstate; // @[VCR.scala 101:23]
  reg [31:0] rdata; // @[VCR.scala 102:22]
  reg [31:0] reg_0; // @[VCR.scala 108:37]
  reg [31:0] reg_1; // @[VCR.scala 108:37]
  reg [31:0] reg_2; // @[VCR.scala 108:37]
  reg [31:0] reg_3; // @[VCR.scala 108:37]
  reg [31:0] reg_4; // @[VCR.scala 108:37]
  reg [31:0] reg_5; // @[VCR.scala 108:37]
  reg [31:0] reg_6; // @[VCR.scala 108:37]
  reg [31:0] reg_7; // @[VCR.scala 108:37]
  reg [31:0] reg_8; // @[VCR.scala 108:37]
  reg [31:0] reg_9; // @[VCR.scala 108:37]
  wire [1:0] _GEN_2 = io_host_b_ready ? 2'h0 : wstate; // @[VCR.scala 128:29 129:16 97:23]
  wire  _T_3 = io_host_aw_ready & io_host_aw_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_7 = io_host_ar_valid | rstate; // @[VCR.scala 143:30 144:16 101:23]
  wire  _T_6 = io_host_w_ready & io_host_w_valid; // @[Decoupled.scala 50:35]
  wire  _T_33 = io_host_ar_ready & io_host_ar_valid; // @[Decoupled.scala 50:35]
  wire [31:0] _rdata_T_1 = 16'h0 == io_host_ar_bits_addr ? reg_0 : 32'h0; // @[Mux.scala 81:58]
  wire [31:0] _rdata_T_3 = 16'h4 == io_host_ar_bits_addr ? reg_1 : _rdata_T_1; // @[Mux.scala 81:58]
  wire [31:0] _rdata_T_5 = 16'h8 == io_host_ar_bits_addr ? reg_2 : _rdata_T_3; // @[Mux.scala 81:58]
  wire [31:0] _rdata_T_7 = 16'hc == io_host_ar_bits_addr ? reg_3 : _rdata_T_5; // @[Mux.scala 81:58]
  wire [31:0] _rdata_T_9 = 16'h10 == io_host_ar_bits_addr ? reg_4 : _rdata_T_7; // @[Mux.scala 81:58]
  wire [31:0] _rdata_T_11 = 16'h14 == io_host_ar_bits_addr ? reg_5 : _rdata_T_9; // @[Mux.scala 81:58]
  wire [31:0] _rdata_T_13 = 16'h18 == io_host_ar_bits_addr ? reg_6 : _rdata_T_11; // @[Mux.scala 81:58]
  wire [31:0] _rdata_T_15 = 16'h1c == io_host_ar_bits_addr ? reg_7 : _rdata_T_13; // @[Mux.scala 81:58]
  assign io_host_aw_ready = wstate == 2'h0; // @[VCR.scala 136:30]
  assign io_host_w_ready = wstate == 2'h1; // @[VCR.scala 137:29]
  assign io_host_b_valid = wstate == 2'h2; // @[VCR.scala 138:29]
  assign io_host_ar_ready = ~rstate; // @[VCR.scala 154:30]
  assign io_host_r_valid = rstate; // @[VCR.scala 155:29]
  assign io_host_r_bits_data = rdata; // @[VCR.scala 156:23]
  assign io_vcr_launch = reg_0[0]; // @[VCR.scala 183:26]
  assign io_vcr_vals_0 = reg_2; // @[VCR.scala 186:20]
  assign io_vcr_ptrs_0 = reg_3; // @[VCR.scala 191:22]
  assign io_vcr_ptrs_1 = reg_4; // @[VCR.scala 191:22]
  assign io_vcr_ptrs_2 = reg_5; // @[VCR.scala 191:22]
  assign io_vcr_ptrs_3 = reg_6; // @[VCR.scala 191:22]
  assign io_vcr_ptrs_4 = reg_7; // @[VCR.scala 191:22]
  assign io_vcr_ptrs_5 = reg_8; // @[VCR.scala 191:22]
  always @(posedge clock) begin
    if (reset) begin // @[VCR.scala 94:22]
      waddr <= 16'hffff; // @[VCR.scala 94:22]
    end else if (_T_3) begin // @[VCR.scala 134:25]
      waddr <= io_host_aw_bits_addr; // @[VCR.scala 134:33]
    end
    if (reset) begin // @[VCR.scala 97:23]
      wstate <= 2'h0; // @[VCR.scala 97:23]
    end else if (2'h0 == wstate) begin // @[VCR.scala 116:18]
      if (io_host_aw_valid) begin // @[VCR.scala 118:30]
        wstate <= 2'h1; // @[VCR.scala 119:16]
      end
    end else if (2'h1 == wstate) begin // @[VCR.scala 116:18]
      if (io_host_w_valid) begin // @[VCR.scala 123:29]
        wstate <= 2'h2; // @[VCR.scala 124:16]
      end
    end else if (2'h2 == wstate) begin // @[VCR.scala 116:18]
      wstate <= _GEN_2;
    end
    if (reset) begin // @[VCR.scala 101:23]
      rstate <= 1'h0; // @[VCR.scala 101:23]
    end else if (~rstate) begin // @[VCR.scala 141:18]
      rstate <= _GEN_7;
    end else if (rstate) begin // @[VCR.scala 141:18]
      if (io_host_r_ready) begin // @[VCR.scala 148:29]
        rstate <= 1'h0; // @[VCR.scala 149:16]
      end
    end
    if (reset) begin // @[VCR.scala 102:22]
      rdata <= 32'h0; // @[VCR.scala 102:22]
    end else if (_T_33) begin // @[VCR.scala 179:25]
      if (16'h24 == io_host_ar_bits_addr) begin // @[Mux.scala 81:58]
        rdata <= reg_9;
      end else if (16'h20 == io_host_ar_bits_addr) begin // @[Mux.scala 81:58]
        rdata <= reg_8;
      end else begin
        rdata <= _rdata_T_15;
      end
    end
    if (reset) begin // @[VCR.scala 108:37]
      reg_0 <= 32'h0; // @[VCR.scala 108:37]
    end else if (io_vcr_finish) begin // @[VCR.scala 159:23]
      reg_0 <= 32'h2; // @[VCR.scala 160:12]
    end else if (_T_6 & 16'h0 == waddr) begin // @[VCR.scala 161:53]
      reg_0 <= io_host_w_bits_data; // @[VCR.scala 162:12]
    end
    if (reset) begin // @[VCR.scala 108:37]
      reg_1 <= 32'h0; // @[VCR.scala 108:37]
    end else if (io_vcr_ecnt_0_valid) begin // @[VCR.scala 166:32]
      reg_1 <= io_vcr_ecnt_0_bits; // @[VCR.scala 167:19]
    end else if (_T_6 & 16'h4 == waddr) begin // @[VCR.scala 168:60]
      reg_1 <= io_host_w_bits_data; // @[VCR.scala 169:19]
    end
    if (reset) begin // @[VCR.scala 108:37]
      reg_2 <= 32'h0; // @[VCR.scala 108:37]
    end else if (_T_6 & 16'h8 == waddr) begin // @[VCR.scala 174:54]
      reg_2 <= io_host_w_bits_data; // @[VCR.scala 175:19]
    end
    if (reset) begin // @[VCR.scala 108:37]
      reg_3 <= 32'h0; // @[VCR.scala 108:37]
    end else if (_T_6 & 16'hc == waddr) begin // @[VCR.scala 174:54]
      reg_3 <= io_host_w_bits_data; // @[VCR.scala 175:19]
    end
    if (reset) begin // @[VCR.scala 108:37]
      reg_4 <= 32'h0; // @[VCR.scala 108:37]
    end else if (_T_6 & 16'h10 == waddr) begin // @[VCR.scala 174:54]
      reg_4 <= io_host_w_bits_data; // @[VCR.scala 175:19]
    end
    if (reset) begin // @[VCR.scala 108:37]
      reg_5 <= 32'h0; // @[VCR.scala 108:37]
    end else if (_T_6 & 16'h14 == waddr) begin // @[VCR.scala 174:54]
      reg_5 <= io_host_w_bits_data; // @[VCR.scala 175:19]
    end
    if (reset) begin // @[VCR.scala 108:37]
      reg_6 <= 32'h0; // @[VCR.scala 108:37]
    end else if (_T_6 & 16'h18 == waddr) begin // @[VCR.scala 174:54]
      reg_6 <= io_host_w_bits_data; // @[VCR.scala 175:19]
    end
    if (reset) begin // @[VCR.scala 108:37]
      reg_7 <= 32'h0; // @[VCR.scala 108:37]
    end else if (_T_6 & 16'h1c == waddr) begin // @[VCR.scala 174:54]
      reg_7 <= io_host_w_bits_data; // @[VCR.scala 175:19]
    end
    if (reset) begin // @[VCR.scala 108:37]
      reg_8 <= 32'h0; // @[VCR.scala 108:37]
    end else if (_T_6 & 16'h20 == waddr) begin // @[VCR.scala 174:54]
      reg_8 <= io_host_w_bits_data; // @[VCR.scala 175:19]
    end
    if (reset) begin // @[VCR.scala 108:37]
      reg_9 <= 32'h0; // @[VCR.scala 108:37]
    end else if (io_vcr_ucnt_0_valid) begin // @[VCR.scala 200:32]
      reg_9 <= io_vcr_ucnt_0_bits; // @[VCR.scala 201:19]
    end else if (_T_6 & 16'h24 == waddr) begin // @[VCR.scala 202:60]
      reg_9 <= io_host_w_bits_data; // @[VCR.scala 203:19]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  waddr = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  wstate = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  rstate = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  rdata = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  reg_0 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  reg_1 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  reg_2 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  reg_3 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  reg_4 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  reg_5 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  reg_6 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  reg_7 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  reg_8 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  reg_9 = _RAND_13[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_addr,
  input  [3:0]  io_enq_bits_len,
  input  [20:0] io_enq_bits_tag,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_addr,
  output [3:0]  io_deq_bits_len,
  output [20:0] io_deq_bits_tag
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram_addr [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_addr_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_addr_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [31:0] ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [31:0] ram_addr_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_addr_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_addr_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_addr_MPORT_en; // @[Decoupled.scala 259:95]
  reg [3:0] ram_len [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_len_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_len_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [3:0] ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [3:0] ram_len_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_len_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_len_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_len_MPORT_en; // @[Decoupled.scala 259:95]
  reg [20:0] ram_tag [0:0]; // @[Decoupled.scala 259:95]
  wire  ram_tag_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire  ram_tag_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [20:0] ram_tag_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [20:0] ram_tag_MPORT_data; // @[Decoupled.scala 259:95]
  wire  ram_tag_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_tag_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_tag_MPORT_en; // @[Decoupled.scala 259:95]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  empty = ~maybe_full; // @[Decoupled.scala 264:28]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign ram_addr_io_deq_bits_MPORT_en = 1'h1;
  assign ram_addr_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_addr_io_deq_bits_MPORT_data = ram_addr[ram_addr_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_addr_MPORT_data = io_enq_bits_addr;
  assign ram_addr_MPORT_addr = 1'h0;
  assign ram_addr_MPORT_mask = 1'h1;
  assign ram_addr_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_len_io_deq_bits_MPORT_en = 1'h1;
  assign ram_len_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_len_io_deq_bits_MPORT_data = ram_len[ram_len_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_len_MPORT_data = io_enq_bits_len;
  assign ram_len_MPORT_addr = 1'h0;
  assign ram_len_MPORT_mask = 1'h1;
  assign ram_len_MPORT_en = io_enq_ready & io_enq_valid;
  assign ram_tag_io_deq_bits_MPORT_en = 1'h1;
  assign ram_tag_io_deq_bits_MPORT_addr = 1'h0;
  assign ram_tag_io_deq_bits_MPORT_data = ram_tag[ram_tag_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_tag_MPORT_data = io_enq_bits_tag;
  assign ram_tag_MPORT_addr = 1'h0;
  assign ram_tag_MPORT_mask = 1'h1;
  assign ram_tag_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~maybe_full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits_addr = ram_addr_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_len = ram_len_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  assign io_deq_bits_tag = ram_tag_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_addr_MPORT_en & ram_addr_MPORT_mask) begin
      ram_addr[ram_addr_MPORT_addr] <= ram_addr_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_len_MPORT_en & ram_len_MPORT_mask) begin
      ram_len[ram_len_MPORT_addr] <= ram_len_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (ram_tag_MPORT_en & ram_tag_MPORT_mask) begin
      ram_tag[ram_tag_MPORT_addr] <= ram_tag_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_addr[initvar] = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_len[initvar] = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    ram_tag[initvar] = _RAND_2[20:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module VME(
  input         clock,
  input         reset,
  input         io_mem_aw_ready,
  output        io_mem_aw_valid,
  output [31:0] io_mem_aw_bits_addr,
  output [3:0]  io_mem_aw_bits_len,
  input         io_mem_w_ready,
  output        io_mem_w_valid,
  output [63:0] io_mem_w_bits_data,
  output        io_mem_w_bits_last,
  output        io_mem_b_ready,
  input         io_mem_b_valid,
  input         io_mem_ar_ready,
  output        io_mem_ar_valid,
  output [31:0] io_mem_ar_bits_addr,
  output [7:0]  io_mem_ar_bits_id,
  output [3:0]  io_mem_ar_bits_len,
  input         io_mem_r_valid,
  input  [63:0] io_mem_r_bits_data,
  input         io_mem_r_bits_last,
  input  [7:0]  io_mem_r_bits_id,
  output        io_vme_rd_0_cmd_ready,
  input         io_vme_rd_0_cmd_valid,
  input  [31:0] io_vme_rd_0_cmd_bits_addr,
  input  [3:0]  io_vme_rd_0_cmd_bits_len,
  input         io_vme_rd_0_data_ready,
  output        io_vme_rd_0_data_valid,
  output [63:0] io_vme_rd_0_data_bits_data,
  output        io_vme_rd_1_cmd_ready,
  input         io_vme_rd_1_cmd_valid,
  input  [31:0] io_vme_rd_1_cmd_bits_addr,
  input  [3:0]  io_vme_rd_1_cmd_bits_len,
  input  [20:0] io_vme_rd_1_cmd_bits_tag,
  output        io_vme_rd_1_data_valid,
  output [63:0] io_vme_rd_1_data_bits_data,
  output [20:0] io_vme_rd_1_data_bits_tag,
  output        io_vme_rd_1_data_bits_last,
  output        io_vme_rd_2_cmd_ready,
  input         io_vme_rd_2_cmd_valid,
  input  [31:0] io_vme_rd_2_cmd_bits_addr,
  input  [3:0]  io_vme_rd_2_cmd_bits_len,
  input  [20:0] io_vme_rd_2_cmd_bits_tag,
  output        io_vme_rd_2_data_valid,
  output [63:0] io_vme_rd_2_data_bits_data,
  output [20:0] io_vme_rd_2_data_bits_tag,
  output        io_vme_rd_3_cmd_ready,
  input         io_vme_rd_3_cmd_valid,
  input  [31:0] io_vme_rd_3_cmd_bits_addr,
  input  [3:0]  io_vme_rd_3_cmd_bits_len,
  input  [20:0] io_vme_rd_3_cmd_bits_tag,
  output        io_vme_rd_3_data_valid,
  output [63:0] io_vme_rd_3_data_bits_data,
  output [20:0] io_vme_rd_3_data_bits_tag,
  output        io_vme_rd_4_cmd_ready,
  input         io_vme_rd_4_cmd_valid,
  input  [31:0] io_vme_rd_4_cmd_bits_addr,
  input  [3:0]  io_vme_rd_4_cmd_bits_len,
  input  [20:0] io_vme_rd_4_cmd_bits_tag,
  output        io_vme_rd_4_data_valid,
  output [63:0] io_vme_rd_4_data_bits_data,
  output [20:0] io_vme_rd_4_data_bits_tag,
  output        io_vme_wr_0_cmd_ready,
  input         io_vme_wr_0_cmd_valid,
  input  [31:0] io_vme_wr_0_cmd_bits_addr,
  input  [3:0]  io_vme_wr_0_cmd_bits_len,
  output        io_vme_wr_0_data_ready,
  input         io_vme_wr_0_data_valid,
  input  [63:0] io_vme_wr_0_data_bits_data,
  output        io_vme_wr_0_ack
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] vmeTag_array_client_id [0:15]; // @[VME.scala 189:33]
  wire  vmeTag_array_client_id_localTag_out_MPORT_en; // @[VME.scala 189:33]
  wire [3:0] vmeTag_array_client_id_localTag_out_MPORT_addr; // @[VME.scala 189:33]
  wire [2:0] vmeTag_array_client_id_localTag_out_MPORT_data; // @[VME.scala 189:33]
  wire [2:0] vmeTag_array_client_id_rdwrPort_data; // @[VME.scala 189:33]
  wire [3:0] vmeTag_array_client_id_rdwrPort_addr; // @[VME.scala 189:33]
  wire  vmeTag_array_client_id_rdwrPort_mask; // @[VME.scala 189:33]
  wire  vmeTag_array_client_id_rdwrPort_en; // @[VME.scala 189:33]
  reg  vmeTag_array_client_id_localTag_out_MPORT_en_pipe_0;
  reg [3:0] vmeTag_array_client_id_localTag_out_MPORT_addr_pipe_0;
  reg [20:0] vmeTag_array_client_tag [0:15]; // @[VME.scala 189:33]
  wire  vmeTag_array_client_tag_localTag_out_MPORT_en; // @[VME.scala 189:33]
  wire [3:0] vmeTag_array_client_tag_localTag_out_MPORT_addr; // @[VME.scala 189:33]
  wire [20:0] vmeTag_array_client_tag_localTag_out_MPORT_data; // @[VME.scala 189:33]
  wire [20:0] vmeTag_array_client_tag_rdwrPort_data; // @[VME.scala 189:33]
  wire [3:0] vmeTag_array_client_tag_rdwrPort_addr; // @[VME.scala 189:33]
  wire  vmeTag_array_client_tag_rdwrPort_mask; // @[VME.scala 189:33]
  wire  vmeTag_array_client_tag_rdwrPort_en; // @[VME.scala 189:33]
  reg  vmeTag_array_client_tag_localTag_out_MPORT_en_pipe_0;
  reg [3:0] vmeTag_array_client_tag_localTag_out_MPORT_addr_pipe_0;
  wire  VMEcmd_Qs_0_clock; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_0_reset; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_0_io_enq_ready; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_0_io_enq_valid; // @[VME.scala 216:45]
  wire [31:0] VMEcmd_Qs_0_io_enq_bits_addr; // @[VME.scala 216:45]
  wire [3:0] VMEcmd_Qs_0_io_enq_bits_len; // @[VME.scala 216:45]
  wire [20:0] VMEcmd_Qs_0_io_enq_bits_tag; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_0_io_deq_ready; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_0_io_deq_valid; // @[VME.scala 216:45]
  wire [31:0] VMEcmd_Qs_0_io_deq_bits_addr; // @[VME.scala 216:45]
  wire [3:0] VMEcmd_Qs_0_io_deq_bits_len; // @[VME.scala 216:45]
  wire [20:0] VMEcmd_Qs_0_io_deq_bits_tag; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_1_clock; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_1_reset; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_1_io_enq_ready; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_1_io_enq_valid; // @[VME.scala 216:45]
  wire [31:0] VMEcmd_Qs_1_io_enq_bits_addr; // @[VME.scala 216:45]
  wire [3:0] VMEcmd_Qs_1_io_enq_bits_len; // @[VME.scala 216:45]
  wire [20:0] VMEcmd_Qs_1_io_enq_bits_tag; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_1_io_deq_ready; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_1_io_deq_valid; // @[VME.scala 216:45]
  wire [31:0] VMEcmd_Qs_1_io_deq_bits_addr; // @[VME.scala 216:45]
  wire [3:0] VMEcmd_Qs_1_io_deq_bits_len; // @[VME.scala 216:45]
  wire [20:0] VMEcmd_Qs_1_io_deq_bits_tag; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_2_clock; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_2_reset; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_2_io_enq_ready; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_2_io_enq_valid; // @[VME.scala 216:45]
  wire [31:0] VMEcmd_Qs_2_io_enq_bits_addr; // @[VME.scala 216:45]
  wire [3:0] VMEcmd_Qs_2_io_enq_bits_len; // @[VME.scala 216:45]
  wire [20:0] VMEcmd_Qs_2_io_enq_bits_tag; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_2_io_deq_ready; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_2_io_deq_valid; // @[VME.scala 216:45]
  wire [31:0] VMEcmd_Qs_2_io_deq_bits_addr; // @[VME.scala 216:45]
  wire [3:0] VMEcmd_Qs_2_io_deq_bits_len; // @[VME.scala 216:45]
  wire [20:0] VMEcmd_Qs_2_io_deq_bits_tag; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_3_clock; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_3_reset; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_3_io_enq_ready; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_3_io_enq_valid; // @[VME.scala 216:45]
  wire [31:0] VMEcmd_Qs_3_io_enq_bits_addr; // @[VME.scala 216:45]
  wire [3:0] VMEcmd_Qs_3_io_enq_bits_len; // @[VME.scala 216:45]
  wire [20:0] VMEcmd_Qs_3_io_enq_bits_tag; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_3_io_deq_ready; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_3_io_deq_valid; // @[VME.scala 216:45]
  wire [31:0] VMEcmd_Qs_3_io_deq_bits_addr; // @[VME.scala 216:45]
  wire [3:0] VMEcmd_Qs_3_io_deq_bits_len; // @[VME.scala 216:45]
  wire [20:0] VMEcmd_Qs_3_io_deq_bits_tag; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_4_clock; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_4_reset; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_4_io_enq_ready; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_4_io_enq_valid; // @[VME.scala 216:45]
  wire [31:0] VMEcmd_Qs_4_io_enq_bits_addr; // @[VME.scala 216:45]
  wire [3:0] VMEcmd_Qs_4_io_enq_bits_len; // @[VME.scala 216:45]
  wire [20:0] VMEcmd_Qs_4_io_enq_bits_tag; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_4_io_deq_ready; // @[VME.scala 216:45]
  wire  VMEcmd_Qs_4_io_deq_valid; // @[VME.scala 216:45]
  wire [31:0] VMEcmd_Qs_4_io_deq_bits_addr; // @[VME.scala 216:45]
  wire [3:0] VMEcmd_Qs_4_io_deq_bits_len; // @[VME.scala 216:45]
  wire [20:0] VMEcmd_Qs_4_io_deq_bits_tag; // @[VME.scala 216:45]
  reg [15:0] availableEntries; // @[VME.scala 197:33]
  wire  oneHotIdx_0 = availableEntries[0]; // @[VME.scala 224:11]
  wire  oneHotIdx_1 = availableEntries[1] & ~(|oneHotIdx_0); // @[VME.scala 227:20]
  wire  oneHotIdx_2 = availableEntries[2] & ~(|availableEntries[1:0]); // @[VME.scala 227:20]
  wire  oneHotIdx_3 = availableEntries[3] & ~(|availableEntries[2:0]); // @[VME.scala 227:20]
  wire  oneHotIdx_4 = availableEntries[4] & ~(|availableEntries[3:0]); // @[VME.scala 227:20]
  wire  oneHotIdx_5 = availableEntries[5] & ~(|availableEntries[4:0]); // @[VME.scala 227:20]
  wire  oneHotIdx_6 = availableEntries[6] & ~(|availableEntries[5:0]); // @[VME.scala 227:20]
  wire  oneHotIdx_7 = availableEntries[7] & ~(|availableEntries[6:0]); // @[VME.scala 227:20]
  wire  oneHotIdx_8 = availableEntries[8] & ~(|availableEntries[7:0]); // @[VME.scala 227:20]
  wire  oneHotIdx_9 = availableEntries[9] & ~(|availableEntries[8:0]); // @[VME.scala 227:20]
  wire  oneHotIdx_10 = availableEntries[10] & ~(|availableEntries[9:0]); // @[VME.scala 227:20]
  wire  oneHotIdx_11 = availableEntries[11] & ~(|availableEntries[10:0]); // @[VME.scala 227:20]
  wire  oneHotIdx_12 = availableEntries[12] & ~(|availableEntries[11:0]); // @[VME.scala 227:20]
  wire  oneHotIdx_13 = availableEntries[13] & ~(|availableEntries[12:0]); // @[VME.scala 227:20]
  wire  oneHotIdx_14 = availableEntries[14] & ~(|availableEntries[13:0]); // @[VME.scala 227:20]
  wire  oneHotIdx_15 = availableEntries[15] & ~(|availableEntries[14:0]); // @[VME.scala 227:20]
  wire [7:0] oHot_lo = {oneHotIdx_7,oneHotIdx_6,oneHotIdx_5,oneHotIdx_4,oneHotIdx_3,oneHotIdx_2,oneHotIdx_1,oneHotIdx_0}
    ; // @[VME.scala 230:35]
  wire [15:0] resetEntry = {oneHotIdx_15,oneHotIdx_14,oneHotIdx_13,oneHotIdx_12,oneHotIdx_11,oneHotIdx_10,oneHotIdx_9,
    oneHotIdx_8,oHot_lo}; // @[VME.scala 230:35]
  wire [15:0] _newVec_T = ~resetEntry; // @[VME.scala 231:22]
  wire [15:0] newEntry = availableEntries & _newVec_T; // @[VME.scala 231:20]
  wire [3:0] _bitPostn_T = oneHotIdx_14 ? 4'he : 4'hf; // @[Mux.scala 47:70]
  wire [3:0] _bitPostn_T_1 = oneHotIdx_13 ? 4'hd : _bitPostn_T; // @[Mux.scala 47:70]
  wire [3:0] _bitPostn_T_2 = oneHotIdx_12 ? 4'hc : _bitPostn_T_1; // @[Mux.scala 47:70]
  wire [3:0] _bitPostn_T_3 = oneHotIdx_11 ? 4'hb : _bitPostn_T_2; // @[Mux.scala 47:70]
  wire [3:0] _bitPostn_T_4 = oneHotIdx_10 ? 4'ha : _bitPostn_T_3; // @[Mux.scala 47:70]
  wire [3:0] _bitPostn_T_5 = oneHotIdx_9 ? 4'h9 : _bitPostn_T_4; // @[Mux.scala 47:70]
  wire [3:0] _bitPostn_T_6 = oneHotIdx_8 ? 4'h8 : _bitPostn_T_5; // @[Mux.scala 47:70]
  wire [3:0] _bitPostn_T_7 = oneHotIdx_7 ? 4'h7 : _bitPostn_T_6; // @[Mux.scala 47:70]
  wire [3:0] _bitPostn_T_8 = oneHotIdx_6 ? 4'h6 : _bitPostn_T_7; // @[Mux.scala 47:70]
  wire [3:0] _bitPostn_T_9 = oneHotIdx_5 ? 4'h5 : _bitPostn_T_8; // @[Mux.scala 47:70]
  wire [3:0] _bitPostn_T_10 = oneHotIdx_4 ? 4'h4 : _bitPostn_T_9; // @[Mux.scala 47:70]
  wire [3:0] _bitPostn_T_11 = oneHotIdx_3 ? 4'h3 : _bitPostn_T_10; // @[Mux.scala 47:70]
  wire [3:0] _bitPostn_T_12 = oneHotIdx_2 ? 4'h2 : _bitPostn_T_11; // @[Mux.scala 47:70]
  wire [3:0] _bitPostn_T_13 = oneHotIdx_1 ? 4'h1 : _bitPostn_T_12; // @[Mux.scala 47:70]
  wire [3:0] firstPostn = oneHotIdx_0 ? 4'h0 : _bitPostn_T_13; // @[Mux.scala 47:70]
  wire  _T = io_mem_r_bits_last & io_mem_r_valid; // @[VME.scala 201:27]
  wire [7:0] updateEntry_lo = {8'h7 == io_mem_r_bits_id,8'h6 == io_mem_r_bits_id,8'h5 == io_mem_r_bits_id,8'h4 ==
    io_mem_r_bits_id,8'h3 == io_mem_r_bits_id,8'h2 == io_mem_r_bits_id,8'h1 == io_mem_r_bits_id,8'h0 == io_mem_r_bits_id
    }; // @[VME.scala 213:108]
  wire [15:0] _updateEntry_T_16 = {8'hf == io_mem_r_bits_id,8'he == io_mem_r_bits_id,8'hd == io_mem_r_bits_id,8'hc ==
    io_mem_r_bits_id,8'hb == io_mem_r_bits_id,8'ha == io_mem_r_bits_id,8'h9 == io_mem_r_bits_id,8'h8 == io_mem_r_bits_id
    ,updateEntry_lo}; // @[VME.scala 213:108]
  wire [15:0] updateEntry = reset ? 16'h0 : _updateEntry_T_16; // @[VME.scala 208:21 210:15 213:15]
  wire [15:0] _availableEntriesNext_T = updateEntry | availableEntries; // @[VME.scala 202:39]
  wire  _T_1 = availableEntries != 16'h0; // @[VME.scala 203:53]
  wire  any_cmd_valid = VMEcmd_Qs_0_io_deq_valid | VMEcmd_Qs_1_io_deq_valid | VMEcmd_Qs_2_io_deq_valid |
    VMEcmd_Qs_3_io_deq_valid | VMEcmd_Qs_4_io_deq_valid; // @[VME.scala 243:69]
  wire  availableEntriesEn = io_mem_ar_ready & any_cmd_valid; // @[VME.scala 244:41]
  wire  _T_4 = ~_T; // @[VME.scala 203:64]
  wire [2:0] _vme_select_T = VMEcmd_Qs_4_io_deq_valid ? 3'h4 : 3'h5; // @[Mux.scala 47:70]
  wire [2:0] _vme_select_T_1 = VMEcmd_Qs_3_io_deq_valid ? 3'h3 : _vme_select_T; // @[Mux.scala 47:70]
  wire [2:0] _vme_select_T_2 = VMEcmd_Qs_2_io_deq_valid ? 3'h2 : _vme_select_T_1; // @[Mux.scala 47:70]
  wire [2:0] _vme_select_T_3 = VMEcmd_Qs_1_io_deq_valid ? 3'h1 : _vme_select_T_2; // @[Mux.scala 47:70]
  wire [2:0] vme_select = VMEcmd_Qs_0_io_deq_valid ? 3'h0 : _vme_select_T_3; // @[Mux.scala 47:70]
  wire  _VMEcmd_Qs_0_io_deq_ready_T = vme_select == 3'h0; // @[VME.scala 250:17]
  wire  _VMEcmd_Qs_0_io_deq_ready_T_1 = io_mem_ar_ready & _VMEcmd_Qs_0_io_deq_ready_T; // @[VME.scala 249:50]
  wire  _VMEcmd_Qs_1_io_deq_ready_T = vme_select == 3'h1; // @[VME.scala 250:17]
  wire  _VMEcmd_Qs_1_io_deq_ready_T_1 = io_mem_ar_ready & _VMEcmd_Qs_1_io_deq_ready_T; // @[VME.scala 249:50]
  wire  _VMEcmd_Qs_2_io_deq_ready_T = vme_select == 3'h2; // @[VME.scala 250:17]
  wire  _VMEcmd_Qs_2_io_deq_ready_T_1 = io_mem_ar_ready & _VMEcmd_Qs_2_io_deq_ready_T; // @[VME.scala 249:50]
  wire  _VMEcmd_Qs_3_io_deq_ready_T = vme_select == 3'h3; // @[VME.scala 250:17]
  wire  _VMEcmd_Qs_3_io_deq_ready_T_1 = io_mem_ar_ready & _VMEcmd_Qs_3_io_deq_ready_T; // @[VME.scala 249:50]
  wire  _VMEcmd_Qs_4_io_deq_ready_T = vme_select == 3'h4; // @[VME.scala 250:17]
  wire  _VMEcmd_Qs_4_io_deq_ready_T_1 = io_mem_ar_ready & _VMEcmd_Qs_4_io_deq_ready_T; // @[VME.scala 249:50]
  wire  _any_cmd_ready_T_3 = VMEcmd_Qs_0_io_deq_ready | VMEcmd_Qs_1_io_deq_ready | VMEcmd_Qs_2_io_deq_ready |
    VMEcmd_Qs_3_io_deq_ready; // @[VME.scala 259:69]
  wire [20:0] _GEN_16 = VMEcmd_Qs_4_io_deq_ready ? VMEcmd_Qs_4_io_deq_bits_tag : 21'h0; // @[VME.scala 272:24 276:36 282:39]
  wire [20:0] _GEN_23 = VMEcmd_Qs_3_io_deq_ready ? VMEcmd_Qs_3_io_deq_bits_tag : _GEN_16; // @[VME.scala 276:36 282:39]
  wire [20:0] _GEN_30 = VMEcmd_Qs_2_io_deq_ready ? VMEcmd_Qs_2_io_deq_bits_tag : _GEN_23; // @[VME.scala 276:36 282:39]
  wire [20:0] _GEN_37 = VMEcmd_Qs_1_io_deq_ready ? VMEcmd_Qs_1_io_deq_bits_tag : _GEN_30; // @[VME.scala 276:36 282:39]
  wire [2:0] _GEN_15 = VMEcmd_Qs_4_io_deq_ready ? 3'h4 : 3'h0; // @[VME.scala 272:24 276:36 281:39]
  wire [2:0] _GEN_22 = VMEcmd_Qs_3_io_deq_ready ? 3'h3 : _GEN_15; // @[VME.scala 276:36 281:39]
  wire [2:0] _GEN_29 = VMEcmd_Qs_2_io_deq_ready ? 3'h2 : _GEN_22; // @[VME.scala 276:36 281:39]
  wire [2:0] _GEN_36 = VMEcmd_Qs_1_io_deq_ready ? 3'h1 : _GEN_29; // @[VME.scala 276:36 281:39]
  wire [31:0] _GEN_11 = VMEcmd_Qs_4_io_deq_ready ? VMEcmd_Qs_4_io_deq_bits_addr : 32'h0; // @[VME.scala 268:23 276:36 277:27]
  wire [3:0] _GEN_12 = VMEcmd_Qs_4_io_deq_ready ? VMEcmd_Qs_4_io_deq_bits_len : 4'h0; // @[VME.scala 269:23 276:36 278:27]
  wire  _GEN_13 = VMEcmd_Qs_4_io_deq_ready & VMEcmd_Qs_4_io_deq_valid; // @[VME.scala 270:23 276:36 279:27]
  wire [3:0] _GEN_14 = VMEcmd_Qs_4_io_deq_ready ? firstPostn : 4'h0; // @[VME.scala 271:23 276:36 280:27]
  wire [31:0] _GEN_18 = VMEcmd_Qs_3_io_deq_ready ? VMEcmd_Qs_3_io_deq_bits_addr : _GEN_11; // @[VME.scala 276:36 277:27]
  wire [3:0] _GEN_19 = VMEcmd_Qs_3_io_deq_ready ? VMEcmd_Qs_3_io_deq_bits_len : _GEN_12; // @[VME.scala 276:36 278:27]
  wire  _GEN_20 = VMEcmd_Qs_3_io_deq_ready ? VMEcmd_Qs_3_io_deq_valid : _GEN_13; // @[VME.scala 276:36 279:27]
  wire [3:0] _GEN_21 = VMEcmd_Qs_3_io_deq_ready ? firstPostn : _GEN_14; // @[VME.scala 276:36 280:27]
  wire [31:0] _GEN_25 = VMEcmd_Qs_2_io_deq_ready ? VMEcmd_Qs_2_io_deq_bits_addr : _GEN_18; // @[VME.scala 276:36 277:27]
  wire [3:0] _GEN_26 = VMEcmd_Qs_2_io_deq_ready ? VMEcmd_Qs_2_io_deq_bits_len : _GEN_19; // @[VME.scala 276:36 278:27]
  wire  _GEN_27 = VMEcmd_Qs_2_io_deq_ready ? VMEcmd_Qs_2_io_deq_valid : _GEN_20; // @[VME.scala 276:36 279:27]
  wire [3:0] _GEN_28 = VMEcmd_Qs_2_io_deq_ready ? firstPostn : _GEN_21; // @[VME.scala 276:36 280:27]
  wire [31:0] _GEN_32 = VMEcmd_Qs_1_io_deq_ready ? VMEcmd_Qs_1_io_deq_bits_addr : _GEN_25; // @[VME.scala 276:36 277:27]
  wire [3:0] _GEN_33 = VMEcmd_Qs_1_io_deq_ready ? VMEcmd_Qs_1_io_deq_bits_len : _GEN_26; // @[VME.scala 276:36 278:27]
  wire  _GEN_34 = VMEcmd_Qs_1_io_deq_ready ? VMEcmd_Qs_1_io_deq_valid : _GEN_27; // @[VME.scala 276:36 279:27]
  wire [3:0] _GEN_35 = VMEcmd_Qs_1_io_deq_ready ? firstPostn : _GEN_28; // @[VME.scala 276:36 280:27]
  wire [3:0] _GEN_42 = VMEcmd_Qs_0_io_deq_ready ? firstPostn : _GEN_35; // @[VME.scala 276:36 280:27]
  reg  io_vme_rd_0_data_valid_REG; // @[VME.scala 297:41]
  wire [2:0] localTag_out_client_id = vmeTag_array_client_id_localTag_out_MPORT_data; // @[VME.scala 194:27 293:24]
  wire  _io_vme_rd_0_data_valid_T_1 = io_vme_rd_0_data_valid_REG & localTag_out_client_id == 3'h0; // @[VME.scala 297:75]
  reg [63:0] io_vme_rd_0_data_bits_data_REG; // @[VME.scala 301:43]
  reg  io_vme_rd_1_data_valid_REG; // @[VME.scala 297:41]
  reg [63:0] io_vme_rd_1_data_bits_data_REG; // @[VME.scala 301:43]
  reg  io_vme_rd_1_data_bits_last_REG; // @[VME.scala 302:43]
  reg  io_vme_rd_2_data_valid_REG; // @[VME.scala 297:41]
  reg [63:0] io_vme_rd_2_data_bits_data_REG; // @[VME.scala 301:43]
  reg  io_vme_rd_3_data_valid_REG; // @[VME.scala 297:41]
  reg [63:0] io_vme_rd_3_data_bits_data_REG; // @[VME.scala 301:43]
  reg  io_vme_rd_4_data_valid_REG; // @[VME.scala 297:41]
  reg [63:0] io_vme_rd_4_data_bits_data_REG; // @[VME.scala 301:43]
  reg [3:0] wr_len; // @[VME.scala 307:23]
  reg [31:0] wr_addr; // @[VME.scala 308:24]
  reg [1:0] wstate; // @[VME.scala 310:23]
  reg [3:0] wr_cnt; // @[VME.scala 311:23]
  wire  _io_vme_wr_0_cmd_ready_T = wstate == 2'h0; // @[VME.scala 312:36]
  wire  _io_vme_wr_0_data_ready_T = wstate == 2'h2; // @[VME.scala 314:37]
  wire  _io_mem_w_bits_last_T = wr_cnt == wr_len; // @[VME.scala 322:32]
  wire  _T_32 = io_vme_wr_0_cmd_ready & io_vme_wr_0_cmd_valid; // @[Decoupled.scala 50:35]
  wire  _T_34 = io_mem_w_ready & io_mem_w_valid; // @[Decoupled.scala 50:35]
  wire [3:0] _wr_cnt_T_1 = wr_cnt + 4'h1; // @[VME.scala 333:22]
  wire [1:0] _GEN_52 = io_vme_wr_0_data_valid & io_mem_w_ready & _io_mem_w_bits_last_T ? 2'h3 : wstate; // @[VME.scala 347:76 348:16 310:23]
  wire [1:0] _GEN_53 = io_mem_b_valid ? 2'h0 : wstate; // @[VME.scala 352:28 353:16 310:23]
  wire [1:0] _GEN_54 = 2'h3 == wstate ? _GEN_53 : wstate; // @[VME.scala 335:17 310:23]
  Queue VMEcmd_Qs_0 ( // @[VME.scala 216:45]
    .clock(VMEcmd_Qs_0_clock),
    .reset(VMEcmd_Qs_0_reset),
    .io_enq_ready(VMEcmd_Qs_0_io_enq_ready),
    .io_enq_valid(VMEcmd_Qs_0_io_enq_valid),
    .io_enq_bits_addr(VMEcmd_Qs_0_io_enq_bits_addr),
    .io_enq_bits_len(VMEcmd_Qs_0_io_enq_bits_len),
    .io_enq_bits_tag(VMEcmd_Qs_0_io_enq_bits_tag),
    .io_deq_ready(VMEcmd_Qs_0_io_deq_ready),
    .io_deq_valid(VMEcmd_Qs_0_io_deq_valid),
    .io_deq_bits_addr(VMEcmd_Qs_0_io_deq_bits_addr),
    .io_deq_bits_len(VMEcmd_Qs_0_io_deq_bits_len),
    .io_deq_bits_tag(VMEcmd_Qs_0_io_deq_bits_tag)
  );
  Queue VMEcmd_Qs_1 ( // @[VME.scala 216:45]
    .clock(VMEcmd_Qs_1_clock),
    .reset(VMEcmd_Qs_1_reset),
    .io_enq_ready(VMEcmd_Qs_1_io_enq_ready),
    .io_enq_valid(VMEcmd_Qs_1_io_enq_valid),
    .io_enq_bits_addr(VMEcmd_Qs_1_io_enq_bits_addr),
    .io_enq_bits_len(VMEcmd_Qs_1_io_enq_bits_len),
    .io_enq_bits_tag(VMEcmd_Qs_1_io_enq_bits_tag),
    .io_deq_ready(VMEcmd_Qs_1_io_deq_ready),
    .io_deq_valid(VMEcmd_Qs_1_io_deq_valid),
    .io_deq_bits_addr(VMEcmd_Qs_1_io_deq_bits_addr),
    .io_deq_bits_len(VMEcmd_Qs_1_io_deq_bits_len),
    .io_deq_bits_tag(VMEcmd_Qs_1_io_deq_bits_tag)
  );
  Queue VMEcmd_Qs_2 ( // @[VME.scala 216:45]
    .clock(VMEcmd_Qs_2_clock),
    .reset(VMEcmd_Qs_2_reset),
    .io_enq_ready(VMEcmd_Qs_2_io_enq_ready),
    .io_enq_valid(VMEcmd_Qs_2_io_enq_valid),
    .io_enq_bits_addr(VMEcmd_Qs_2_io_enq_bits_addr),
    .io_enq_bits_len(VMEcmd_Qs_2_io_enq_bits_len),
    .io_enq_bits_tag(VMEcmd_Qs_2_io_enq_bits_tag),
    .io_deq_ready(VMEcmd_Qs_2_io_deq_ready),
    .io_deq_valid(VMEcmd_Qs_2_io_deq_valid),
    .io_deq_bits_addr(VMEcmd_Qs_2_io_deq_bits_addr),
    .io_deq_bits_len(VMEcmd_Qs_2_io_deq_bits_len),
    .io_deq_bits_tag(VMEcmd_Qs_2_io_deq_bits_tag)
  );
  Queue VMEcmd_Qs_3 ( // @[VME.scala 216:45]
    .clock(VMEcmd_Qs_3_clock),
    .reset(VMEcmd_Qs_3_reset),
    .io_enq_ready(VMEcmd_Qs_3_io_enq_ready),
    .io_enq_valid(VMEcmd_Qs_3_io_enq_valid),
    .io_enq_bits_addr(VMEcmd_Qs_3_io_enq_bits_addr),
    .io_enq_bits_len(VMEcmd_Qs_3_io_enq_bits_len),
    .io_enq_bits_tag(VMEcmd_Qs_3_io_enq_bits_tag),
    .io_deq_ready(VMEcmd_Qs_3_io_deq_ready),
    .io_deq_valid(VMEcmd_Qs_3_io_deq_valid),
    .io_deq_bits_addr(VMEcmd_Qs_3_io_deq_bits_addr),
    .io_deq_bits_len(VMEcmd_Qs_3_io_deq_bits_len),
    .io_deq_bits_tag(VMEcmd_Qs_3_io_deq_bits_tag)
  );
  Queue VMEcmd_Qs_4 ( // @[VME.scala 216:45]
    .clock(VMEcmd_Qs_4_clock),
    .reset(VMEcmd_Qs_4_reset),
    .io_enq_ready(VMEcmd_Qs_4_io_enq_ready),
    .io_enq_valid(VMEcmd_Qs_4_io_enq_valid),
    .io_enq_bits_addr(VMEcmd_Qs_4_io_enq_bits_addr),
    .io_enq_bits_len(VMEcmd_Qs_4_io_enq_bits_len),
    .io_enq_bits_tag(VMEcmd_Qs_4_io_enq_bits_tag),
    .io_deq_ready(VMEcmd_Qs_4_io_deq_ready),
    .io_deq_valid(VMEcmd_Qs_4_io_deq_valid),
    .io_deq_bits_addr(VMEcmd_Qs_4_io_deq_bits_addr),
    .io_deq_bits_len(VMEcmd_Qs_4_io_deq_bits_len),
    .io_deq_bits_tag(VMEcmd_Qs_4_io_deq_bits_tag)
  );
  assign vmeTag_array_client_id_localTag_out_MPORT_en = vmeTag_array_client_id_localTag_out_MPORT_en_pipe_0;
  assign vmeTag_array_client_id_localTag_out_MPORT_addr = vmeTag_array_client_id_localTag_out_MPORT_addr_pipe_0;
  assign vmeTag_array_client_id_localTag_out_MPORT_data =
    vmeTag_array_client_id[vmeTag_array_client_id_localTag_out_MPORT_addr]; // @[VME.scala 189:33]
  assign vmeTag_array_client_id_rdwrPort_data = VMEcmd_Qs_0_io_deq_ready ? 3'h0 : _GEN_36;
  assign vmeTag_array_client_id_rdwrPort_addr = oneHotIdx_0 ? 4'h0 : _bitPostn_T_13;
  assign vmeTag_array_client_id_rdwrPort_mask = 1'h1;
  assign vmeTag_array_client_id_rdwrPort_en = _any_cmd_ready_T_3 | VMEcmd_Qs_4_io_deq_ready;
  assign vmeTag_array_client_tag_localTag_out_MPORT_en = vmeTag_array_client_tag_localTag_out_MPORT_en_pipe_0;
  assign vmeTag_array_client_tag_localTag_out_MPORT_addr = vmeTag_array_client_tag_localTag_out_MPORT_addr_pipe_0;
  assign vmeTag_array_client_tag_localTag_out_MPORT_data =
    vmeTag_array_client_tag[vmeTag_array_client_tag_localTag_out_MPORT_addr]; // @[VME.scala 189:33]
  assign vmeTag_array_client_tag_rdwrPort_data = VMEcmd_Qs_0_io_deq_ready ? VMEcmd_Qs_0_io_deq_bits_tag : _GEN_37;
  assign vmeTag_array_client_tag_rdwrPort_addr = oneHotIdx_0 ? 4'h0 : _bitPostn_T_13;
  assign vmeTag_array_client_tag_rdwrPort_mask = 1'h1;
  assign vmeTag_array_client_tag_rdwrPort_en = _any_cmd_ready_T_3 | VMEcmd_Qs_4_io_deq_ready;
  assign io_mem_aw_valid = wstate == 2'h1; // @[VME.scala 315:29]
  assign io_mem_aw_bits_addr = wr_addr; // @[VME.scala 316:23]
  assign io_mem_aw_bits_len = wr_len; // @[VME.scala 317:22]
  assign io_mem_w_valid = _io_vme_wr_0_data_ready_T & io_vme_wr_0_data_valid; // @[VME.scala 319:43]
  assign io_mem_w_bits_data = io_vme_wr_0_data_bits_data; // @[VME.scala 320:22]
  assign io_mem_w_bits_last = wr_cnt == wr_len; // @[VME.scala 322:32]
  assign io_mem_b_ready = wstate == 2'h3; // @[VME.scala 324:28]
  assign io_mem_ar_valid = VMEcmd_Qs_0_io_deq_ready ? VMEcmd_Qs_0_io_deq_valid : _GEN_34; // @[VME.scala 276:36 279:27]
  assign io_mem_ar_bits_addr = VMEcmd_Qs_0_io_deq_ready ? VMEcmd_Qs_0_io_deq_bits_addr : _GEN_32; // @[VME.scala 276:36 277:27]
  assign io_mem_ar_bits_id = {{4'd0}, _GEN_42};
  assign io_mem_ar_bits_len = VMEcmd_Qs_0_io_deq_ready ? VMEcmd_Qs_0_io_deq_bits_len : _GEN_33; // @[VME.scala 276:36 278:27]
  assign io_vme_rd_0_cmd_ready = VMEcmd_Qs_0_io_enq_ready; // @[VME.scala 252:28]
  assign io_vme_rd_0_data_valid = _io_vme_rd_0_data_valid_T_1 & io_vme_rd_0_data_ready; // @[VME.scala 298:5]
  assign io_vme_rd_0_data_bits_data = io_vme_rd_0_data_bits_data_REG; // @[VME.scala 301:33]
  assign io_vme_rd_1_cmd_ready = VMEcmd_Qs_1_io_enq_ready; // @[VME.scala 252:28]
  assign io_vme_rd_1_data_valid = io_vme_rd_1_data_valid_REG & localTag_out_client_id == 3'h1; // @[VME.scala 297:75]
  assign io_vme_rd_1_data_bits_data = io_vme_rd_1_data_bits_data_REG; // @[VME.scala 301:33]
  assign io_vme_rd_1_data_bits_tag = vmeTag_array_client_tag_localTag_out_MPORT_data; // @[VME.scala 194:27 293:24]
  assign io_vme_rd_1_data_bits_last = io_vme_rd_1_data_bits_last_REG; // @[VME.scala 302:33]
  assign io_vme_rd_2_cmd_ready = VMEcmd_Qs_2_io_enq_ready; // @[VME.scala 252:28]
  assign io_vme_rd_2_data_valid = io_vme_rd_2_data_valid_REG & localTag_out_client_id == 3'h2; // @[VME.scala 297:75]
  assign io_vme_rd_2_data_bits_data = io_vme_rd_2_data_bits_data_REG; // @[VME.scala 301:33]
  assign io_vme_rd_2_data_bits_tag = vmeTag_array_client_tag_localTag_out_MPORT_data; // @[VME.scala 194:27 293:24]
  assign io_vme_rd_3_cmd_ready = VMEcmd_Qs_3_io_enq_ready; // @[VME.scala 252:28]
  assign io_vme_rd_3_data_valid = io_vme_rd_3_data_valid_REG & localTag_out_client_id == 3'h3; // @[VME.scala 297:75]
  assign io_vme_rd_3_data_bits_data = io_vme_rd_3_data_bits_data_REG; // @[VME.scala 301:33]
  assign io_vme_rd_3_data_bits_tag = vmeTag_array_client_tag_localTag_out_MPORT_data; // @[VME.scala 194:27 293:24]
  assign io_vme_rd_4_cmd_ready = VMEcmd_Qs_4_io_enq_ready; // @[VME.scala 252:28]
  assign io_vme_rd_4_data_valid = io_vme_rd_4_data_valid_REG & localTag_out_client_id == 3'h4; // @[VME.scala 297:75]
  assign io_vme_rd_4_data_bits_data = io_vme_rd_4_data_bits_data_REG; // @[VME.scala 301:33]
  assign io_vme_rd_4_data_bits_tag = vmeTag_array_client_tag_localTag_out_MPORT_data; // @[VME.scala 194:27 293:24]
  assign io_vme_wr_0_cmd_ready = wstate == 2'h0; // @[VME.scala 312:36]
  assign io_vme_wr_0_data_ready = wstate == 2'h2 & io_mem_w_ready; // @[VME.scala 314:52]
  assign io_vme_wr_0_ack = io_mem_b_ready & io_mem_b_valid; // @[Decoupled.scala 50:35]
  assign VMEcmd_Qs_0_clock = clock;
  assign VMEcmd_Qs_0_reset = reset;
  assign VMEcmd_Qs_0_io_enq_valid = io_vme_rd_0_cmd_valid & VMEcmd_Qs_0_io_enq_ready; // @[VME.scala 247:58]
  assign VMEcmd_Qs_0_io_enq_bits_addr = io_vme_rd_0_cmd_bits_addr; // @[VME.scala 248:31]
  assign VMEcmd_Qs_0_io_enq_bits_len = io_vme_rd_0_cmd_bits_len; // @[VME.scala 248:31]
  assign VMEcmd_Qs_0_io_enq_bits_tag = 21'h0; // @[VME.scala 248:31]
  assign VMEcmd_Qs_0_io_deq_ready = _VMEcmd_Qs_0_io_deq_ready_T_1 & _T_1 & _T_4; // @[VME.scala 250:62]
  assign VMEcmd_Qs_1_clock = clock;
  assign VMEcmd_Qs_1_reset = reset;
  assign VMEcmd_Qs_1_io_enq_valid = io_vme_rd_1_cmd_valid & VMEcmd_Qs_1_io_enq_ready; // @[VME.scala 247:58]
  assign VMEcmd_Qs_1_io_enq_bits_addr = io_vme_rd_1_cmd_bits_addr; // @[VME.scala 248:31]
  assign VMEcmd_Qs_1_io_enq_bits_len = io_vme_rd_1_cmd_bits_len; // @[VME.scala 248:31]
  assign VMEcmd_Qs_1_io_enq_bits_tag = io_vme_rd_1_cmd_bits_tag; // @[VME.scala 248:31]
  assign VMEcmd_Qs_1_io_deq_ready = _VMEcmd_Qs_1_io_deq_ready_T_1 & _T_1 & _T_4; // @[VME.scala 250:62]
  assign VMEcmd_Qs_2_clock = clock;
  assign VMEcmd_Qs_2_reset = reset;
  assign VMEcmd_Qs_2_io_enq_valid = io_vme_rd_2_cmd_valid & VMEcmd_Qs_2_io_enq_ready; // @[VME.scala 247:58]
  assign VMEcmd_Qs_2_io_enq_bits_addr = io_vme_rd_2_cmd_bits_addr; // @[VME.scala 248:31]
  assign VMEcmd_Qs_2_io_enq_bits_len = io_vme_rd_2_cmd_bits_len; // @[VME.scala 248:31]
  assign VMEcmd_Qs_2_io_enq_bits_tag = io_vme_rd_2_cmd_bits_tag; // @[VME.scala 248:31]
  assign VMEcmd_Qs_2_io_deq_ready = _VMEcmd_Qs_2_io_deq_ready_T_1 & _T_1 & _T_4; // @[VME.scala 250:62]
  assign VMEcmd_Qs_3_clock = clock;
  assign VMEcmd_Qs_3_reset = reset;
  assign VMEcmd_Qs_3_io_enq_valid = io_vme_rd_3_cmd_valid & VMEcmd_Qs_3_io_enq_ready; // @[VME.scala 247:58]
  assign VMEcmd_Qs_3_io_enq_bits_addr = io_vme_rd_3_cmd_bits_addr; // @[VME.scala 248:31]
  assign VMEcmd_Qs_3_io_enq_bits_len = io_vme_rd_3_cmd_bits_len; // @[VME.scala 248:31]
  assign VMEcmd_Qs_3_io_enq_bits_tag = io_vme_rd_3_cmd_bits_tag; // @[VME.scala 248:31]
  assign VMEcmd_Qs_3_io_deq_ready = _VMEcmd_Qs_3_io_deq_ready_T_1 & _T_1 & _T_4; // @[VME.scala 250:62]
  assign VMEcmd_Qs_4_clock = clock;
  assign VMEcmd_Qs_4_reset = reset;
  assign VMEcmd_Qs_4_io_enq_valid = io_vme_rd_4_cmd_valid & VMEcmd_Qs_4_io_enq_ready; // @[VME.scala 247:58]
  assign VMEcmd_Qs_4_io_enq_bits_addr = io_vme_rd_4_cmd_bits_addr; // @[VME.scala 248:31]
  assign VMEcmd_Qs_4_io_enq_bits_len = io_vme_rd_4_cmd_bits_len; // @[VME.scala 248:31]
  assign VMEcmd_Qs_4_io_enq_bits_tag = io_vme_rd_4_cmd_bits_tag; // @[VME.scala 248:31]
  assign VMEcmd_Qs_4_io_deq_ready = _VMEcmd_Qs_4_io_deq_ready_T_1 & _T_1 & _T_4; // @[VME.scala 250:62]
  always @(posedge clock) begin
    if (vmeTag_array_client_id_rdwrPort_en & vmeTag_array_client_id_rdwrPort_mask) begin
      vmeTag_array_client_id[vmeTag_array_client_id_rdwrPort_addr] <= vmeTag_array_client_id_rdwrPort_data; // @[VME.scala 189:33]
    end
    vmeTag_array_client_id_localTag_out_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      vmeTag_array_client_id_localTag_out_MPORT_addr_pipe_0 <= io_mem_r_bits_id[3:0];
    end
    if (vmeTag_array_client_tag_rdwrPort_en & vmeTag_array_client_tag_rdwrPort_mask) begin
      vmeTag_array_client_tag[vmeTag_array_client_tag_rdwrPort_addr] <= vmeTag_array_client_tag_rdwrPort_data; // @[VME.scala 189:33]
    end
    vmeTag_array_client_tag_localTag_out_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      vmeTag_array_client_tag_localTag_out_MPORT_addr_pipe_0 <= io_mem_r_bits_id[3:0];
    end
    if (reset) begin // @[VME.scala 208:21]
      availableEntries <= 16'hffff; // @[VME.scala 209:20]
    end else if (io_mem_r_bits_last & io_mem_r_valid) begin // @[VME.scala 201:44]
      availableEntries <= _availableEntriesNext_T; // @[VME.scala 202:24]
    end else if (availableEntriesEn & availableEntries != 16'h0 & ~_T) begin // @[VME.scala 203:103]
      availableEntries <= newEntry; // @[VME.scala 204:23]
    end
    if (reset) begin // @[VME.scala 297:41]
      io_vme_rd_0_data_valid_REG <= 1'h0; // @[VME.scala 297:41]
    end else begin
      io_vme_rd_0_data_valid_REG <= io_mem_r_valid; // @[VME.scala 297:41]
    end
    if (reset) begin // @[VME.scala 301:43]
      io_vme_rd_0_data_bits_data_REG <= 64'h0; // @[VME.scala 301:43]
    end else begin
      io_vme_rd_0_data_bits_data_REG <= io_mem_r_bits_data; // @[VME.scala 301:43]
    end
    if (reset) begin // @[VME.scala 297:41]
      io_vme_rd_1_data_valid_REG <= 1'h0; // @[VME.scala 297:41]
    end else begin
      io_vme_rd_1_data_valid_REG <= io_mem_r_valid; // @[VME.scala 297:41]
    end
    if (reset) begin // @[VME.scala 301:43]
      io_vme_rd_1_data_bits_data_REG <= 64'h0; // @[VME.scala 301:43]
    end else begin
      io_vme_rd_1_data_bits_data_REG <= io_mem_r_bits_data; // @[VME.scala 301:43]
    end
    if (reset) begin // @[VME.scala 302:43]
      io_vme_rd_1_data_bits_last_REG <= 1'h0; // @[VME.scala 302:43]
    end else begin
      io_vme_rd_1_data_bits_last_REG <= io_mem_r_bits_last; // @[VME.scala 302:43]
    end
    if (reset) begin // @[VME.scala 297:41]
      io_vme_rd_2_data_valid_REG <= 1'h0; // @[VME.scala 297:41]
    end else begin
      io_vme_rd_2_data_valid_REG <= io_mem_r_valid; // @[VME.scala 297:41]
    end
    if (reset) begin // @[VME.scala 301:43]
      io_vme_rd_2_data_bits_data_REG <= 64'h0; // @[VME.scala 301:43]
    end else begin
      io_vme_rd_2_data_bits_data_REG <= io_mem_r_bits_data; // @[VME.scala 301:43]
    end
    if (reset) begin // @[VME.scala 297:41]
      io_vme_rd_3_data_valid_REG <= 1'h0; // @[VME.scala 297:41]
    end else begin
      io_vme_rd_3_data_valid_REG <= io_mem_r_valid; // @[VME.scala 297:41]
    end
    if (reset) begin // @[VME.scala 301:43]
      io_vme_rd_3_data_bits_data_REG <= 64'h0; // @[VME.scala 301:43]
    end else begin
      io_vme_rd_3_data_bits_data_REG <= io_mem_r_bits_data; // @[VME.scala 301:43]
    end
    if (reset) begin // @[VME.scala 297:41]
      io_vme_rd_4_data_valid_REG <= 1'h0; // @[VME.scala 297:41]
    end else begin
      io_vme_rd_4_data_valid_REG <= io_mem_r_valid; // @[VME.scala 297:41]
    end
    if (reset) begin // @[VME.scala 301:43]
      io_vme_rd_4_data_bits_data_REG <= 64'h0; // @[VME.scala 301:43]
    end else begin
      io_vme_rd_4_data_bits_data_REG <= io_mem_r_bits_data; // @[VME.scala 301:43]
    end
    if (reset) begin // @[VME.scala 307:23]
      wr_len <= 4'h0; // @[VME.scala 307:23]
    end else if (_T_32) begin // @[VME.scala 325:31]
      wr_len <= io_vme_wr_0_cmd_bits_len; // @[VME.scala 326:12]
    end
    if (reset) begin // @[VME.scala 308:24]
      wr_addr <= 32'h0; // @[VME.scala 308:24]
    end else if (_T_32) begin // @[VME.scala 325:31]
      wr_addr <= io_vme_wr_0_cmd_bits_addr; // @[VME.scala 327:13]
    end
    if (reset) begin // @[VME.scala 310:23]
      wstate <= 2'h0; // @[VME.scala 310:23]
    end else if (2'h0 == wstate) begin // @[VME.scala 335:17]
      if (io_vme_wr_0_cmd_valid) begin // @[VME.scala 337:35]
        wstate <= 2'h1; // @[VME.scala 338:16]
      end
    end else if (2'h1 == wstate) begin // @[VME.scala 335:17]
      if (io_mem_aw_ready) begin // @[VME.scala 342:28]
        wstate <= 2'h2; // @[VME.scala 343:16]
      end
    end else if (2'h2 == wstate) begin // @[VME.scala 335:17]
      wstate <= _GEN_52;
    end else begin
      wstate <= _GEN_54;
    end
    if (reset) begin // @[VME.scala 311:23]
      wr_cnt <= 4'h0; // @[VME.scala 311:23]
    end else if (_io_vme_wr_0_cmd_ready_T) begin // @[VME.scala 329:31]
      wr_cnt <= 4'h0; // @[VME.scala 330:12]
    end else if (_T_34) begin // @[VME.scala 332:27]
      wr_cnt <= _wr_cnt_T_1; // @[VME.scala 333:12]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(io_vme_rd_0_data_ready | ~io_vme_rd_0_data_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at VME.scala:300 assert(io.vme.rd(i).data.ready || ~io.vme.rd(i).data.valid)\n"); // @[VME.scala 300:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    vmeTag_array_client_id[initvar] = _RAND_0[2:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    vmeTag_array_client_tag[initvar] = _RAND_3[20:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  vmeTag_array_client_id_localTag_out_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  vmeTag_array_client_id_localTag_out_MPORT_addr_pipe_0 = _RAND_2[3:0];
  _RAND_4 = {1{`RANDOM}};
  vmeTag_array_client_tag_localTag_out_MPORT_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  vmeTag_array_client_tag_localTag_out_MPORT_addr_pipe_0 = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  availableEntries = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  io_vme_rd_0_data_valid_REG = _RAND_7[0:0];
  _RAND_8 = {2{`RANDOM}};
  io_vme_rd_0_data_bits_data_REG = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  io_vme_rd_1_data_valid_REG = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  io_vme_rd_1_data_bits_data_REG = _RAND_10[63:0];
  _RAND_11 = {1{`RANDOM}};
  io_vme_rd_1_data_bits_last_REG = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  io_vme_rd_2_data_valid_REG = _RAND_12[0:0];
  _RAND_13 = {2{`RANDOM}};
  io_vme_rd_2_data_bits_data_REG = _RAND_13[63:0];
  _RAND_14 = {1{`RANDOM}};
  io_vme_rd_3_data_valid_REG = _RAND_14[0:0];
  _RAND_15 = {2{`RANDOM}};
  io_vme_rd_3_data_bits_data_REG = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  io_vme_rd_4_data_valid_REG = _RAND_16[0:0];
  _RAND_17 = {2{`RANDOM}};
  io_vme_rd_4_data_bits_data_REG = _RAND_17[63:0];
  _RAND_18 = {1{`RANDOM}};
  wr_len = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  wr_addr = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  wstate = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  wr_cnt = _RAND_21[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(io_vme_rd_0_data_ready | ~io_vme_rd_0_data_valid); // @[VME.scala 300:11]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[VME.scala 300:11]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[VME.scala 300:11]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[VME.scala 300:11]
    end
    //
    if (~reset) begin
      assert(1'h1); // @[VME.scala 300:11]
    end
  end
endmodule
module TwoPortMem(
  input          clock,
  input          io_wr_en,
  input  [15:0]  io_wr_addr,
  input  [127:0] io_wr_data,
  input          io_rd_en,
  input  [15:0]  io_rd_addr,
  output [127:0] io_rd_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] mem [0:7]; // @[SyncQueue.scala 496:24]
  wire  mem_io_rd_data_MPORT_en; // @[SyncQueue.scala 496:24]
  wire [2:0] mem_io_rd_data_MPORT_addr; // @[SyncQueue.scala 496:24]
  wire [127:0] mem_io_rd_data_MPORT_data; // @[SyncQueue.scala 496:24]
  wire [127:0] mem_MPORT_data; // @[SyncQueue.scala 496:24]
  wire [2:0] mem_MPORT_addr; // @[SyncQueue.scala 496:24]
  wire  mem_MPORT_mask; // @[SyncQueue.scala 496:24]
  wire  mem_MPORT_en; // @[SyncQueue.scala 496:24]
  reg  mem_io_rd_data_MPORT_en_pipe_0;
  reg [2:0] mem_io_rd_data_MPORT_addr_pipe_0;
  assign mem_io_rd_data_MPORT_en = mem_io_rd_data_MPORT_en_pipe_0;
  assign mem_io_rd_data_MPORT_addr = mem_io_rd_data_MPORT_addr_pipe_0;
  assign mem_io_rd_data_MPORT_data = mem[mem_io_rd_data_MPORT_addr]; // @[SyncQueue.scala 496:24]
  assign mem_MPORT_data = io_wr_data;
  assign mem_MPORT_addr = io_wr_addr[2:0];
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wr_en;
  assign io_rd_data = mem_io_rd_data_MPORT_data; // @[SyncQueue.scala 502:20 503:16]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SyncQueue.scala 496:24]
    end
    mem_io_rd_data_MPORT_en_pipe_0 <= io_rd_en;
    if (io_rd_en) begin
      mem_io_rd_data_MPORT_addr_pipe_0 <= io_rd_addr[2:0];
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    mem[initvar] = _RAND_0[127:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_rd_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_rd_data_MPORT_addr_pipe_0 = _RAND_2[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module OneCycleQueue(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [127:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [127:0] io_deq_bits,
  output [3:0]   io_count
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ram0_clock; // @[SyncQueue.scala 377:20]
  wire  ram0_io_wr_en; // @[SyncQueue.scala 377:20]
  wire [15:0] ram0_io_wr_addr; // @[SyncQueue.scala 377:20]
  wire [127:0] ram0_io_wr_data; // @[SyncQueue.scala 377:20]
  wire  ram0_io_rd_en; // @[SyncQueue.scala 377:20]
  wire [15:0] ram0_io_rd_addr; // @[SyncQueue.scala 377:20]
  wire [127:0] ram0_io_rd_data; // @[SyncQueue.scala 377:20]
  reg [2:0] value; // @[Counter.scala 62:40]
  reg [2:0] value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[SyncQueue.scala 380:27]
  wire  ptr_match = value == value_1; // @[SyncQueue.scala 383:33]
  wire  empty = ptr_match & ~maybe_full; // @[SyncQueue.scala 384:25]
  wire  full = ptr_match & maybe_full; // @[SyncQueue.scala 385:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  wrap = value_1 == 3'h7; // @[Counter.scala 74:24]
  wire [2:0] _value_T_1 = value_1 + 3'h1; // @[Counter.scala 78:24]
  wire [2:0] _value_T_3 = value + 3'h1; // @[Counter.scala 78:24]
  wire  _firstRead_T_1 = do_enq & io_count == 4'h0; // @[SyncQueue.scala 403:43]
  reg  firstRead; // @[Reg.scala 28:20]
  wire  _io_deq_valid_T_1 = ~firstRead; // @[SyncQueue.scala 404:29]
  wire [2:0] _GEN_4 = wrap ? 3'h0 : _value_T_1; // @[SyncQueue.scala 413:17 414:14 416:14]
  wire [2:0] _GEN_5 = do_deq ? _GEN_4 : value_1; // @[SyncQueue.scala 411:23 419:12]
  wire [2:0] rdAddr = firstRead ? value_1 : _GEN_5; // @[SyncQueue.scala 409:19 410:12]
  wire [2:0] ptr_diff = value - value_1; // @[SyncQueue.scala 430:32]
  wire [3:0] _io_count_T_1 = maybe_full & ptr_match ? 4'h8 : 4'h0; // @[SyncQueue.scala 432:20]
  wire [3:0] _GEN_7 = {{1'd0}, ptr_diff}; // @[SyncQueue.scala 432:62]
  TwoPortMem ram0 ( // @[SyncQueue.scala 377:20]
    .clock(ram0_clock),
    .io_wr_en(ram0_io_wr_en),
    .io_wr_addr(ram0_io_wr_addr),
    .io_wr_data(ram0_io_wr_data),
    .io_rd_en(ram0_io_rd_en),
    .io_rd_addr(ram0_io_rd_addr),
    .io_rd_data(ram0_io_rd_data)
  );
  assign io_enq_ready = ~full; // @[SyncQueue.scala 405:19]
  assign io_deq_valid = ~empty & ~firstRead; // @[SyncQueue.scala 404:26]
  assign io_deq_bits = ram0_io_rd_data; // @[SyncQueue.scala 426:15]
  assign io_count = _io_count_T_1 | _GEN_7; // @[SyncQueue.scala 432:62]
  assign ram0_clock = clock;
  assign ram0_io_wr_en = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  assign ram0_io_wr_addr = {{13'd0}, value}; // @[SyncQueue.scala 423:19]
  assign ram0_io_wr_data = io_enq_bits; // @[SyncQueue.scala 422:19]
  assign ram0_io_rd_en = do_deq | firstRead; // @[SyncQueue.scala 424:27]
  assign ram0_io_rd_addr = {{13'd0}, rdAddr}; // @[SyncQueue.scala 425:19]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 62:40]
      value <= 3'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[SyncQueue.scala 399:17]
      value <= _value_T_3; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 3'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[SyncQueue.scala 391:16]
      value_1 <= _value_T_1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[SyncQueue.scala 380:27]
      maybe_full <= 1'h0; // @[SyncQueue.scala 380:27]
    end else if (do_enq != do_deq) begin // @[SyncQueue.scala 395:27]
      maybe_full <= do_enq; // @[SyncQueue.scala 396:16]
    end
    if (reset) begin // @[Reg.scala 28:20]
      firstRead <= 1'h0; // @[Reg.scala 28:20]
    end else begin
      firstRead <= _firstRead_T_1;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_io_deq_valid_T_1 | ~do_deq)) begin
          $fwrite(32'h80000002,
            "Assertion failed: -F- Cannot have deq with first read as queue output is not valid yet\n    at SyncQueue.scala:406 assert(!firstRead || !do_deq, \"-F- Cannot have deq with first read as queue output is not valid yet\")\n"
            ); // @[SyncQueue.scala 406:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  value_1 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  firstRead = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(_io_deq_valid_T_1 | ~do_deq); // @[SyncQueue.scala 406:9]
    end
  end
endmodule
module Queue_5(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [127:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [127:0] io_deq_bits
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [127:0] _RAND_1;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] ram [0:2]; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [1:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [127:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [127:0] ram_MPORT_data; // @[Decoupled.scala 259:95]
  wire [1:0] ram_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 259:95]
  reg [1:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [1:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  wrap = enq_ptr_value == 2'h2; // @[Counter.scala 74:24]
  wire [1:0] _value_T_1 = enq_ptr_value + 2'h1; // @[Counter.scala 78:24]
  wire  wrap_1 = deq_ptr_value == 2'h2; // @[Counter.scala 74:24]
  wire [1:0] _value_T_3 = deq_ptr_value + 2'h1; // @[Counter.scala 78:24]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `else
  assign ram_io_deq_bits_MPORT_data = ram_io_deq_bits_MPORT_addr >= 2'h3 ? _RAND_1[127:0] :
    ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 2'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      if (wrap) begin // @[Counter.scala 88:20]
        enq_ptr_value <= 2'h0; // @[Counter.scala 88:28]
      end else begin
        enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
      end
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 2'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      if (wrap_1) begin // @[Counter.scala 88:20]
        deq_ptr_value <= 2'h0; // @[Counter.scala 88:28]
      end else begin
        deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
      end
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {4{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 3; initvar = initvar+1)
    ram[initvar] = _RAND_0[127:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  enq_ptr_value = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  deq_ptr_value = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  maybe_full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module SyncQueue2PortMemImpl(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [127:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [127:0] io_deq_bits,
  output [3:0]   io_count
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  memoryQueue_clock; // @[SyncQueue.scala 172:27]
  wire  memoryQueue_reset; // @[SyncQueue.scala 172:27]
  wire  memoryQueue_io_enq_ready; // @[SyncQueue.scala 172:27]
  wire  memoryQueue_io_enq_valid; // @[SyncQueue.scala 172:27]
  wire [127:0] memoryQueue_io_enq_bits; // @[SyncQueue.scala 172:27]
  wire  memoryQueue_io_deq_ready; // @[SyncQueue.scala 172:27]
  wire  memoryQueue_io_deq_valid; // @[SyncQueue.scala 172:27]
  wire [127:0] memoryQueue_io_deq_bits; // @[SyncQueue.scala 172:27]
  wire [3:0] memoryQueue_io_count; // @[SyncQueue.scala 172:27]
  wire  buffer_clock; // @[SyncQueue.scala 173:22]
  wire  buffer_reset; // @[SyncQueue.scala 173:22]
  wire  buffer_io_enq_ready; // @[SyncQueue.scala 173:22]
  wire  buffer_io_enq_valid; // @[SyncQueue.scala 173:22]
  wire [127:0] buffer_io_enq_bits; // @[SyncQueue.scala 173:22]
  wire  buffer_io_deq_ready; // @[SyncQueue.scala 173:22]
  wire  buffer_io_deq_valid; // @[SyncQueue.scala 173:22]
  wire [127:0] buffer_io_deq_bits; // @[SyncQueue.scala 173:22]
  wire  memoryQueueHasValues = memoryQueue_io_count != 4'h0; // @[SyncQueue.scala 175:51]
  wire  _memoryQueue_io_enq_valid_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _countNext_T_1 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _countNext_T_2 = _memoryQueue_io_enq_valid_T | _countNext_T_1; // @[SyncQueue.scala 190:26]
  reg [3:0] countNext; // @[Reg.scala 28:20]
  wire  _T_3 = _memoryQueue_io_enq_valid_T & ~_countNext_T_1; // @[SyncQueue.scala 191:21]
  wire [3:0] _count_T_1 = countNext + 4'h1; // @[SyncQueue.scala 193:24]
  wire  _T_11 = ~_memoryQueue_io_enq_valid_T & _countNext_T_1; // @[SyncQueue.scala 194:28]
  wire [3:0] _count_T_3 = countNext - 4'h1; // @[SyncQueue.scala 196:24]
  wire  _T_6 = ~reset; // @[SyncQueue.scala 192:11]
  OneCycleQueue memoryQueue ( // @[SyncQueue.scala 172:27]
    .clock(memoryQueue_clock),
    .reset(memoryQueue_reset),
    .io_enq_ready(memoryQueue_io_enq_ready),
    .io_enq_valid(memoryQueue_io_enq_valid),
    .io_enq_bits(memoryQueue_io_enq_bits),
    .io_deq_ready(memoryQueue_io_deq_ready),
    .io_deq_valid(memoryQueue_io_deq_valid),
    .io_deq_bits(memoryQueue_io_deq_bits),
    .io_count(memoryQueue_io_count)
  );
  Queue_5 buffer ( // @[SyncQueue.scala 173:22]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .io_enq_ready(buffer_io_enq_ready),
    .io_enq_valid(buffer_io_enq_valid),
    .io_enq_bits(buffer_io_enq_bits),
    .io_deq_ready(buffer_io_deq_ready),
    .io_deq_valid(buffer_io_deq_valid),
    .io_deq_bits(buffer_io_deq_bits)
  );
  assign io_enq_ready = countNext != 4'h8; // @[SyncQueue.scala 202:30]
  assign io_deq_valid = countNext != 4'h0; // @[SyncQueue.scala 203:30]
  assign io_deq_bits = buffer_io_deq_bits; // @[SyncQueue.scala 181:10]
  assign io_count = countNext; // @[SyncQueue.scala 201:12]
  assign memoryQueue_clock = clock;
  assign memoryQueue_reset = reset;
  assign memoryQueue_io_enq_valid = _memoryQueue_io_enq_valid_T & (~buffer_io_enq_ready | memoryQueueHasValues); // @[SyncQueue.scala 183:43]
  assign memoryQueue_io_enq_bits = io_enq_bits; // @[SyncQueue.scala 182:27]
  assign memoryQueue_io_deq_ready = buffer_io_enq_ready; // @[SyncQueue.scala 184:28]
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_io_enq_valid = memoryQueueHasValues ? memoryQueue_io_deq_valid : io_enq_valid; // @[SyncQueue.scala 176:26]
  assign buffer_io_enq_bits = memoryQueueHasValues ? memoryQueue_io_deq_bits : io_enq_bits; // @[SyncQueue.scala 177:25]
  assign buffer_io_deq_ready = io_deq_ready; // @[SyncQueue.scala 181:10]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      countNext <= 4'h0; // @[Reg.scala 28:20]
    end else if (_countNext_T_2) begin // @[Reg.scala 29:18]
      if (_memoryQueue_io_enq_valid_T & ~_countNext_T_1) begin // @[SyncQueue.scala 191:38]
        countNext <= _count_T_1; // @[SyncQueue.scala 193:11]
      end else if (~_memoryQueue_io_enq_valid_T & _countNext_T_1) begin // @[SyncQueue.scala 194:44]
        countNext <= _count_T_3; // @[SyncQueue.scala 196:11]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~reset & ~(countNext < 4'h8)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at SyncQueue.scala:192 assert(countNext < entries.U)\n"); // @[SyncQueue.scala 192:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_3 & _T_11 & _T_6 & ~(countNext > 4'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at SyncQueue.scala:195 assert(countNext > 0.U)\n"); // @[SyncQueue.scala 195:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6 & ~(io_deq_valid == buffer_io_deq_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at SyncQueue.scala:204 assert(io.deq.valid === buffer.io.deq.valid)\n"); // @[SyncQueue.scala 204:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6 & ~(io_enq_ready == buffer_io_enq_ready | memoryQueue_io_enq_ready)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at SyncQueue.scala:205 assert(io.enq.ready === buffer.io.enq.ready || memoryQueue.io.enq.ready)\n"
            ); // @[SyncQueue.scala 205:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  countNext = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_3 & ~reset) begin
      assert(countNext < 4'h8); // @[SyncQueue.scala 192:11]
    end
    //
    if (~_T_3 & _T_11 & _T_6) begin
      assert(countNext > 4'h0); // @[SyncQueue.scala 195:11]
    end
    //
    if (_T_6) begin
      assert(io_deq_valid == buffer_io_deq_valid); // @[SyncQueue.scala 204:9]
    end
    //
    if (_T_6) begin
      assert(io_enq_ready == buffer_io_enq_ready | memoryQueue_io_enq_ready); // @[SyncQueue.scala 205:9]
    end
  end
endmodule
module SyncQueue2PortMem(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [127:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [127:0] io_deq_bits,
  output [3:0]   io_count
);
  wire  queue_clock; // @[SyncQueue.scala 151:23]
  wire  queue_reset; // @[SyncQueue.scala 151:23]
  wire  queue_io_enq_ready; // @[SyncQueue.scala 151:23]
  wire  queue_io_enq_valid; // @[SyncQueue.scala 151:23]
  wire [127:0] queue_io_enq_bits; // @[SyncQueue.scala 151:23]
  wire  queue_io_deq_ready; // @[SyncQueue.scala 151:23]
  wire  queue_io_deq_valid; // @[SyncQueue.scala 151:23]
  wire [127:0] queue_io_deq_bits; // @[SyncQueue.scala 151:23]
  wire [3:0] queue_io_count; // @[SyncQueue.scala 151:23]
  SyncQueue2PortMemImpl queue ( // @[SyncQueue.scala 151:23]
    .clock(queue_clock),
    .reset(queue_reset),
    .io_enq_ready(queue_io_enq_ready),
    .io_enq_valid(queue_io_enq_valid),
    .io_enq_bits(queue_io_enq_bits),
    .io_deq_ready(queue_io_deq_ready),
    .io_deq_valid(queue_io_deq_valid),
    .io_deq_bits(queue_io_deq_bits),
    .io_count(queue_io_count)
  );
  assign io_enq_ready = queue_io_enq_ready; // @[SyncQueue.scala 152:8]
  assign io_deq_valid = queue_io_deq_valid; // @[SyncQueue.scala 152:8]
  assign io_deq_bits = queue_io_deq_bits; // @[SyncQueue.scala 152:8]
  assign io_count = queue_io_count; // @[SyncQueue.scala 152:8]
  assign queue_clock = clock;
  assign queue_reset = reset;
  assign queue_io_enq_valid = io_enq_valid; // @[SyncQueue.scala 152:8]
  assign queue_io_enq_bits = io_enq_bits; // @[SyncQueue.scala 152:8]
  assign queue_io_deq_ready = io_deq_ready; // @[SyncQueue.scala 152:8]
endmodule
module SyncQueue(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [127:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [127:0] io_deq_bits,
  output [3:0]   io_count
);
  wire  queue_clock; // @[SyncQueue.scala 47:23]
  wire  queue_reset; // @[SyncQueue.scala 47:23]
  wire  queue_io_enq_ready; // @[SyncQueue.scala 47:23]
  wire  queue_io_enq_valid; // @[SyncQueue.scala 47:23]
  wire [127:0] queue_io_enq_bits; // @[SyncQueue.scala 47:23]
  wire  queue_io_deq_ready; // @[SyncQueue.scala 47:23]
  wire  queue_io_deq_valid; // @[SyncQueue.scala 47:23]
  wire [127:0] queue_io_deq_bits; // @[SyncQueue.scala 47:23]
  wire [3:0] queue_io_count; // @[SyncQueue.scala 47:23]
  SyncQueue2PortMem queue ( // @[SyncQueue.scala 47:23]
    .clock(queue_clock),
    .reset(queue_reset),
    .io_enq_ready(queue_io_enq_ready),
    .io_enq_valid(queue_io_enq_valid),
    .io_enq_bits(queue_io_enq_bits),
    .io_deq_ready(queue_io_deq_ready),
    .io_deq_valid(queue_io_deq_valid),
    .io_deq_bits(queue_io_deq_bits),
    .io_count(queue_io_count)
  );
  assign io_enq_ready = queue_io_enq_ready; // @[SyncQueue.scala 48:8]
  assign io_deq_valid = queue_io_deq_valid; // @[SyncQueue.scala 48:8]
  assign io_deq_bits = queue_io_deq_bits; // @[SyncQueue.scala 48:8]
  assign io_count = queue_io_count; // @[SyncQueue.scala 48:8]
  assign queue_clock = clock;
  assign queue_reset = reset;
  assign queue_io_enq_valid = io_enq_valid; // @[SyncQueue.scala 48:8]
  assign queue_io_enq_bits = io_enq_bits; // @[SyncQueue.scala 48:8]
  assign queue_io_deq_ready = io_deq_ready; // @[SyncQueue.scala 48:8]
endmodule
module FetchDecode(
  input  [127:0] io_inst,
  output         io_isLoad,
  output         io_isCompute,
  output         io_isStore
);
  wire [127:0] _csignals_T = io_inst & 128'h387; // @[Lookup.scala 31:38]
  wire  _csignals_T_1 = 128'h0 == _csignals_T; // @[Lookup.scala 31:38]
  wire  _csignals_T_3 = 128'h80 == _csignals_T; // @[Lookup.scala 31:38]
  wire  _csignals_T_5 = 128'h100 == _csignals_T; // @[Lookup.scala 31:38]
  wire  _csignals_T_7 = 128'h180 == _csignals_T; // @[Lookup.scala 31:38]
  wire [127:0] _csignals_T_8 = io_inst & 128'h7; // @[Lookup.scala 31:38]
  wire  _csignals_T_9 = 128'h1 == _csignals_T_8; // @[Lookup.scala 31:38]
  wire  _csignals_T_11 = 128'h2 == _csignals_T_8; // @[Lookup.scala 31:38]
  wire  _csignals_T_13 = 128'h3 == _csignals_T_8; // @[Lookup.scala 31:38]
  wire [127:0] _csignals_T_14 = io_inst & 128'h7000000000000000000000000007; // @[Lookup.scala 31:38]
  wire  _csignals_T_15 = 128'h4 == _csignals_T_14; // @[Lookup.scala 31:38]
  wire  _csignals_T_17 = 128'h1000000000000000000000000004 == _csignals_T_14; // @[Lookup.scala 31:38]
  wire  _csignals_T_19 = 128'h2000000000000000000000000004 == _csignals_T_14; // @[Lookup.scala 31:38]
  wire  _csignals_T_21 = 128'h3000000000000000000000000004 == _csignals_T_14; // @[Lookup.scala 31:38]
  wire  cs_val_inst = _csignals_T_1 | (_csignals_T_3 | (_csignals_T_5 | (_csignals_T_7 | (_csignals_T_9 | (
    _csignals_T_11 | (_csignals_T_13 | (_csignals_T_15 | (_csignals_T_17 | (_csignals_T_19 | _csignals_T_21))))))))); // @[Lookup.scala 34:39]
  wire [2:0] _csignals_T_32 = _csignals_T_21 ? 3'h2 : 3'h5; // @[Lookup.scala 34:39]
  wire [2:0] _csignals_T_33 = _csignals_T_19 ? 3'h2 : _csignals_T_32; // @[Lookup.scala 34:39]
  wire [2:0] _csignals_T_34 = _csignals_T_17 ? 3'h2 : _csignals_T_33; // @[Lookup.scala 34:39]
  wire [2:0] _csignals_T_35 = _csignals_T_15 ? 3'h2 : _csignals_T_34; // @[Lookup.scala 34:39]
  wire [2:0] _csignals_T_36 = _csignals_T_13 ? 3'h2 : _csignals_T_35; // @[Lookup.scala 34:39]
  wire [2:0] _csignals_T_37 = _csignals_T_11 ? 3'h2 : _csignals_T_36; // @[Lookup.scala 34:39]
  wire [2:0] _csignals_T_38 = _csignals_T_9 ? 3'h1 : _csignals_T_37; // @[Lookup.scala 34:39]
  wire [2:0] _csignals_T_39 = _csignals_T_7 ? 3'h2 : _csignals_T_38; // @[Lookup.scala 34:39]
  wire [2:0] _csignals_T_40 = _csignals_T_5 ? 3'h0 : _csignals_T_39; // @[Lookup.scala 34:39]
  wire [2:0] _csignals_T_41 = _csignals_T_3 ? 3'h0 : _csignals_T_40; // @[Lookup.scala 34:39]
  wire [2:0] cs_op_type = _csignals_T_1 ? 3'h2 : _csignals_T_41; // @[Lookup.scala 34:39]
  assign io_isLoad = cs_val_inst & cs_op_type == 3'h0; // @[Decode.scala 155:28]
  assign io_isCompute = cs_val_inst & cs_op_type == 3'h2; // @[Decode.scala 156:31]
  assign io_isStore = cs_val_inst & cs_op_type == 3'h1; // @[Decode.scala 157:29]
endmodule
module Fetch64Bit(
  input          clock,
  input          reset,
  input          io_launch,
  input  [31:0]  io_ins_baddr,
  input  [31:0]  io_ins_count,
  input          io_vme_rd_cmd_ready,
  output         io_vme_rd_cmd_valid,
  output [31:0]  io_vme_rd_cmd_bits_addr,
  output [3:0]   io_vme_rd_cmd_bits_len,
  output         io_vme_rd_data_ready,
  input          io_vme_rd_data_valid,
  input  [63:0]  io_vme_rd_data_bits_data,
  input          io_inst_ld_ready,
  output         io_inst_ld_valid,
  output [127:0] io_inst_ld_bits,
  input          io_inst_co_ready,
  output         io_inst_co_valid,
  output [127:0] io_inst_co_bits,
  input          io_inst_st_ready,
  output         io_inst_st_valid,
  output [127:0] io_inst_st_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  inst_q_clock; // @[FetchVME64.scala 58:22]
  wire  inst_q_reset; // @[FetchVME64.scala 58:22]
  wire  inst_q_io_enq_ready; // @[FetchVME64.scala 58:22]
  wire  inst_q_io_enq_valid; // @[FetchVME64.scala 58:22]
  wire [127:0] inst_q_io_enq_bits; // @[FetchVME64.scala 58:22]
  wire  inst_q_io_deq_ready; // @[FetchVME64.scala 58:22]
  wire  inst_q_io_deq_valid; // @[FetchVME64.scala 58:22]
  wire [127:0] inst_q_io_deq_bits; // @[FetchVME64.scala 58:22]
  wire [3:0] inst_q_io_count; // @[FetchVME64.scala 58:22]
  wire [127:0] dec_io_inst; // @[FetchVME64.scala 59:19]
  wire  dec_io_isLoad; // @[FetchVME64.scala 59:19]
  wire  dec_io_isCompute; // @[FetchVME64.scala 59:19]
  wire  dec_io_isStore; // @[FetchVME64.scala 59:19]
  reg  s1_launch; // @[FetchVME64.scala 61:26]
  wire  pulse = io_launch & ~s1_launch; // @[FetchVME64.scala 62:25]
  reg [31:0] raddr; // @[FetchVME64.scala 64:18]
  reg [3:0] rlen; // @[FetchVME64.scala 65:17]
  reg [3:0] ilen; // @[FetchVME64.scala 66:17]
  reg [31:0] xrem; // @[FetchVME64.scala 68:17]
  wire [32:0] _xsize_T = {io_ins_count, 1'h0}; // @[FetchVME64.scala 69:29]
  wire [32:0] xsize = _xsize_T - 33'h1; // @[FetchVME64.scala 69:37]
  reg [2:0] state; // @[FetchVME64.scala 74:22]
  wire [32:0] _ilen_T = {{1'd0}, xsize[32:1]}; // @[FetchVME64.scala 83:25]
  wire [4:0] _rlen_T_1 = 5'h10 - 5'h1; // @[FetchVME64.scala 86:24]
  wire [4:0] _ilen_T_3 = 5'h8 - 5'h1; // @[FetchVME64.scala 87:33]
  wire [32:0] _xrem_T_1 = xsize - 33'h10; // @[FetchVME64.scala 88:25]
  wire [32:0] _GEN_0 = xsize < 33'h10 ? xsize : {{28'd0}, _rlen_T_1}; // @[FetchVME64.scala 81:28 82:16 86:16]
  wire [32:0] _GEN_1 = xsize < 33'h10 ? _ilen_T : {{28'd0}, _ilen_T_3}; // @[FetchVME64.scala 81:28 83:16 87:16]
  wire [32:0] _GEN_2 = xsize < 33'h10 ? 33'h0 : _xrem_T_1; // @[FetchVME64.scala 81:28 84:16 88:16]
  wire [32:0] _GEN_4 = pulse ? _GEN_0 : {{29'd0}, rlen}; // @[FetchVME64.scala 65:17 79:19]
  wire [32:0] _GEN_5 = pulse ? _GEN_1 : {{29'd0}, ilen}; // @[FetchVME64.scala 66:17 79:19]
  wire [32:0] _GEN_6 = pulse ? _GEN_2 : {{1'd0}, xrem}; // @[FetchVME64.scala 68:17 79:19]
  wire [2:0] _GEN_8 = io_vme_rd_data_valid ? 3'h3 : state; // @[FetchVME64.scala 98:34 99:15 74:22]
  wire [2:0] _GEN_9 = inst_q_io_count == ilen ? 3'h4 : 3'h2; // @[FetchVME64.scala 104:40 105:17 107:17]
  wire [2:0] _GEN_10 = io_vme_rd_data_valid ? _GEN_9 : state; // @[FetchVME64.scala 103:34 74:22]
  wire  _T_7 = inst_q_io_count == 4'h0; // @[FetchVME64.scala 112:28]
  wire [31:0] _ilen_T_4 = {{1'd0}, xrem[31:1]}; // @[FetchVME64.scala 118:24]
  wire [31:0] _xrem_T_3 = xrem - 32'h10; // @[FetchVME64.scala 124:24]
  wire [31:0] _GEN_12 = xrem < 32'h10 ? xrem : {{27'd0}, _rlen_T_1}; // @[FetchVME64.scala 115:33 117:16 122:16]
  wire [31:0] _GEN_13 = xrem < 32'h10 ? _ilen_T_4 : {{27'd0}, _ilen_T_3}; // @[FetchVME64.scala 115:33 118:16 123:16]
  wire [31:0] _GEN_14 = xrem < 32'h10 ? 32'h0 : _xrem_T_3; // @[FetchVME64.scala 115:33 119:16 124:16]
  wire [2:0] _GEN_15 = xrem == 32'h0 ? 3'h0 : 3'h1; // @[FetchVME64.scala 113:28 114:17]
  wire [31:0] _GEN_16 = xrem == 32'h0 ? {{28'd0}, rlen} : _GEN_12; // @[FetchVME64.scala 113:28 65:17]
  wire [31:0] _GEN_17 = xrem == 32'h0 ? {{28'd0}, ilen} : _GEN_13; // @[FetchVME64.scala 113:28 66:17]
  wire [31:0] _GEN_18 = xrem == 32'h0 ? xrem : _GEN_14; // @[FetchVME64.scala 113:28 68:17]
  wire [2:0] _GEN_19 = inst_q_io_count == 4'h0 ? _GEN_15 : state; // @[FetchVME64.scala 112:37 74:22]
  wire [31:0] _GEN_20 = inst_q_io_count == 4'h0 ? _GEN_16 : {{28'd0}, rlen}; // @[FetchVME64.scala 112:37 65:17]
  wire [31:0] _GEN_21 = inst_q_io_count == 4'h0 ? _GEN_17 : {{28'd0}, ilen}; // @[FetchVME64.scala 112:37 66:17]
  wire [31:0] _GEN_22 = inst_q_io_count == 4'h0 ? _GEN_18 : xrem; // @[FetchVME64.scala 112:37 68:17]
  wire [2:0] _GEN_23 = 3'h4 == state ? _GEN_19 : state; // @[FetchVME64.scala 77:17 74:22]
  wire [31:0] _GEN_24 = 3'h4 == state ? _GEN_20 : {{28'd0}, rlen}; // @[FetchVME64.scala 65:17 77:17]
  wire [31:0] _GEN_25 = 3'h4 == state ? _GEN_21 : {{28'd0}, ilen}; // @[FetchVME64.scala 66:17 77:17]
  wire [31:0] _GEN_26 = 3'h4 == state ? _GEN_22 : xrem; // @[FetchVME64.scala 68:17 77:17]
  wire [2:0] _GEN_27 = 3'h3 == state ? _GEN_10 : _GEN_23; // @[FetchVME64.scala 77:17]
  wire [31:0] _GEN_28 = 3'h3 == state ? {{28'd0}, rlen} : _GEN_24; // @[FetchVME64.scala 65:17 77:17]
  wire [31:0] _GEN_29 = 3'h3 == state ? {{28'd0}, ilen} : _GEN_25; // @[FetchVME64.scala 66:17 77:17]
  wire [31:0] _GEN_30 = 3'h3 == state ? xrem : _GEN_26; // @[FetchVME64.scala 68:17 77:17]
  wire [31:0] _GEN_32 = 3'h2 == state ? {{28'd0}, rlen} : _GEN_28; // @[FetchVME64.scala 65:17 77:17]
  wire [31:0] _GEN_33 = 3'h2 == state ? {{28'd0}, ilen} : _GEN_29; // @[FetchVME64.scala 66:17 77:17]
  wire [31:0] _GEN_34 = 3'h2 == state ? xrem : _GEN_30; // @[FetchVME64.scala 68:17 77:17]
  wire [31:0] _GEN_36 = 3'h1 == state ? {{28'd0}, rlen} : _GEN_32; // @[FetchVME64.scala 65:17 77:17]
  wire [31:0] _GEN_37 = 3'h1 == state ? {{28'd0}, ilen} : _GEN_33; // @[FetchVME64.scala 66:17 77:17]
  wire [31:0] _GEN_38 = 3'h1 == state ? xrem : _GEN_34; // @[FetchVME64.scala 68:17 77:17]
  wire [32:0] _GEN_40 = 3'h0 == state ? _GEN_4 : {{1'd0}, _GEN_36}; // @[FetchVME64.scala 77:17]
  wire [32:0] _GEN_41 = 3'h0 == state ? _GEN_5 : {{1'd0}, _GEN_37}; // @[FetchVME64.scala 77:17]
  wire [32:0] _GEN_42 = 3'h0 == state ? _GEN_6 : {{1'd0}, _GEN_38}; // @[FetchVME64.scala 77:17]
  wire  _T_11 = state == 3'h4; // @[FetchVME64.scala 133:20]
  wire [31:0] _raddr_T_1 = raddr + 32'h80; // @[FetchVME64.scala 134:20]
  reg [63:0] lsb; // @[FetchVME64.scala 144:16]
  wire [2:0] deq_sel = {dec_io_isCompute,dec_io_isStore,dec_io_isLoad}; // @[Cat.scala 31:58]
  wire  _deq_ready_T_3 = 3'h2 == deq_sel ? io_inst_st_ready : 3'h1 == deq_sel & io_inst_ld_ready; // @[Mux.scala 81:58]
  wire  deq_ready = 3'h4 == deq_sel ? io_inst_co_ready : _deq_ready_T_3; // @[Mux.scala 81:58]
  SyncQueue inst_q ( // @[FetchVME64.scala 58:22]
    .clock(inst_q_clock),
    .reset(inst_q_reset),
    .io_enq_ready(inst_q_io_enq_ready),
    .io_enq_valid(inst_q_io_enq_valid),
    .io_enq_bits(inst_q_io_enq_bits),
    .io_deq_ready(inst_q_io_deq_ready),
    .io_deq_valid(inst_q_io_deq_valid),
    .io_deq_bits(inst_q_io_deq_bits),
    .io_count(inst_q_io_count)
  );
  FetchDecode dec ( // @[FetchVME64.scala 59:19]
    .io_inst(dec_io_inst),
    .io_isLoad(dec_io_isLoad),
    .io_isCompute(dec_io_isCompute),
    .io_isStore(dec_io_isStore)
  );
  assign io_vme_rd_cmd_valid = state == 3'h1; // @[FetchVME64.scala 137:32]
  assign io_vme_rd_cmd_bits_addr = raddr; // @[FetchVME64.scala 138:27]
  assign io_vme_rd_cmd_bits_len = rlen; // @[FetchVME64.scala 139:26]
  assign io_vme_rd_data_ready = inst_q_io_enq_ready; // @[FetchVME64.scala 142:24]
  assign io_inst_ld_valid = dec_io_isLoad & inst_q_io_deq_valid & _T_11; // @[FetchVME64.scala 157:59]
  assign io_inst_ld_bits = inst_q_io_deq_bits; // @[FetchVME64.scala 164:19]
  assign io_inst_co_valid = dec_io_isCompute & inst_q_io_deq_valid & _T_11; // @[FetchVME64.scala 158:62]
  assign io_inst_co_bits = inst_q_io_deq_bits; // @[FetchVME64.scala 165:19]
  assign io_inst_st_valid = dec_io_isStore & inst_q_io_deq_valid & _T_11; // @[FetchVME64.scala 159:60]
  assign io_inst_st_bits = inst_q_io_deq_bits; // @[FetchVME64.scala 166:19]
  assign inst_q_clock = clock;
  assign inst_q_reset = reset;
  assign inst_q_io_enq_valid = io_vme_rd_data_valid & state == 3'h3; // @[FetchVME64.scala 150:47]
  assign inst_q_io_enq_bits = {io_vme_rd_data_bits_data,lsb}; // @[Cat.scala 31:58]
  assign inst_q_io_deq_ready = deq_ready & inst_q_io_deq_valid & _T_11; // @[FetchVME64.scala 180:58]
  assign dec_io_inst = inst_q_io_deq_bits; // @[FetchVME64.scala 154:15]
  always @(posedge clock) begin
    if (reset) begin // @[FetchVME64.scala 61:26]
      s1_launch <= 1'h0; // @[FetchVME64.scala 61:26]
    end else begin
      s1_launch <= io_launch; // @[FetchVME64.scala 61:26]
    end
    if (state == 3'h0) begin // @[FetchVME64.scala 131:25]
      raddr <= io_ins_baddr; // @[FetchVME64.scala 132:11]
    end else if (state == 3'h4 & _T_7 & xrem != 32'h0) begin // @[FetchVME64.scala 133:75]
      raddr <= _raddr_T_1; // @[FetchVME64.scala 134:11]
    end
    rlen <= _GEN_40[3:0];
    ilen <= _GEN_41[3:0];
    xrem <= _GEN_42[31:0];
    if (reset) begin // @[FetchVME64.scala 74:22]
      state <= 3'h0; // @[FetchVME64.scala 74:22]
    end else if (3'h0 == state) begin // @[FetchVME64.scala 77:17]
      if (pulse) begin // @[FetchVME64.scala 79:19]
        state <= 3'h1; // @[FetchVME64.scala 80:15]
      end
    end else if (3'h1 == state) begin // @[FetchVME64.scala 77:17]
      if (io_vme_rd_cmd_ready) begin // @[FetchVME64.scala 93:33]
        state <= 3'h2; // @[FetchVME64.scala 94:15]
      end
    end else if (3'h2 == state) begin // @[FetchVME64.scala 77:17]
      state <= _GEN_8;
    end else begin
      state <= _GEN_27;
    end
    if (state == 3'h2) begin // @[FetchVME64.scala 148:28]
      lsb <= io_vme_rd_data_bits_data; // @[FetchVME64.scala 148:34]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~(inst_q_io_deq_valid & _T_11) | dec_io_isLoad | dec_io_isCompute | dec_io_isStore)) begin
          $fwrite(32'h80000002,
            "Assertion failed: -F- Fetch: Unknown instruction type\n    at FetchVME64.scala:161 assert(!(inst_q.io.deq.valid & state === sDrain) || dec.io.isLoad || dec.io.isCompute || dec.io.isStore,\n"
            ); // @[FetchVME64.scala 161:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  s1_launch = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  raddr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  rlen = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  ilen = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  xrem = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  state = _RAND_5[2:0];
  _RAND_6 = {2{`RANDOM}};
  lsb = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~(inst_q_io_deq_valid & _T_11) | dec_io_isLoad | dec_io_isCompute | dec_io_isStore); // @[FetchVME64.scala 161:9]
    end
  end
endmodule
module Fetch(
  input          clock,
  input          reset,
  input          io_launch,
  input  [31:0]  io_ins_baddr,
  input  [31:0]  io_ins_count,
  input          io_vme_rd_cmd_ready,
  output         io_vme_rd_cmd_valid,
  output [31:0]  io_vme_rd_cmd_bits_addr,
  output [3:0]   io_vme_rd_cmd_bits_len,
  output         io_vme_rd_data_ready,
  input          io_vme_rd_data_valid,
  input  [63:0]  io_vme_rd_data_bits_data,
  input          io_inst_ld_ready,
  output         io_inst_ld_valid,
  output [127:0] io_inst_ld_bits,
  input          io_inst_co_ready,
  output         io_inst_co_valid,
  output [127:0] io_inst_co_bits,
  input          io_inst_st_ready,
  output         io_inst_st_valid,
  output [127:0] io_inst_st_bits
);
  wire  fetch_clock; // @[Fetch.scala 70:23]
  wire  fetch_reset; // @[Fetch.scala 70:23]
  wire  fetch_io_launch; // @[Fetch.scala 70:23]
  wire [31:0] fetch_io_ins_baddr; // @[Fetch.scala 70:23]
  wire [31:0] fetch_io_ins_count; // @[Fetch.scala 70:23]
  wire  fetch_io_vme_rd_cmd_ready; // @[Fetch.scala 70:23]
  wire  fetch_io_vme_rd_cmd_valid; // @[Fetch.scala 70:23]
  wire [31:0] fetch_io_vme_rd_cmd_bits_addr; // @[Fetch.scala 70:23]
  wire [3:0] fetch_io_vme_rd_cmd_bits_len; // @[Fetch.scala 70:23]
  wire  fetch_io_vme_rd_data_ready; // @[Fetch.scala 70:23]
  wire  fetch_io_vme_rd_data_valid; // @[Fetch.scala 70:23]
  wire [63:0] fetch_io_vme_rd_data_bits_data; // @[Fetch.scala 70:23]
  wire  fetch_io_inst_ld_ready; // @[Fetch.scala 70:23]
  wire  fetch_io_inst_ld_valid; // @[Fetch.scala 70:23]
  wire [127:0] fetch_io_inst_ld_bits; // @[Fetch.scala 70:23]
  wire  fetch_io_inst_co_ready; // @[Fetch.scala 70:23]
  wire  fetch_io_inst_co_valid; // @[Fetch.scala 70:23]
  wire [127:0] fetch_io_inst_co_bits; // @[Fetch.scala 70:23]
  wire  fetch_io_inst_st_ready; // @[Fetch.scala 70:23]
  wire  fetch_io_inst_st_valid; // @[Fetch.scala 70:23]
  wire [127:0] fetch_io_inst_st_bits; // @[Fetch.scala 70:23]
  Fetch64Bit fetch ( // @[Fetch.scala 70:23]
    .clock(fetch_clock),
    .reset(fetch_reset),
    .io_launch(fetch_io_launch),
    .io_ins_baddr(fetch_io_ins_baddr),
    .io_ins_count(fetch_io_ins_count),
    .io_vme_rd_cmd_ready(fetch_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(fetch_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(fetch_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(fetch_io_vme_rd_cmd_bits_len),
    .io_vme_rd_data_ready(fetch_io_vme_rd_data_ready),
    .io_vme_rd_data_valid(fetch_io_vme_rd_data_valid),
    .io_vme_rd_data_bits_data(fetch_io_vme_rd_data_bits_data),
    .io_inst_ld_ready(fetch_io_inst_ld_ready),
    .io_inst_ld_valid(fetch_io_inst_ld_valid),
    .io_inst_ld_bits(fetch_io_inst_ld_bits),
    .io_inst_co_ready(fetch_io_inst_co_ready),
    .io_inst_co_valid(fetch_io_inst_co_valid),
    .io_inst_co_bits(fetch_io_inst_co_bits),
    .io_inst_st_ready(fetch_io_inst_st_ready),
    .io_inst_st_valid(fetch_io_inst_st_valid),
    .io_inst_st_bits(fetch_io_inst_st_bits)
  );
  assign io_vme_rd_cmd_valid = fetch_io_vme_rd_cmd_valid; // @[Fetch.scala 71:8]
  assign io_vme_rd_cmd_bits_addr = fetch_io_vme_rd_cmd_bits_addr; // @[Fetch.scala 71:8]
  assign io_vme_rd_cmd_bits_len = fetch_io_vme_rd_cmd_bits_len; // @[Fetch.scala 71:8]
  assign io_vme_rd_data_ready = fetch_io_vme_rd_data_ready; // @[Fetch.scala 71:8]
  assign io_inst_ld_valid = fetch_io_inst_ld_valid; // @[Fetch.scala 71:8]
  assign io_inst_ld_bits = fetch_io_inst_ld_bits; // @[Fetch.scala 71:8]
  assign io_inst_co_valid = fetch_io_inst_co_valid; // @[Fetch.scala 71:8]
  assign io_inst_co_bits = fetch_io_inst_co_bits; // @[Fetch.scala 71:8]
  assign io_inst_st_valid = fetch_io_inst_st_valid; // @[Fetch.scala 71:8]
  assign io_inst_st_bits = fetch_io_inst_st_bits; // @[Fetch.scala 71:8]
  assign fetch_clock = clock;
  assign fetch_reset = reset;
  assign fetch_io_launch = io_launch; // @[Fetch.scala 71:8]
  assign fetch_io_ins_baddr = io_ins_baddr; // @[Fetch.scala 71:8]
  assign fetch_io_ins_count = io_ins_count; // @[Fetch.scala 71:8]
  assign fetch_io_vme_rd_cmd_ready = io_vme_rd_cmd_ready; // @[Fetch.scala 71:8]
  assign fetch_io_vme_rd_data_valid = io_vme_rd_data_valid; // @[Fetch.scala 71:8]
  assign fetch_io_vme_rd_data_bits_data = io_vme_rd_data_bits_data; // @[Fetch.scala 71:8]
  assign fetch_io_inst_ld_ready = io_inst_ld_ready; // @[Fetch.scala 71:8]
  assign fetch_io_inst_co_ready = io_inst_co_ready; // @[Fetch.scala 71:8]
  assign fetch_io_inst_st_ready = io_inst_st_ready; // @[Fetch.scala 71:8]
endmodule
module Semaphore(
  input   clock,
  input   reset,
  input   io_spost,
  input   io_swait,
  output  io_sready
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] cnt; // @[Semaphore.scala 38:20]
  wire [7:0] _cnt_T_1 = cnt + 8'h1; // @[Semaphore.scala 40:16]
  wire [7:0] _cnt_T_3 = cnt - 8'h1; // @[Semaphore.scala 42:59]
  assign io_sready = cnt != 8'h0; // @[Semaphore.scala 43:20]
  always @(posedge clock) begin
    if (reset) begin // @[Semaphore.scala 38:20]
      cnt <= 8'h0; // @[Semaphore.scala 38:20]
    end else if (~io_spost & io_swait & cnt != 8'h0) begin // @[Semaphore.scala 42:46]
      cnt <= _cnt_T_3; // @[Semaphore.scala 42:52]
    end else if (io_spost & ~io_swait & cnt != 8'hff) begin // @[Semaphore.scala 39:74]
      cnt <= _cnt_T_1; // @[Semaphore.scala 40:9]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue_6(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [127:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [127:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] ram [0:31]; // @[Decoupled.scala 259:95]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:95]
  wire [4:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:95]
  wire [127:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:95]
  wire [127:0] ram_MPORT_data; // @[Decoupled.scala 259:95]
  wire [4:0] ram_MPORT_addr; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_mask; // @[Decoupled.scala 259:95]
  wire  ram_MPORT_en; // @[Decoupled.scala 259:95]
  reg [4:0] enq_ptr_value; // @[Counter.scala 62:40]
  reg [4:0] deq_ptr_value; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = enq_ptr_value == deq_ptr_value; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [4:0] _value_T_1 = enq_ptr_value + 5'h1; // @[Counter.scala 78:24]
  wire [4:0] _value_T_3 = deq_ptr_value + 5'h1; // @[Counter.scala 78:24]
  assign ram_io_deq_bits_MPORT_en = 1'h1;
  assign ram_io_deq_bits_MPORT_addr = deq_ptr_value;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:95]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = enq_ptr_value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 296:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 259:95]
    end
    if (reset) begin // @[Counter.scala 62:40]
      enq_ptr_value <= 5'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      enq_ptr_value <= _value_T_1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      deq_ptr_value <= 5'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      deq_ptr_value <= _value_T_3; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    ram[initvar] = _RAND_0[127:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  enq_ptr_value = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  deq_ptr_value = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  maybe_full = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module LoadDecode(
  input  [127:0] io_inst,
  output         io_push_next,
  output         io_pop_next,
  output         io_isInput,
  output         io_isWeight,
  output         io_isSync
);
  wire [15:0] dec_xsize = io_inst[95:80]; // @[Decode.scala 173:29]
  wire [127:0] _io_isInput_T = io_inst & 128'h387; // @[Decode.scala 176:25]
  wire  _io_isInput_T_1 = 128'h100 == _io_isInput_T; // @[Decode.scala 176:25]
  wire  _io_isInput_T_2 = dec_xsize != 16'h0; // @[Decode.scala 176:46]
  wire  _io_isWeight_T_1 = 128'h80 == _io_isInput_T; // @[Decode.scala 177:26]
  assign io_push_next = io_inst[6]; // @[Decode.scala 173:29]
  assign io_pop_next = io_inst[4]; // @[Decode.scala 173:29]
  assign io_isInput = 128'h100 == _io_isInput_T & dec_xsize != 16'h0; // @[Decode.scala 176:34]
  assign io_isWeight = 128'h80 == _io_isInput_T & _io_isInput_T_2; // @[Decode.scala 177:35]
  assign io_isSync = (_io_isInput_T_1 | _io_isWeight_T_1) & dec_xsize == 16'h0; // @[Decode.scala 178:54]
endmodule
module GenVMECmd(
  input          clock,
  input          reset,
  input          io_start,
  input          io_isBusy,
  input  [127:0] io_inst,
  input  [31:0]  io_baddr,
  input          io_vmeCmd_ready,
  output         io_vmeCmd_valid,
  output [31:0]  io_vmeCmd_bits_addr,
  output [3:0]   io_vmeCmd_bits_len,
  output [20:0]  io_vmeCmd_bits_tag,
  output [4:0]   io_readLen,
  output         io_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] dec_sram_offset = io_inst[25:10]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [31:0] dec_dram_offset = io_inst[57:26]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [15:0] dec_ysize = io_inst[79:64]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [15:0] dec_xsize = io_inst[95:80]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [15:0] dec_xstride = io_inst[111:96]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [3:0] dec_ypad_0 = io_inst[115:112]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [3:0] dec_xpad_0 = io_inst[123:120]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [3:0] dec_xpad_1 = io_inst[127:124]; // @[TensorLoadNarrowVME.scala 566:29]
  reg [31:0] rdCmdExtAddr; // @[TensorLoadNarrowVME.scala 568:25]
  wire [35:0] _xfer_init_addr_T = {dec_dram_offset, 4'h0}; // @[TensorLoadNarrowVME.scala 573:66]
  wire [35:0] _xfer_init_addr_T_1 = 36'hffffffff & _xfer_init_addr_T; // @[TensorLoadNarrowVME.scala 573:47]
  wire [35:0] _GEN_31 = {{4'd0}, io_baddr}; // @[TensorLoadNarrowVME.scala 573:33]
  wire [35:0] xfer_init_addr = _GEN_31 | _xfer_init_addr_T_1; // @[TensorLoadNarrowVME.scala 573:33]
  wire [31:0] _GEN_0 = rdCmdExtAddr % 32'h80; // @[TensorLoadNarrowVME.scala 577:53]
  wire [7:0] _firstMaxTransfer_T = _GEN_0[7:0]; // @[TensorLoadNarrowVME.scala 577:53]
  wire [7:0] _firstMaxTransfer_T_2 = 8'h80 - _firstMaxTransfer_T; // @[TensorLoadNarrowVME.scala 577:38]
  wire [4:0] firstMaxTransfer = _firstMaxTransfer_T_2[7:3]; // @[TensorLoadNarrowVME.scala 577:67]
  reg [6:0] rdCmdStartIdx; // @[TensorLoadNarrowVME.scala 586:26]
  reg  commandsDone; // @[TensorLoadNarrowVME.scala 588:29]
  wire [16:0] blocksReadSize = {dec_xsize, 1'h0}; // @[TensorLoadNarrowVME.scala 590:35]
  reg [16:0] blocksReadNb; // @[TensorLoadNarrowVME.scala 591:25]
  reg [31:0] rdCmdExtAddrRowBegin; // @[TensorLoadNarrowVME.scala 592:33]
  reg  newReadRow; // @[TensorLoadNarrowVME.scala 593:23]
  reg [15:0] srcRowIdx; // @[TensorLoadNarrowVME.scala 596:22]
  wire [15:0] _srcRowIdx_T_1 = srcRowIdx + 16'h1; // @[TensorLoadNarrowVME.scala 600:28]
  wire [16:0] blocksRemained = blocksReadSize - blocksReadNb; // @[TensorLoadNarrowVME.scala 628:39]
  wire [16:0] _GEN_32 = {{12'd0}, firstMaxTransfer}; // @[TensorLoadNarrowVME.scala 630:25]
  wire [16:0] _GEN_8 = blocksRemained < _GEN_32 ? blocksRemained : {{12'd0}, firstMaxTransfer}; // @[TensorLoadNarrowVME.scala 630:45 631:15 633:15]
  wire [16:0] _GEN_9 = blocksRemained < 17'h10 ? blocksRemained : 17'h10; // @[TensorLoadNarrowVME.scala 636:40 637:15 639:15]
  wire [16:0] _GEN_10 = newReadRow ? _GEN_8 : _GEN_9; // @[TensorLoadNarrowVME.scala 629:21]
  wire [4:0] readLen = _GEN_10[4:0]; // @[TensorLoadNarrowVME.scala 587:21]
  wire [16:0] _GEN_33 = {{12'd0}, readLen}; // @[TensorLoadNarrowVME.scala 621:41]
  wire [16:0] _T_8 = blocksReadSize - _GEN_33; // @[TensorLoadNarrowVME.scala 621:41]
  wire [15:0] _T_11 = dec_ysize - 16'h1; // @[TensorLoadNarrowVME.scala 621:80]
  wire  _T_14 = io_vmeCmd_ready & io_vmeCmd_valid; // @[Decoupled.scala 50:35]
  wire  stride = blocksReadNb == _T_8 & srcRowIdx != _T_11 & _T_14; // @[TensorLoadNarrowVME.scala 621:87]
  wire [16:0] nextBlRNb = blocksReadNb + _GEN_33; // @[TensorLoadNarrowVME.scala 611:34]
  wire  _GEN_2 = nextBlRNb == blocksReadSize & srcRowIdx == _T_11 | commandsDone; // @[TensorLoadNarrowVME.scala 606:16 613:74 614:20]
  wire  _GEN_4 = _T_14 ? _GEN_2 : commandsDone; // @[TensorLoadNarrowVME.scala 606:16 610:31]
  wire  _GEN_6 = io_start | stride ? 1'h0 : _GEN_4; // @[TensorLoadNarrowVME.scala 607:29 609:18]
  wire  _T_20 = ~reset; // @[TensorLoadNarrowVME.scala 627:9]
  wire [15:0] _GEN_35 = {{12'd0}, dec_xpad_0}; // @[TensorLoadNarrowVME.scala 643:30]
  wire [15:0] _totalWidth_T_1 = dec_xsize + _GEN_35; // @[TensorLoadNarrowVME.scala 643:30]
  wire [15:0] _GEN_36 = {{12'd0}, dec_xpad_1}; // @[TensorLoadNarrowVME.scala 643:43]
  wire [15:0] totalWidth = _totalWidth_T_1 + _GEN_36; // @[TensorLoadNarrowVME.scala 643:43]
  reg [19:0] currentRowIdx; // @[TensorLoadNarrowVME.scala 647:26]
  wire [19:0] _GEN_37 = {{16'd0}, dec_ypad_0}; // @[TensorLoadNarrowVME.scala 649:39]
  wire [15:0] _GEN_38 = {{12'd0}, dec_ypad_0}; // @[TensorLoadNarrowVME.scala 650:32]
  wire [15:0] _rdCmdStartIdxValid_T_2 = dec_ysize + _GEN_38; // @[TensorLoadNarrowVME.scala 650:32]
  wire [19:0] _GEN_39 = {{4'd0}, _rdCmdStartIdxValid_T_2}; // @[TensorLoadNarrowVME.scala 650:19]
  wire  _rdCmdStartIdxValid_T_3 = currentRowIdx < _GEN_39; // @[TensorLoadNarrowVME.scala 650:19]
  wire  _rdCmdStartIdxValid_T_4 = currentRowIdx >= _GEN_37 & _rdCmdStartIdxValid_T_3; // @[TensorLoadNarrowVME.scala 649:53]
  wire  _rdCmdStartIdxValid_T_5 = _rdCmdStartIdxValid_T_4 & io_isBusy; // @[TensorLoadNarrowVME.scala 650:46]
  wire  _rdCmdStartIdxValid_T_6 = ~commandsDone; // @[TensorLoadNarrowVME.scala 652:5]
  wire  rdCmdStartIdxValid = _rdCmdStartIdxValid_T_5 & _rdCmdStartIdxValid_T_6; // @[TensorLoadNarrowVME.scala 651:15]
  wire [15:0] _rdCmdStartIdx_T_1 = dec_sram_offset + _GEN_35; // @[TensorLoadNarrowVME.scala 655:38]
  wire [15:0] _GEN_42 = {{9'd0}, rdCmdStartIdx}; // @[TensorLoadNarrowVME.scala 657:36]
  wire [15:0] _rdCmdStartIdx_T_3 = _GEN_42 + totalWidth; // @[TensorLoadNarrowVME.scala 657:36]
  wire [19:0] _currentRowIdx_T_1 = currentRowIdx + 20'h1; // @[TensorLoadNarrowVME.scala 658:36]
  wire [15:0] _GEN_11 = io_isBusy & (currentRowIdx < _GEN_37 | stride) ? _rdCmdStartIdx_T_3 : {{9'd0}, rdCmdStartIdx}; // @[TensorLoadNarrowVME.scala 656:68 657:19 586:26]
  wire [15:0] _GEN_14 = io_start ? _rdCmdStartIdx_T_1 : _GEN_11; // @[TensorLoadNarrowVME.scala 653:19 655:19]
  wire  startIssueCmdRead = blocksReadNb == 17'h0 & rdCmdStartIdxValid; // @[TensorLoadNarrowVME.scala 661:29]
  wire [19:0] _memRow_T = {dec_xstride, 4'h0}; // @[TensorLoadNarrowVME.scala 672:56]
  wire [31:0] _GEN_43 = {{12'd0}, _memRow_T}; // @[TensorLoadNarrowVME.scala 672:41]
  wire [31:0] memRow = rdCmdExtAddrRowBegin + _GEN_43; // @[TensorLoadNarrowVME.scala 672:41]
  wire [7:0] _rdCmdExtAddr_T = {readLen, 3'h0}; // @[TensorLoadNarrowVME.scala 679:47]
  wire [31:0] _GEN_44 = {{24'd0}, _rdCmdExtAddr_T}; // @[TensorLoadNarrowVME.scala 679:36]
  wire [31:0] _rdCmdExtAddr_T_2 = rdCmdExtAddr + _GEN_44; // @[TensorLoadNarrowVME.scala 679:36]
  wire [31:0] _GEN_16 = stride ? memRow : _rdCmdExtAddr_T_2; // @[TensorLoadNarrowVME.scala 671:18 673:20 679:20]
  wire [31:0] _GEN_17 = stride ? memRow : rdCmdExtAddrRowBegin; // @[TensorLoadNarrowVME.scala 671:18 664:24 674:28]
  wire [31:0] _GEN_19 = _T_14 ? _GEN_16 : rdCmdExtAddr; // @[TensorLoadNarrowVME.scala 670:31 682:18]
  wire [31:0] _GEN_20 = _T_14 ? _GEN_17 : rdCmdExtAddrRowBegin; // @[TensorLoadNarrowVME.scala 664:24 670:31]
  wire  _GEN_21 = _T_14 ? stride : newReadRow; // @[TensorLoadNarrowVME.scala 670:31 683:16]
  wire [35:0] _GEN_22 = io_start ? xfer_init_addr : {{4'd0}, _GEN_19}; // @[TensorLoadNarrowVME.scala 666:19 667:18]
  wire [35:0] _GEN_23 = io_start ? xfer_init_addr : {{4'd0}, _GEN_20}; // @[TensorLoadNarrowVME.scala 666:19 668:26]
  reg [7:0] rdCmdDestBlockIdxNext; // @[TensorLoadNarrowVME.scala 700:34]
  wire [7:0] _rdCmdDestBlockIdx_T = {rdCmdStartIdx, 1'h0}; // @[TensorLoadNarrowVME.scala 710:42]
  wire [7:0] _GEN_26 = startIssueCmdRead ? _rdCmdDestBlockIdx_T : rdCmdDestBlockIdxNext; // @[TensorLoadNarrowVME.scala 702:21 709:29 710:25]
  wire [7:0] rdCmdDestBlockIdx = rdCmdStartIdxValid ? _GEN_26 : rdCmdDestBlockIdxNext; // @[TensorLoadNarrowVME.scala 702:21 707:28]
  wire [7:0] _GEN_45 = {{3'd0}, readLen}; // @[TensorLoadNarrowVME.scala 711:49]
  wire [7:0] _rdCmdDestBlockIdxNext_T_1 = rdCmdDestBlockIdx + _GEN_45; // @[TensorLoadNarrowVME.scala 711:49]
  wire [7:0] _rdCmdDestBlockIdxNext_T_3 = rdCmdDestBlockIdxNext + _GEN_45; // @[TensorLoadNarrowVME.scala 714:53]
  wire [4:0] _io_vmeCmd_bits_len_T_1 = readLen - 5'h1; // @[TensorLoadNarrowVME.scala 732:33]
  assign io_vmeCmd_valid = _rdCmdStartIdxValid_T_5 & _rdCmdStartIdxValid_T_6; // @[TensorLoadNarrowVME.scala 651:15]
  assign io_vmeCmd_bits_addr = rdCmdExtAddr; // @[TensorLoadNarrowVME.scala 731:23]
  assign io_vmeCmd_bits_len = _io_vmeCmd_bits_len_T_1[3:0]; // @[TensorLoadNarrowVME.scala 732:22]
  assign io_vmeCmd_bits_tag = {{13'd0}, rdCmdDestBlockIdx}; // @[TensorLoadNarrowVME.scala 737:22]
  assign io_readLen = _GEN_10[4:0]; // @[TensorLoadNarrowVME.scala 587:21]
  assign io_done = commandsDone; // @[TensorLoadNarrowVME.scala 739:11]
  always @(posedge clock) begin
    rdCmdExtAddr <= _GEN_22[31:0];
    rdCmdStartIdx <= _GEN_14[6:0];
    commandsDone <= reset | _GEN_6; // @[TensorLoadNarrowVME.scala 588:{29,29}]
    if (io_start | stride) begin // @[TensorLoadNarrowVME.scala 607:29]
      blocksReadNb <= 17'h0; // @[TensorLoadNarrowVME.scala 608:18]
    end else if (_T_14) begin // @[TensorLoadNarrowVME.scala 610:31]
      blocksReadNb <= nextBlRNb; // @[TensorLoadNarrowVME.scala 612:18]
    end
    rdCmdExtAddrRowBegin <= _GEN_23[31:0];
    newReadRow <= io_start | _GEN_21; // @[TensorLoadNarrowVME.scala 666:19 669:16]
    if (io_start) begin // @[TensorLoadNarrowVME.scala 597:19]
      srcRowIdx <= 16'h0; // @[TensorLoadNarrowVME.scala 598:15]
    end else if (stride) begin // @[TensorLoadNarrowVME.scala 599:23]
      srcRowIdx <= _srcRowIdx_T_1; // @[TensorLoadNarrowVME.scala 600:15]
    end
    if (io_start) begin // @[TensorLoadNarrowVME.scala 653:19]
      currentRowIdx <= 20'h0; // @[TensorLoadNarrowVME.scala 654:19]
    end else if (io_isBusy & (currentRowIdx < _GEN_37 | stride)) begin // @[TensorLoadNarrowVME.scala 656:68]
      currentRowIdx <= _currentRowIdx_T_1; // @[TensorLoadNarrowVME.scala 658:19]
    end
    if (rdCmdStartIdxValid) begin // @[TensorLoadNarrowVME.scala 707:28]
      if (startIssueCmdRead) begin // @[TensorLoadNarrowVME.scala 709:29]
        rdCmdDestBlockIdxNext <= _rdCmdDestBlockIdxNext_T_1; // @[TensorLoadNarrowVME.scala 711:28]
      end else if (_T_14) begin // @[TensorLoadNarrowVME.scala 712:33]
        rdCmdDestBlockIdxNext <= _rdCmdDestBlockIdxNext_T_3; // @[TensorLoadNarrowVME.scala 714:28]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~io_isBusy | blocksReadSize >= blocksReadNb)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorLoadNarrowVME.scala:627 assert(!io.isBusy || blocksReadSize >= blocksReadNb)// define how many block to read at this cycle\n"
            ); // @[TensorLoadNarrowVME.scala 627:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_20 & ~(~io_vmeCmd_valid | _rdCmdExtAddr_T <= _firstMaxTransfer_T_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed: -F- inp DRAM page alignment failure. DRAM address + len overlaps mp.lenBits*memBlockSize alignment %x %x\n    at TensorLoadNarrowVME.scala:733 assert(!io.vmeCmd.valid || ((readLen << log2Ceil(mp.dataBits/8)) <= (maxTrBytes - rdCmdExtAddr %% maxTrBytes)),\n"
            ,rdCmdExtAddr,readLen); // @[TensorLoadNarrowVME.scala 733:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rdCmdExtAddr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  rdCmdStartIdx = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  commandsDone = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  blocksReadNb = _RAND_3[16:0];
  _RAND_4 = {1{`RANDOM}};
  rdCmdExtAddrRowBegin = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  newReadRow = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  srcRowIdx = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  currentRowIdx = _RAND_7[19:0];
  _RAND_8 = {1{`RANDOM}};
  rdCmdDestBlockIdxNext = _RAND_8[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~io_isBusy | blocksReadSize >= blocksReadNb); // @[TensorLoadNarrowVME.scala 627:9]
    end
    //
    if (_T_20) begin
      assert(~io_vmeCmd_valid | _rdCmdExtAddr_T <= _firstMaxTransfer_T_2); // @[TensorLoadNarrowVME.scala 733:9]
    end
  end
endmodule
module ReadVMEData(
  input         clock,
  input         reset,
  input         io_start,
  output        io_vmeData_ready,
  input         io_vmeData_valid,
  input  [20:0] io_vmeData_bits_tag,
  output [6:0]  io_idx,
  output        io_col
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [20:0] vmeTagDecodeLast; // @[TensorLoadNarrowVME.scala 502:29]
  wire [19:0] rdDataIdx = io_vmeData_bits_tag[20:1]; // @[TensorLoadNarrowVME.scala 503:31]
  wire  rdDataCol = io_vmeData_bits_tag[0]; // @[TensorLoadNarrowVME.scala 504:65]
  reg  rdDataDestColNext; // @[TensorLoadNarrowVME.scala 505:30]
  reg [15:0] rdDataDestIdxNext; // @[TensorLoadNarrowVME.scala 506:30]
  reg  vmeTagDecodeLastValidNext; // @[TensorLoadNarrowVME.scala 509:42]
  wire  _T = io_vmeData_ready & io_vmeData_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_0 = _T | vmeTagDecodeLastValidNext; // @[TensorLoadNarrowVME.scala 514:31 515:27 517:27]
  wire  _T_3 = io_vmeData_bits_tag != vmeTagDecodeLast; // @[TensorLoadNarrowVME.scala 525:29]
  wire  _T_4 = vmeTagDecodeLastValidNext & _T_3; // @[TensorLoadNarrowVME.scala 524:34]
  wire  _T_5 = ~vmeTagDecodeLastValidNext | _T_4; // @[TensorLoadNarrowVME.scala 523:34]
  wire  rdDataDestCol = _T_5 ? rdDataCol : rdDataDestColNext; // @[TensorLoadNarrowVME.scala 525:59 528:21 533:21]
  wire [15:0] _rdDataDestIdxNext_T_1 = rdDataDestIdxNext + 16'h1; // @[TensorLoadNarrowVME.scala 537:48]
  wire [15:0] _GEN_2 = rdDataDestCol ? _rdDataDestIdxNext_T_1 : rdDataDestIdxNext; // @[TensorLoadNarrowVME.scala 536:54 537:27 506:30]
  wire [19:0] _GEN_5 = _T_5 ? rdDataIdx : {{4'd0}, rdDataDestIdxNext}; // @[TensorLoadNarrowVME.scala 525:59 529:21 535:21]
  wire [19:0] _GEN_7 = _T_5 ? rdDataIdx : {{4'd0}, _GEN_2}; // @[TensorLoadNarrowVME.scala 525:59 531:25]
  wire [19:0] _GEN_12 = _T ? _GEN_7 : {{4'd0}, rdDataDestIdxNext}; // @[TensorLoadNarrowVME.scala 521:25 506:30]
  wire [15:0] rdDataDestIdx = _GEN_5[15:0]; // @[TensorLoadNarrowVME.scala 497:27]
  assign io_vmeData_ready = 1'h1; // @[TensorLoadNarrowVME.scala 498:20]
  assign io_idx = rdDataDestIdx[6:0]; // @[TensorLoadNarrowVME.scala 542:10]
  assign io_col = _T_5 ? rdDataCol : rdDataDestColNext; // @[TensorLoadNarrowVME.scala 525:59 528:21 533:21]
  always @(posedge clock) begin
    if (_T) begin // @[TensorLoadNarrowVME.scala 521:25]
      if (_T_5) begin // @[TensorLoadNarrowVME.scala 525:59]
        vmeTagDecodeLast <= io_vmeData_bits_tag; // @[TensorLoadNarrowVME.scala 527:24]
      end
    end
    if (_T) begin // @[TensorLoadNarrowVME.scala 521:25]
      if (_T_5) begin // @[TensorLoadNarrowVME.scala 525:59]
        rdDataDestColNext <= rdDataCol + 1'h1; // @[TensorLoadNarrowVME.scala 530:25]
      end else begin
        rdDataDestColNext <= rdDataDestColNext + 1'h1; // @[TensorLoadNarrowVME.scala 534:25]
      end
    end
    rdDataDestIdxNext <= _GEN_12[15:0];
    if (reset) begin // @[TensorLoadNarrowVME.scala 509:42]
      vmeTagDecodeLastValidNext <= 1'h0; // @[TensorLoadNarrowVME.scala 509:42]
    end else if (io_start) begin // @[TensorLoadNarrowVME.scala 512:18]
      vmeTagDecodeLastValidNext <= 1'h0; // @[TensorLoadNarrowVME.scala 513:27]
    end else begin
      vmeTagDecodeLastValidNext <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  vmeTagDecodeLast = _RAND_0[20:0];
  _RAND_1 = {1{`RANDOM}};
  rdDataDestColNext = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  rdDataDestIdxNext = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  vmeTagDecodeLastValidNext = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ZeroPadding(
  input          clock,
  input          reset,
  input          io_canWriteMem,
  input  [127:0] io_inst,
  output         io_tensorIdx_valid,
  output [6:0]   io_tensorIdx_bits,
  input          io_start,
  output         io_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] dec_sram_offset = io_inst[25:10]; // @[TensorLoadNarrowVME.scala 329:29]
  wire [15:0] dec_ysize = io_inst[79:64]; // @[TensorLoadNarrowVME.scala 329:29]
  wire [15:0] dec_xsize = io_inst[95:80]; // @[TensorLoadNarrowVME.scala 329:29]
  wire [3:0] dec_ypad_0 = io_inst[115:112]; // @[TensorLoadNarrowVME.scala 329:29]
  wire [3:0] dec_ypad_1 = io_inst[119:116]; // @[TensorLoadNarrowVME.scala 329:29]
  wire [3:0] dec_xpad_0 = io_inst[123:120]; // @[TensorLoadNarrowVME.scala 329:29]
  wire [3:0] dec_xpad_1 = io_inst[127:124]; // @[TensorLoadNarrowVME.scala 329:29]
  reg [2:0] zpState; // @[TensorLoadNarrowVME.scala 335:24]
  reg [23:0] zpColIdx; // @[TensorLoadNarrowVME.scala 337:21]
  reg [23:0] zpRowIdx; // @[TensorLoadNarrowVME.scala 340:21]
  reg [15:0] zpDestRowOffset; // @[TensorLoadNarrowVME.scala 342:28]
  wire [15:0] _GEN_35 = {{12'd0}, dec_ypad_0}; // @[TensorLoadNarrowVME.scala 349:47]
  wire [15:0] _zpLastDataRow_T_1 = _GEN_35 + dec_ysize; // @[TensorLoadNarrowVME.scala 349:47]
  wire [15:0] _zpLastDataRow_T_3 = _zpLastDataRow_T_1 - 16'h1; // @[TensorLoadNarrowVME.scala 349:59]
  wire [23:0] _GEN_36 = {{8'd0}, _zpLastDataRow_T_3}; // @[TensorLoadNarrowVME.scala 349:32]
  wire  zpLastDataRow = zpRowIdx == _GEN_36; // @[TensorLoadNarrowVME.scala 349:32]
  wire [15:0] _GEN_37 = {{12'd0}, dec_xpad_0}; // @[TensorLoadNarrowVME.scala 350:33]
  wire [15:0] _zpTopLastIdx_T_1 = _GEN_37 + dec_xsize; // @[TensorLoadNarrowVME.scala 350:33]
  wire [15:0] _GEN_38 = {{12'd0}, dec_xpad_1}; // @[TensorLoadNarrowVME.scala 350:45]
  wire [15:0] _zpTopLastIdx_T_3 = _zpTopLastIdx_T_1 + _GEN_38; // @[TensorLoadNarrowVME.scala 350:45]
  wire [15:0] zpTopLastIdx = _zpTopLastIdx_T_3 - 16'h1; // @[TensorLoadNarrowVME.scala 350:58]
  wire  _zpWideLineEnd_T = zpState == 3'h4; // @[TensorLoadNarrowVME.scala 351:32]
  wire  _zpWideLineEnd_T_1 = zpState == 3'h3; // @[TensorLoadNarrowVME.scala 351:59]
  wire [23:0] _GEN_39 = {{8'd0}, zpTopLastIdx}; // @[TensorLoadNarrowVME.scala 351:89]
  wire  _zpWideLineEnd_T_3 = zpColIdx == _GEN_39; // @[TensorLoadNarrowVME.scala 351:89]
  wire  zpWideLineEnd = (zpState == 3'h4 | zpState == 3'h3) & zpColIdx == _GEN_39; // @[TensorLoadNarrowVME.scala 351:77]
  wire [3:0] _zpNarwLineEnd_T_2 = dec_xpad_0 - 4'h1; // @[TensorLoadNarrowVME.scala 352:74]
  wire [23:0] _GEN_40 = {{20'd0}, _zpNarwLineEnd_T_2}; // @[TensorLoadNarrowVME.scala 352:59]
  wire  _zpNarwLineEnd_T_3 = zpColIdx == _GEN_40; // @[TensorLoadNarrowVME.scala 352:59]
  wire  zpNarwLineEnd = zpState == 3'h2 & zpColIdx == _GEN_40; // @[TensorLoadNarrowVME.scala 352:47]
  wire  zpFillLineEnd = zpWideLineEnd | zpNarwLineEnd; // @[TensorLoadNarrowVME.scala 353:37]
  wire  _T_1 = dec_xpad_1 != 4'h0; // @[TensorLoadNarrowVME.scala 360:43]
  wire  _T_2 = dec_xpad_0 == 4'h0 & dec_xpad_1 != 4'h0; // @[TensorLoadNarrowVME.scala 360:29]
  wire [15:0] _GEN_0 = dec_xpad_0 == 4'h0 & dec_xpad_1 != 4'h0 & dec_ypad_0 == 4'h0 ? _zpTopLastIdx_T_1 : 16'h0; // @[TensorLoadNarrowVME.scala 359:14 360:74 361:16]
  wire  _T_6 = dec_xpad_0 != 4'h0; // @[TensorLoadNarrowVME.scala 365:27]
  wire  _T_15 = dec_ypad_1 != 4'h0; // @[TensorLoadNarrowVME.scala 371:27]
  wire [2:0] _GEN_1 = dec_ypad_1 != 4'h0 ? 3'h5 : 3'h0; // @[TensorLoadNarrowVME.scala 371:36 372:15 374:15]
  wire [2:0] _GEN_2 = _T_6 & _T_1 ? 3'h4 : _GEN_1; // @[TensorLoadNarrowVME.scala 369:58 370:15]
  wire [2:0] _GEN_3 = _T_2 ? 3'h3 : _GEN_2; // @[TensorLoadNarrowVME.scala 367:58 368:15]
  wire [2:0] _GEN_4 = dec_xpad_0 != 4'h0 & dec_xpad_1 == 4'h0 ? 3'h2 : _GEN_3; // @[TensorLoadNarrowVME.scala 365:58 366:15]
  wire  _T_16 = zpState == 3'h1; // @[TensorLoadNarrowVME.scala 378:14]
  wire  _T_17 = io_canWriteMem & _T_16; // @[TensorLoadNarrowVME.scala 377:20]
  wire [3:0] _T_19 = dec_ypad_0 - 4'h1; // @[TensorLoadNarrowVME.scala 379:29]
  wire [23:0] _GEN_42 = {{20'd0}, _T_19}; // @[TensorLoadNarrowVME.scala 379:14]
  wire  _T_20 = zpRowIdx == _GEN_42; // @[TensorLoadNarrowVME.scala 379:14]
  wire  _T_21 = _T_17 & _T_20; // @[TensorLoadNarrowVME.scala 378:25]
  wire  _T_23 = _T_21 & _zpWideLineEnd_T_3; // @[TensorLoadNarrowVME.scala 379:35]
  wire [15:0] _GEN_6 = _T_2 ? _zpTopLastIdx_T_1 : 16'h0; // @[TensorLoadNarrowVME.scala 383:14 384:52 385:16]
  wire  _T_38 = zpState == 3'h5; // @[TensorLoadNarrowVME.scala 401:15]
  wire  _T_39 = zpFillLineEnd & io_canWriteMem | _T_38; // @[TensorLoadNarrowVME.scala 400:40]
  wire  _T_40 = zpLastDataRow & _T_39; // @[TensorLoadNarrowVME.scala 399:19]
  wire [23:0] _GEN_11 = _T_15 ? 24'h0 : zpColIdx; // @[TensorLoadNarrowVME.scala 344:12 405:30 406:16]
  wire [2:0] _GEN_12 = _T_15 ? 3'h6 : 3'h0; // @[TensorLoadNarrowVME.scala 405:30 407:15 409:15]
  wire  _T_42 = zpState == 3'h6; // @[TensorLoadNarrowVME.scala 413:14]
  wire  _T_43 = io_canWriteMem & _T_42; // @[TensorLoadNarrowVME.scala 412:20]
  wire [15:0] _GEN_46 = {{12'd0}, dec_ypad_1}; // @[TensorLoadNarrowVME.scala 414:41]
  wire [15:0] _T_47 = _zpLastDataRow_T_1 + _GEN_46; // @[TensorLoadNarrowVME.scala 414:41]
  wire [15:0] _T_49 = _T_47 - 16'h1; // @[TensorLoadNarrowVME.scala 414:54]
  wire [23:0] _GEN_47 = {{8'd0}, _T_49}; // @[TensorLoadNarrowVME.scala 414:14]
  wire  _T_50 = zpRowIdx == _GEN_47; // @[TensorLoadNarrowVME.scala 414:14]
  wire  _T_51 = _T_43 & _T_50; // @[TensorLoadNarrowVME.scala 413:25]
  wire  _T_53 = _T_51 & _zpWideLineEnd_T_3; // @[TensorLoadNarrowVME.scala 414:60]
  wire [23:0] _GEN_14 = _T_53 ? 24'h0 : zpColIdx; // @[TensorLoadNarrowVME.scala 344:12 415:32 418:14]
  wire [2:0] _GEN_15 = _T_53 ? 3'h0 : zpState; // @[TensorLoadNarrowVME.scala 415:32 419:13 421:13]
  wire  _GEN_16 = _T_40 | _T_53; // @[TensorLoadNarrowVME.scala 401:63 403:20]
  wire [23:0] _GEN_17 = _T_40 ? _GEN_11 : _GEN_14; // @[TensorLoadNarrowVME.scala 401:63]
  wire  _GEN_19 = _T_23 | _GEN_16; // @[TensorLoadNarrowVME.scala 380:32 381:20]
  wire [23:0] _GEN_20 = _T_23 ? {{8'd0}, _GEN_6} : _GEN_17; // @[TensorLoadNarrowVME.scala 380:32]
  wire [23:0] _GEN_24 = io_start ? {{8'd0}, _GEN_0} : _GEN_20; // @[TensorLoadNarrowVME.scala 355:18]
  wire  zpNewFillBlock = io_start ? 1'h0 : _GEN_19; // @[TensorLoadNarrowVME.scala 346:18 355:18]
  wire  isZeroPadWrite = zpState != 3'h0 & zpState != 3'h5 & io_canWriteMem; // @[TensorLoadNarrowVME.scala 424:68]
  wire [23:0] _GEN_49 = {{8'd0}, zpDestRowOffset}; // @[TensorLoadNarrowVME.scala 425:32]
  wire [23:0] _zpDestIdx_T_1 = _GEN_49 + zpColIdx; // @[TensorLoadNarrowVME.scala 425:32]
  wire  _T_62 = (_T_16 | _zpWideLineEnd_T | _zpWideLineEnd_T_1 | _T_42) & _zpWideLineEnd_T_3; // @[TensorLoadNarrowVME.scala 432:106]
  wire  _T_68 = _T_62 | zpNarwLineEnd; // @[TensorLoadNarrowVME.scala 433:34]
  wire  incrementRow = _T_68 & io_canWriteMem | _T_38; // @[TensorLoadNarrowVME.scala 434:84]
  wire [15:0] _zpDestRowOffset_T_1 = zpDestRowOffset + zpTopLastIdx; // @[TensorLoadNarrowVME.scala 437:40]
  wire [15:0] _zpDestRowOffset_T_3 = _zpDestRowOffset_T_1 + 16'h1; // @[TensorLoadNarrowVME.scala 437:55]
  wire [23:0] _zpRowIdx_T_1 = zpRowIdx + 24'h1; // @[TensorLoadNarrowVME.scala 438:26]
  wire  _T_72 = ~zpNewFillBlock; // @[TensorLoadNarrowVME.scala 440:10]
  wire [15:0] _GEN_27 = _zpWideLineEnd_T_1 ? _zpTopLastIdx_T_1 : 16'h0; // @[TensorLoadNarrowVME.scala 441:38 442:18 444:18]
  wire [23:0] _GEN_54 = {{8'd0}, dec_xsize}; // @[TensorLoadNarrowVME.scala 452:28]
  wire [23:0] _zpColIdx_T_7 = zpColIdx + _GEN_54; // @[TensorLoadNarrowVME.scala 452:28]
  wire [23:0] _zpColIdx_T_9 = _zpColIdx_T_7 + 24'h1; // @[TensorLoadNarrowVME.scala 452:40]
  wire [23:0] _zpColIdx_T_11 = zpColIdx + 24'h1; // @[TensorLoadNarrowVME.scala 455:28]
  wire [15:0] zpDestIdx = _zpDestIdx_T_1[15:0]; // @[TensorLoadNarrowVME.scala 332:23 425:13]
  assign io_tensorIdx_valid = zpState != 3'h0 & zpState != 3'h5 & io_canWriteMem; // @[TensorLoadNarrowVME.scala 424:68]
  assign io_tensorIdx_bits = zpDestIdx[6:0]; // @[TensorLoadNarrowVME.scala 460:21]
  assign io_done = zpState == 3'h0; // @[TensorLoadNarrowVME.scala 458:22]
  always @(posedge clock) begin
    if (reset) begin // @[TensorLoadNarrowVME.scala 335:24]
      zpState <= 3'h0; // @[TensorLoadNarrowVME.scala 335:24]
    end else if (io_start) begin // @[TensorLoadNarrowVME.scala 355:18]
      if (dec_ypad_0 != 4'h0) begin // @[TensorLoadNarrowVME.scala 363:30]
        zpState <= 3'h1; // @[TensorLoadNarrowVME.scala 364:15]
      end else begin
        zpState <= _GEN_4;
      end
    end else if (_T_23) begin // @[TensorLoadNarrowVME.scala 380:32]
      zpState <= _GEN_4;
    end else if (_T_40) begin // @[TensorLoadNarrowVME.scala 401:63]
      zpState <= _GEN_12;
    end else begin
      zpState <= _GEN_15;
    end
    if (isZeroPadWrite & _T_72 & ~incrementRow) begin // @[TensorLoadNarrowVME.scala 450:60]
      if (_zpWideLineEnd_T & _zpNarwLineEnd_T_3) begin // @[TensorLoadNarrowVME.scala 451:68]
        zpColIdx <= _zpColIdx_T_9; // @[TensorLoadNarrowVME.scala 452:16]
      end else begin
        zpColIdx <= _zpColIdx_T_11; // @[TensorLoadNarrowVME.scala 455:16]
      end
    end else if (incrementRow) begin // @[TensorLoadNarrowVME.scala 435:30]
      if (~zpNewFillBlock) begin // @[TensorLoadNarrowVME.scala 440:27]
        zpColIdx <= {{8'd0}, _GEN_27};
      end else begin
        zpColIdx <= _GEN_24;
      end
    end else begin
      zpColIdx <= _GEN_24;
    end
    if (incrementRow) begin // @[TensorLoadNarrowVME.scala 435:30]
      zpRowIdx <= _zpRowIdx_T_1; // @[TensorLoadNarrowVME.scala 438:14]
    end else if (io_start) begin // @[TensorLoadNarrowVME.scala 355:18]
      zpRowIdx <= 24'h0; // @[TensorLoadNarrowVME.scala 356:14]
    end
    if (incrementRow) begin // @[TensorLoadNarrowVME.scala 435:30]
      zpDestRowOffset <= _zpDestRowOffset_T_3; // @[TensorLoadNarrowVME.scala 437:21]
    end else if (io_start) begin // @[TensorLoadNarrowVME.scala 355:18]
      zpDestRowOffset <= dec_sram_offset; // @[TensorLoadNarrowVME.scala 357:21]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  zpState = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  zpColIdx = _RAND_1[23:0];
  _RAND_2 = {1{`RANDOM}};
  zpRowIdx = _RAND_2[23:0];
  _RAND_3 = {1{`RANDOM}};
  zpDestRowOffset = _RAND_3[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TensorLoadNarrowVME(
  input          clock,
  input          reset,
  input          io_start,
  output         io_done,
  input  [127:0] io_inst,
  input  [31:0]  io_baddr,
  input          io_vme_rd_cmd_ready,
  output         io_vme_rd_cmd_valid,
  output [31:0]  io_vme_rd_cmd_bits_addr,
  output [3:0]   io_vme_rd_cmd_bits_len,
  output [20:0]  io_vme_rd_cmd_bits_tag,
  output         io_vme_rd_data_ready,
  input          io_vme_rd_data_valid,
  input  [63:0]  io_vme_rd_data_bits_data,
  input  [20:0]  io_vme_rd_data_bits_tag,
  input          io_tensor_rd_0_idx_valid,
  input  [6:0]   io_tensor_rd_0_idx_bits,
  output         io_tensor_rd_0_data_valid,
  output [7:0]   io_tensor_rd_0_data_bits_0_0,
  output [7:0]   io_tensor_rd_0_data_bits_0_1,
  output [7:0]   io_tensor_rd_0_data_bits_0_2,
  output [7:0]   io_tensor_rd_0_data_bits_0_3,
  output [7:0]   io_tensor_rd_0_data_bits_0_4,
  output [7:0]   io_tensor_rd_0_data_bits_0_5,
  output [7:0]   io_tensor_rd_0_data_bits_0_6,
  output [7:0]   io_tensor_rd_0_data_bits_0_7,
  output [7:0]   io_tensor_rd_0_data_bits_0_8,
  output [7:0]   io_tensor_rd_0_data_bits_0_9,
  output [7:0]   io_tensor_rd_0_data_bits_0_10,
  output [7:0]   io_tensor_rd_0_data_bits_0_11,
  output [7:0]   io_tensor_rd_0_data_bits_0_12,
  output [7:0]   io_tensor_rd_0_data_bits_0_13,
  output [7:0]   io_tensor_rd_0_data_bits_0_14,
  output [7:0]   io_tensor_rd_0_data_bits_0_15
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [127:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_REG_INIT
  wire  vmeCmd_clock; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_reset; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_start; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_isBusy; // @[TensorLoadNarrowVME.scala 75:23]
  wire [127:0] vmeCmd_io_inst; // @[TensorLoadNarrowVME.scala 75:23]
  wire [31:0] vmeCmd_io_baddr; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_vmeCmd_ready; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_vmeCmd_valid; // @[TensorLoadNarrowVME.scala 75:23]
  wire [31:0] vmeCmd_io_vmeCmd_bits_addr; // @[TensorLoadNarrowVME.scala 75:23]
  wire [3:0] vmeCmd_io_vmeCmd_bits_len; // @[TensorLoadNarrowVME.scala 75:23]
  wire [20:0] vmeCmd_io_vmeCmd_bits_tag; // @[TensorLoadNarrowVME.scala 75:23]
  wire [4:0] vmeCmd_io_readLen; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_done; // @[TensorLoadNarrowVME.scala 75:23]
  wire  readData_clock; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_reset; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_io_start; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_io_vmeData_ready; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_io_vmeData_valid; // @[TensorLoadNarrowVME.scala 105:24]
  wire [20:0] readData_io_vmeData_bits_tag; // @[TensorLoadNarrowVME.scala 105:24]
  wire [6:0] readData_io_idx; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_io_col; // @[TensorLoadNarrowVME.scala 105:24]
  wire  fillPadding_clock; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_reset; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_io_canWriteMem; // @[TensorLoadNarrowVME.scala 119:27]
  wire [127:0] fillPadding_io_inst; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_io_tensorIdx_valid; // @[TensorLoadNarrowVME.scala 119:27]
  wire [6:0] fillPadding_io_tensorIdx_bits; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_io_start; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_io_done; // @[TensorLoadNarrowVME.scala 119:27]
  reg [63:0] tensorFile_0 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_0_MPORT_2_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_0_MPORT_2_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_0_MPORT_2_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_0_MPORT_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_0_MPORT_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_0_MPORT_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_0_MPORT_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_0_MPORT_2_en_pipe_0;
  reg [6:0] tensorFile_0_MPORT_2_addr_pipe_0;
  reg [63:0] tensorFile_1 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_1_MPORT_3_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_1_MPORT_3_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_1_MPORT_3_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_1_MPORT_1_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_1_MPORT_1_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_1_MPORT_1_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_1_MPORT_1_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_1_MPORT_3_en_pipe_0;
  reg [6:0] tensorFile_1_MPORT_3_addr_pipe_0;
  reg  state; // @[TensorLoadNarrowVME.scala 54:22]
  reg [7:0] blocksInFlight; // @[TensorLoadNarrowVME.scala 87:27]
  wire  loadDone = blocksInFlight == 8'h0 & vmeCmd_io_done & state; // @[TensorLoadNarrowVME.scala 292:57]
  wire  localDone = loadDone & fillPadding_io_done; // @[TensorLoadNarrowVME.scala 293:25]
  wire  _GEN_0 = localDone ? 1'h0 : state; // @[TensorLoadNarrowVME.scala 61:25 62:11 54:22]
  wire  _GEN_1 = io_start | _GEN_0; // @[TensorLoadNarrowVME.scala 59:18 60:11]
  reg [63:0] vmeDataBitsPipe_data; // @[TensorLoadNarrowVME.scala 67:32]
  reg [20:0] vmeDataBitsPipe_tag; // @[TensorLoadNarrowVME.scala 67:32]
  reg  vmeDataValidPipe; // @[TensorLoadNarrowVME.scala 68:33]
  reg  vmeDataReadyPipe; // @[TensorLoadNarrowVME.scala 69:33]
  wire  vmeDataFirePipe = vmeDataValidPipe & vmeDataReadyPipe; // @[TensorLoadNarrowVME.scala 70:42]
  wire  _T = io_vme_rd_cmd_ready & io_vme_rd_cmd_valid; // @[Decoupled.scala 50:35]
  wire  _T_1 = state & _T; // @[TensorLoadNarrowVME.scala 90:21]
  wire  _T_3 = state & _T & ~vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 90:43]
  wire [7:0] _GEN_22 = {{3'd0}, vmeCmd_io_readLen}; // @[TensorLoadNarrowVME.scala 91:38]
  wire [7:0] _blocksInFlight_T_1 = blocksInFlight + _GEN_22; // @[TensorLoadNarrowVME.scala 91:38]
  wire  _T_6 = _T_1 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 92:43]
  wire [7:0] _blocksInFlight_T_5 = _blocksInFlight_T_1 - 8'h1; // @[TensorLoadNarrowVME.scala 93:48]
  wire  _T_10 = state & ~_T & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 94:44]
  wire  _T_13 = ~reset; // @[TensorLoadNarrowVME.scala 95:11]
  wire [7:0] _blocksInFlight_T_7 = blocksInFlight - 8'h1; // @[TensorLoadNarrowVME.scala 96:38]
  reg [127:0] fillPadding_io_inst_REG; // @[TensorLoadNarrowVME.scala 121:33]
  reg  fillPadding_io_start_REG; // @[TensorLoadNarrowVME.scala 122:34]
  wire [6:0] waddrTensInstrTmp = fillPadding_io_tensorIdx_valid ? fillPadding_io_tensorIdx_bits : readData_io_idx; // @[TensorLoadNarrowVME.scala 166:30]
  wire  _waddr_0_T = ~state; // @[TensorLoadNarrowVME.scala 186:27]
  wire  wenTensInstr_0 = fillPadding_io_tensorIdx_valid | ~readData_io_col & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_1 = fillPadding_io_tensorIdx_valid | readData_io_col & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire [63:0] wdataTensInstr_0 = fillPadding_io_tensorIdx_valid ? 64'h0 : vmeDataBitsPipe_data; // @[TensorLoadNarrowVME.scala 234:29]
  reg  rvalid; // @[Reg.scala 28:20]
  wire [63:0] _WIRE_2_1 = tensorFile_1_MPORT_3_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_2_0 = tensorFile_0_MPORT_2_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [127:0] _T_24 = {_WIRE_2_1,_WIRE_2_0}; // @[TensorLoadNarrowVME.scala 288:18]
  GenVMECmd vmeCmd ( // @[TensorLoadNarrowVME.scala 75:23]
    .clock(vmeCmd_clock),
    .reset(vmeCmd_reset),
    .io_start(vmeCmd_io_start),
    .io_isBusy(vmeCmd_io_isBusy),
    .io_inst(vmeCmd_io_inst),
    .io_baddr(vmeCmd_io_baddr),
    .io_vmeCmd_ready(vmeCmd_io_vmeCmd_ready),
    .io_vmeCmd_valid(vmeCmd_io_vmeCmd_valid),
    .io_vmeCmd_bits_addr(vmeCmd_io_vmeCmd_bits_addr),
    .io_vmeCmd_bits_len(vmeCmd_io_vmeCmd_bits_len),
    .io_vmeCmd_bits_tag(vmeCmd_io_vmeCmd_bits_tag),
    .io_readLen(vmeCmd_io_readLen),
    .io_done(vmeCmd_io_done)
  );
  ReadVMEData readData ( // @[TensorLoadNarrowVME.scala 105:24]
    .clock(readData_clock),
    .reset(readData_reset),
    .io_start(readData_io_start),
    .io_vmeData_ready(readData_io_vmeData_ready),
    .io_vmeData_valid(readData_io_vmeData_valid),
    .io_vmeData_bits_tag(readData_io_vmeData_bits_tag),
    .io_idx(readData_io_idx),
    .io_col(readData_io_col)
  );
  ZeroPadding fillPadding ( // @[TensorLoadNarrowVME.scala 119:27]
    .clock(fillPadding_clock),
    .reset(fillPadding_reset),
    .io_canWriteMem(fillPadding_io_canWriteMem),
    .io_inst(fillPadding_io_inst),
    .io_tensorIdx_valid(fillPadding_io_tensorIdx_valid),
    .io_tensorIdx_bits(fillPadding_io_tensorIdx_bits),
    .io_start(fillPadding_io_start),
    .io_done(fillPadding_io_done)
  );
  assign tensorFile_0_MPORT_2_en = tensorFile_0_MPORT_2_en_pipe_0;
  assign tensorFile_0_MPORT_2_addr = tensorFile_0_MPORT_2_addr_pipe_0;
  assign tensorFile_0_MPORT_2_data = tensorFile_0[tensorFile_0_MPORT_2_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_0_MPORT_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_0_MPORT_addr = _waddr_0_T ? 7'h0 : waddrTensInstrTmp;
  assign tensorFile_0_MPORT_mask = 1'h1;
  assign tensorFile_0_MPORT_en = _waddr_0_T ? 1'h0 : wenTensInstr_0;
  assign tensorFile_1_MPORT_3_en = tensorFile_1_MPORT_3_en_pipe_0;
  assign tensorFile_1_MPORT_3_addr = tensorFile_1_MPORT_3_addr_pipe_0;
  assign tensorFile_1_MPORT_3_data = tensorFile_1[tensorFile_1_MPORT_3_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_1_MPORT_1_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_1_MPORT_1_addr = _waddr_0_T ? 7'h0 : waddrTensInstrTmp;
  assign tensorFile_1_MPORT_1_mask = 1'h1;
  assign tensorFile_1_MPORT_1_en = _waddr_0_T ? 1'h0 : wenTensInstr_1;
  assign io_done = loadDone & fillPadding_io_done; // @[TensorLoadNarrowVME.scala 293:25]
  assign io_vme_rd_cmd_valid = vmeCmd_io_vmeCmd_valid; // @[TensorLoadNarrowVME.scala 80:20]
  assign io_vme_rd_cmd_bits_addr = vmeCmd_io_vmeCmd_bits_addr; // @[TensorLoadNarrowVME.scala 80:20]
  assign io_vme_rd_cmd_bits_len = vmeCmd_io_vmeCmd_bits_len; // @[TensorLoadNarrowVME.scala 80:20]
  assign io_vme_rd_cmd_bits_tag = vmeCmd_io_vmeCmd_bits_tag; // @[TensorLoadNarrowVME.scala 80:20]
  assign io_vme_rd_data_ready = 1'h1; // @[TensorLoadNarrowVME.scala 111:24]
  assign io_tensor_rd_0_data_valid = rvalid; // @[TensorLoadNarrowVME.scala 278:36]
  assign io_tensor_rd_0_data_bits_0_0 = _T_24[7:0]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_1 = _T_24[15:8]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_2 = _T_24[23:16]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_3 = _T_24[31:24]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_4 = _T_24[39:32]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_5 = _T_24[47:40]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_6 = _T_24[55:48]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_7 = _T_24[63:56]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_8 = _T_24[71:64]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_9 = _T_24[79:72]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_10 = _T_24[87:80]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_11 = _T_24[95:88]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_12 = _T_24[103:96]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_13 = _T_24[111:104]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_14 = _T_24[119:112]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_15 = _T_24[127:120]; // @[TensorLoadNarrowVME.scala 288:18]
  assign vmeCmd_clock = clock;
  assign vmeCmd_reset = reset;
  assign vmeCmd_io_start = io_start; // @[TensorLoadNarrowVME.scala 76:19]
  assign vmeCmd_io_isBusy = state; // @[TensorLoadNarrowVME.scala 56:22]
  assign vmeCmd_io_inst = io_inst; // @[TensorLoadNarrowVME.scala 78:18]
  assign vmeCmd_io_baddr = io_baddr; // @[TensorLoadNarrowVME.scala 79:19]
  assign vmeCmd_io_vmeCmd_ready = io_vme_rd_cmd_ready; // @[TensorLoadNarrowVME.scala 80:20]
  assign readData_clock = clock;
  assign readData_reset = reset;
  assign readData_io_start = io_start; // @[TensorLoadNarrowVME.scala 106:21]
  assign readData_io_vmeData_valid = vmeDataValidPipe; // @[TensorLoadNarrowVME.scala 107:29]
  assign readData_io_vmeData_bits_tag = vmeDataBitsPipe_tag; // @[TensorLoadNarrowVME.scala 108:28]
  assign fillPadding_clock = clock;
  assign fillPadding_reset = reset;
  assign fillPadding_io_canWriteMem = ~vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 120:33]
  assign fillPadding_io_inst = fillPadding_io_inst_REG; // @[TensorLoadNarrowVME.scala 121:23]
  assign fillPadding_io_start = fillPadding_io_start_REG; // @[TensorLoadNarrowVME.scala 122:24]
  always @(posedge clock) begin
    if (tensorFile_0_MPORT_en & tensorFile_0_MPORT_mask) begin
      tensorFile_0[tensorFile_0_MPORT_addr] <= tensorFile_0_MPORT_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_0_MPORT_2_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_0_MPORT_2_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_1_MPORT_1_en & tensorFile_1_MPORT_1_mask) begin
      tensorFile_1[tensorFile_1_MPORT_1_addr] <= tensorFile_1_MPORT_1_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_1_MPORT_3_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_1_MPORT_3_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (reset) begin // @[TensorLoadNarrowVME.scala 54:22]
      state <= 1'h0; // @[TensorLoadNarrowVME.scala 54:22]
    end else begin
      state <= _GEN_1;
    end
    if (io_start) begin // @[TensorLoadNarrowVME.scala 88:18]
      blocksInFlight <= 8'h0; // @[TensorLoadNarrowVME.scala 89:20]
    end else if (state & _T & ~vmeDataFirePipe) begin // @[TensorLoadNarrowVME.scala 90:64]
      blocksInFlight <= _blocksInFlight_T_1; // @[TensorLoadNarrowVME.scala 91:20]
    end else if (_T_1 & vmeDataFirePipe) begin // @[TensorLoadNarrowVME.scala 92:63]
      blocksInFlight <= _blocksInFlight_T_5; // @[TensorLoadNarrowVME.scala 93:20]
    end else if (state & ~_T & vmeDataFirePipe) begin // @[TensorLoadNarrowVME.scala 94:64]
      blocksInFlight <= _blocksInFlight_T_7; // @[TensorLoadNarrowVME.scala 96:20]
    end
    vmeDataBitsPipe_data <= io_vme_rd_data_bits_data; // @[TensorLoadNarrowVME.scala 67:32]
    vmeDataBitsPipe_tag <= io_vme_rd_data_bits_tag; // @[TensorLoadNarrowVME.scala 67:32]
    if (reset) begin // @[TensorLoadNarrowVME.scala 68:33]
      vmeDataValidPipe <= 1'h0; // @[TensorLoadNarrowVME.scala 68:33]
    end else begin
      vmeDataValidPipe <= io_vme_rd_data_valid; // @[TensorLoadNarrowVME.scala 68:33]
    end
    if (reset) begin // @[TensorLoadNarrowVME.scala 69:33]
      vmeDataReadyPipe <= 1'h0; // @[TensorLoadNarrowVME.scala 69:33]
    end else begin
      vmeDataReadyPipe <= io_vme_rd_data_ready; // @[TensorLoadNarrowVME.scala 69:33]
    end
    fillPadding_io_inst_REG <= io_inst; // @[TensorLoadNarrowVME.scala 121:33]
    if (reset) begin // @[TensorLoadNarrowVME.scala 122:34]
      fillPadding_io_start_REG <= 1'h0; // @[TensorLoadNarrowVME.scala 122:34]
    end else begin
      fillPadding_io_start_REG <= io_start; // @[TensorLoadNarrowVME.scala 122:34]
    end
    if (reset) begin // @[Reg.scala 28:20]
      rvalid <= 1'h0; // @[Reg.scala 28:20]
    end else begin
      rvalid <= io_tensor_rd_0_idx_valid;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~io_start & ~_T_3 & ~_T_6 & _T_10 & ~reset & ~(blocksInFlight > 8'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TensorLoadNarrowVME.scala:95 assert(blocksInFlight > 0.U)\n"); // @[TensorLoadNarrowVME.scala 95:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_0[initvar] = _RAND_0[63:0];
  _RAND_3 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_1[initvar] = _RAND_3[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tensorFile_0_MPORT_2_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  tensorFile_0_MPORT_2_addr_pipe_0 = _RAND_2[6:0];
  _RAND_4 = {1{`RANDOM}};
  tensorFile_1_MPORT_3_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  tensorFile_1_MPORT_3_addr_pipe_0 = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  blocksInFlight = _RAND_7[7:0];
  _RAND_8 = {2{`RANDOM}};
  vmeDataBitsPipe_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  vmeDataBitsPipe_tag = _RAND_9[20:0];
  _RAND_10 = {1{`RANDOM}};
  vmeDataValidPipe = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  vmeDataReadyPipe = _RAND_11[0:0];
  _RAND_12 = {4{`RANDOM}};
  fillPadding_io_inst_REG = _RAND_12[127:0];
  _RAND_13 = {1{`RANDOM}};
  fillPadding_io_start_REG = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  rvalid = _RAND_14[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~io_start & ~_T_3 & ~_T_6 & _T_10 & ~reset) begin
      assert(blocksInFlight > 8'h0); // @[TensorLoadNarrowVME.scala 95:11]
    end
    //
    if (_T_13) begin
      assert(1'h1); // @[TensorLoadNarrowVME.scala 109:9]
    end
  end
endmodule
module TensorLoadInp(
  input          clock,
  input          reset,
  input          io_start,
  output         io_done,
  input  [127:0] io_inst,
  input  [31:0]  io_baddr,
  input          io_vme_rd_cmd_ready,
  output         io_vme_rd_cmd_valid,
  output [31:0]  io_vme_rd_cmd_bits_addr,
  output [3:0]   io_vme_rd_cmd_bits_len,
  output [20:0]  io_vme_rd_cmd_bits_tag,
  input          io_vme_rd_data_valid,
  input  [63:0]  io_vme_rd_data_bits_data,
  input  [20:0]  io_vme_rd_data_bits_tag,
  input          io_tensor_rd_0_idx_valid,
  input  [6:0]   io_tensor_rd_0_idx_bits,
  output         io_tensor_rd_0_data_valid,
  output [7:0]   io_tensor_rd_0_data_bits_0_0,
  output [7:0]   io_tensor_rd_0_data_bits_0_1,
  output [7:0]   io_tensor_rd_0_data_bits_0_2,
  output [7:0]   io_tensor_rd_0_data_bits_0_3,
  output [7:0]   io_tensor_rd_0_data_bits_0_4,
  output [7:0]   io_tensor_rd_0_data_bits_0_5,
  output [7:0]   io_tensor_rd_0_data_bits_0_6,
  output [7:0]   io_tensor_rd_0_data_bits_0_7,
  output [7:0]   io_tensor_rd_0_data_bits_0_8,
  output [7:0]   io_tensor_rd_0_data_bits_0_9,
  output [7:0]   io_tensor_rd_0_data_bits_0_10,
  output [7:0]   io_tensor_rd_0_data_bits_0_11,
  output [7:0]   io_tensor_rd_0_data_bits_0_12,
  output [7:0]   io_tensor_rd_0_data_bits_0_13,
  output [7:0]   io_tensor_rd_0_data_bits_0_14,
  output [7:0]   io_tensor_rd_0_data_bits_0_15
);
  wire  tensorLoad_clock; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_reset; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_start; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_done; // @[TensorLoad.scala 71:28]
  wire [127:0] tensorLoad_io_inst; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_baddr; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_vme_rd_cmd_ready; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_vme_rd_cmd_valid; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_vme_rd_cmd_bits_addr; // @[TensorLoad.scala 71:28]
  wire [3:0] tensorLoad_io_vme_rd_cmd_bits_len; // @[TensorLoad.scala 71:28]
  wire [20:0] tensorLoad_io_vme_rd_cmd_bits_tag; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_vme_rd_data_ready; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_vme_rd_data_valid; // @[TensorLoad.scala 71:28]
  wire [63:0] tensorLoad_io_vme_rd_data_bits_data; // @[TensorLoad.scala 71:28]
  wire [20:0] tensorLoad_io_vme_rd_data_bits_tag; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_tensor_rd_0_idx_valid; // @[TensorLoad.scala 71:28]
  wire [6:0] tensorLoad_io_tensor_rd_0_idx_bits; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_tensor_rd_0_data_valid; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_15; // @[TensorLoad.scala 71:28]
  TensorLoadNarrowVME tensorLoad ( // @[TensorLoad.scala 71:28]
    .clock(tensorLoad_clock),
    .reset(tensorLoad_reset),
    .io_start(tensorLoad_io_start),
    .io_done(tensorLoad_io_done),
    .io_inst(tensorLoad_io_inst),
    .io_baddr(tensorLoad_io_baddr),
    .io_vme_rd_cmd_ready(tensorLoad_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(tensorLoad_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(tensorLoad_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(tensorLoad_io_vme_rd_cmd_bits_len),
    .io_vme_rd_cmd_bits_tag(tensorLoad_io_vme_rd_cmd_bits_tag),
    .io_vme_rd_data_ready(tensorLoad_io_vme_rd_data_ready),
    .io_vme_rd_data_valid(tensorLoad_io_vme_rd_data_valid),
    .io_vme_rd_data_bits_data(tensorLoad_io_vme_rd_data_bits_data),
    .io_vme_rd_data_bits_tag(tensorLoad_io_vme_rd_data_bits_tag),
    .io_tensor_rd_0_idx_valid(tensorLoad_io_tensor_rd_0_idx_valid),
    .io_tensor_rd_0_idx_bits(tensorLoad_io_tensor_rd_0_idx_bits),
    .io_tensor_rd_0_data_valid(tensorLoad_io_tensor_rd_0_data_valid),
    .io_tensor_rd_0_data_bits_0_0(tensorLoad_io_tensor_rd_0_data_bits_0_0),
    .io_tensor_rd_0_data_bits_0_1(tensorLoad_io_tensor_rd_0_data_bits_0_1),
    .io_tensor_rd_0_data_bits_0_2(tensorLoad_io_tensor_rd_0_data_bits_0_2),
    .io_tensor_rd_0_data_bits_0_3(tensorLoad_io_tensor_rd_0_data_bits_0_3),
    .io_tensor_rd_0_data_bits_0_4(tensorLoad_io_tensor_rd_0_data_bits_0_4),
    .io_tensor_rd_0_data_bits_0_5(tensorLoad_io_tensor_rd_0_data_bits_0_5),
    .io_tensor_rd_0_data_bits_0_6(tensorLoad_io_tensor_rd_0_data_bits_0_6),
    .io_tensor_rd_0_data_bits_0_7(tensorLoad_io_tensor_rd_0_data_bits_0_7),
    .io_tensor_rd_0_data_bits_0_8(tensorLoad_io_tensor_rd_0_data_bits_0_8),
    .io_tensor_rd_0_data_bits_0_9(tensorLoad_io_tensor_rd_0_data_bits_0_9),
    .io_tensor_rd_0_data_bits_0_10(tensorLoad_io_tensor_rd_0_data_bits_0_10),
    .io_tensor_rd_0_data_bits_0_11(tensorLoad_io_tensor_rd_0_data_bits_0_11),
    .io_tensor_rd_0_data_bits_0_12(tensorLoad_io_tensor_rd_0_data_bits_0_12),
    .io_tensor_rd_0_data_bits_0_13(tensorLoad_io_tensor_rd_0_data_bits_0_13),
    .io_tensor_rd_0_data_bits_0_14(tensorLoad_io_tensor_rd_0_data_bits_0_14),
    .io_tensor_rd_0_data_bits_0_15(tensorLoad_io_tensor_rd_0_data_bits_0_15)
  );
  assign io_done = tensorLoad_io_done; // @[TensorLoad.scala 72:8]
  assign io_vme_rd_cmd_valid = tensorLoad_io_vme_rd_cmd_valid; // @[TensorLoad.scala 72:8]
  assign io_vme_rd_cmd_bits_addr = tensorLoad_io_vme_rd_cmd_bits_addr; // @[TensorLoad.scala 72:8]
  assign io_vme_rd_cmd_bits_len = tensorLoad_io_vme_rd_cmd_bits_len; // @[TensorLoad.scala 72:8]
  assign io_vme_rd_cmd_bits_tag = tensorLoad_io_vme_rd_cmd_bits_tag; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_valid = tensorLoad_io_tensor_rd_0_data_valid; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_0 = tensorLoad_io_tensor_rd_0_data_bits_0_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_1 = tensorLoad_io_tensor_rd_0_data_bits_0_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_2 = tensorLoad_io_tensor_rd_0_data_bits_0_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_3 = tensorLoad_io_tensor_rd_0_data_bits_0_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_4 = tensorLoad_io_tensor_rd_0_data_bits_0_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_5 = tensorLoad_io_tensor_rd_0_data_bits_0_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_6 = tensorLoad_io_tensor_rd_0_data_bits_0_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_7 = tensorLoad_io_tensor_rd_0_data_bits_0_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_8 = tensorLoad_io_tensor_rd_0_data_bits_0_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_9 = tensorLoad_io_tensor_rd_0_data_bits_0_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_10 = tensorLoad_io_tensor_rd_0_data_bits_0_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_11 = tensorLoad_io_tensor_rd_0_data_bits_0_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_12 = tensorLoad_io_tensor_rd_0_data_bits_0_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_13 = tensorLoad_io_tensor_rd_0_data_bits_0_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_14 = tensorLoad_io_tensor_rd_0_data_bits_0_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_15 = tensorLoad_io_tensor_rd_0_data_bits_0_15; // @[TensorLoad.scala 72:8]
  assign tensorLoad_clock = clock;
  assign tensorLoad_reset = reset;
  assign tensorLoad_io_start = io_start; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_inst = io_inst; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_baddr = io_baddr; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_vme_rd_cmd_ready = io_vme_rd_cmd_ready; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_vme_rd_data_valid = io_vme_rd_data_valid; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_vme_rd_data_bits_data = io_vme_rd_data_bits_data; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_vme_rd_data_bits_tag = io_vme_rd_data_bits_tag; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_rd_0_idx_valid = io_tensor_rd_0_idx_valid; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_rd_0_idx_bits = io_tensor_rd_0_idx_bits; // @[TensorLoad.scala 72:8]
endmodule
module GenVMECmd_1(
  input          clock,
  input          reset,
  input          io_start,
  input          io_isBusy,
  input  [127:0] io_inst,
  input  [31:0]  io_baddr,
  input          io_vmeCmd_ready,
  output         io_vmeCmd_valid,
  output [31:0]  io_vmeCmd_bits_addr,
  output [3:0]   io_vmeCmd_bits_len,
  output [20:0]  io_vmeCmd_bits_tag,
  output [4:0]   io_readLen,
  output         io_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] dec_sram_offset = io_inst[25:10]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [31:0] dec_dram_offset = io_inst[57:26]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [15:0] dec_ysize = io_inst[79:64]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [15:0] dec_xsize = io_inst[95:80]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [15:0] dec_xstride = io_inst[111:96]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [3:0] dec_ypad_0 = io_inst[115:112]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [3:0] dec_xpad_0 = io_inst[123:120]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [3:0] dec_xpad_1 = io_inst[127:124]; // @[TensorLoadNarrowVME.scala 566:29]
  reg [31:0] rdCmdExtAddr; // @[TensorLoadNarrowVME.scala 568:25]
  wire [40:0] _xfer_init_addr_T = {dec_dram_offset, 9'h0}; // @[TensorLoadNarrowVME.scala 573:66]
  wire [40:0] _xfer_init_addr_T_1 = 41'hffffffff & _xfer_init_addr_T; // @[TensorLoadNarrowVME.scala 573:47]
  wire [40:0] _GEN_31 = {{9'd0}, io_baddr}; // @[TensorLoadNarrowVME.scala 573:33]
  wire [40:0] xfer_init_addr = _GEN_31 | _xfer_init_addr_T_1; // @[TensorLoadNarrowVME.scala 573:33]
  wire [31:0] _GEN_0 = rdCmdExtAddr % 32'h80; // @[TensorLoadNarrowVME.scala 577:53]
  wire [7:0] _firstMaxTransfer_T = _GEN_0[7:0]; // @[TensorLoadNarrowVME.scala 577:53]
  wire [7:0] _firstMaxTransfer_T_2 = 8'h80 - _firstMaxTransfer_T; // @[TensorLoadNarrowVME.scala 577:38]
  wire [4:0] firstMaxTransfer = _firstMaxTransfer_T_2[7:3]; // @[TensorLoadNarrowVME.scala 577:67]
  reg [5:0] rdCmdStartIdx; // @[TensorLoadNarrowVME.scala 586:26]
  reg  commandsDone; // @[TensorLoadNarrowVME.scala 588:29]
  wire [21:0] blocksReadSize = {dec_xsize, 6'h0}; // @[TensorLoadNarrowVME.scala 590:35]
  reg [21:0] blocksReadNb; // @[TensorLoadNarrowVME.scala 591:25]
  reg [31:0] rdCmdExtAddrRowBegin; // @[TensorLoadNarrowVME.scala 592:33]
  reg  newReadRow; // @[TensorLoadNarrowVME.scala 593:23]
  reg [15:0] srcRowIdx; // @[TensorLoadNarrowVME.scala 596:22]
  wire [15:0] _srcRowIdx_T_1 = srcRowIdx + 16'h1; // @[TensorLoadNarrowVME.scala 600:28]
  wire [21:0] blocksRemained = blocksReadSize - blocksReadNb; // @[TensorLoadNarrowVME.scala 628:39]
  wire [21:0] _GEN_32 = {{17'd0}, firstMaxTransfer}; // @[TensorLoadNarrowVME.scala 630:25]
  wire [21:0] _GEN_8 = blocksRemained < _GEN_32 ? blocksRemained : {{17'd0}, firstMaxTransfer}; // @[TensorLoadNarrowVME.scala 630:45 631:15 633:15]
  wire [21:0] _GEN_9 = blocksRemained < 22'h10 ? blocksRemained : 22'h10; // @[TensorLoadNarrowVME.scala 636:40 637:15 639:15]
  wire [21:0] _GEN_10 = newReadRow ? _GEN_8 : _GEN_9; // @[TensorLoadNarrowVME.scala 629:21]
  wire [4:0] readLen = _GEN_10[4:0]; // @[TensorLoadNarrowVME.scala 587:21]
  wire [21:0] _GEN_33 = {{17'd0}, readLen}; // @[TensorLoadNarrowVME.scala 621:41]
  wire [21:0] _T_8 = blocksReadSize - _GEN_33; // @[TensorLoadNarrowVME.scala 621:41]
  wire [15:0] _T_11 = dec_ysize - 16'h1; // @[TensorLoadNarrowVME.scala 621:80]
  wire  _T_14 = io_vmeCmd_ready & io_vmeCmd_valid; // @[Decoupled.scala 50:35]
  wire  stride = blocksReadNb == _T_8 & srcRowIdx != _T_11 & _T_14; // @[TensorLoadNarrowVME.scala 621:87]
  wire [21:0] nextBlRNb = blocksReadNb + _GEN_33; // @[TensorLoadNarrowVME.scala 611:34]
  wire  _GEN_2 = nextBlRNb == blocksReadSize & srcRowIdx == _T_11 | commandsDone; // @[TensorLoadNarrowVME.scala 606:16 613:74 614:20]
  wire  _GEN_4 = _T_14 ? _GEN_2 : commandsDone; // @[TensorLoadNarrowVME.scala 606:16 610:31]
  wire  _GEN_6 = io_start | stride ? 1'h0 : _GEN_4; // @[TensorLoadNarrowVME.scala 607:29 609:18]
  wire  _T_20 = ~reset; // @[TensorLoadNarrowVME.scala 627:9]
  wire [15:0] _GEN_35 = {{12'd0}, dec_xpad_0}; // @[TensorLoadNarrowVME.scala 643:30]
  wire [15:0] _totalWidth_T_1 = dec_xsize + _GEN_35; // @[TensorLoadNarrowVME.scala 643:30]
  wire [15:0] _GEN_36 = {{12'd0}, dec_xpad_1}; // @[TensorLoadNarrowVME.scala 643:43]
  wire [15:0] totalWidth = _totalWidth_T_1 + _GEN_36; // @[TensorLoadNarrowVME.scala 643:43]
  reg [19:0] currentRowIdx; // @[TensorLoadNarrowVME.scala 647:26]
  wire [19:0] _GEN_37 = {{16'd0}, dec_ypad_0}; // @[TensorLoadNarrowVME.scala 649:39]
  wire [15:0] _GEN_38 = {{12'd0}, dec_ypad_0}; // @[TensorLoadNarrowVME.scala 650:32]
  wire [15:0] _rdCmdStartIdxValid_T_2 = dec_ysize + _GEN_38; // @[TensorLoadNarrowVME.scala 650:32]
  wire [19:0] _GEN_39 = {{4'd0}, _rdCmdStartIdxValid_T_2}; // @[TensorLoadNarrowVME.scala 650:19]
  wire  _rdCmdStartIdxValid_T_3 = currentRowIdx < _GEN_39; // @[TensorLoadNarrowVME.scala 650:19]
  wire  _rdCmdStartIdxValid_T_4 = currentRowIdx >= _GEN_37 & _rdCmdStartIdxValid_T_3; // @[TensorLoadNarrowVME.scala 649:53]
  wire  _rdCmdStartIdxValid_T_5 = _rdCmdStartIdxValid_T_4 & io_isBusy; // @[TensorLoadNarrowVME.scala 650:46]
  wire  _rdCmdStartIdxValid_T_6 = ~commandsDone; // @[TensorLoadNarrowVME.scala 652:5]
  wire  rdCmdStartIdxValid = _rdCmdStartIdxValid_T_5 & _rdCmdStartIdxValid_T_6; // @[TensorLoadNarrowVME.scala 651:15]
  wire [15:0] _rdCmdStartIdx_T_1 = dec_sram_offset + _GEN_35; // @[TensorLoadNarrowVME.scala 655:38]
  wire [15:0] _GEN_42 = {{10'd0}, rdCmdStartIdx}; // @[TensorLoadNarrowVME.scala 657:36]
  wire [15:0] _rdCmdStartIdx_T_3 = _GEN_42 + totalWidth; // @[TensorLoadNarrowVME.scala 657:36]
  wire [19:0] _currentRowIdx_T_1 = currentRowIdx + 20'h1; // @[TensorLoadNarrowVME.scala 658:36]
  wire [15:0] _GEN_11 = io_isBusy & (currentRowIdx < _GEN_37 | stride) ? _rdCmdStartIdx_T_3 : {{10'd0}, rdCmdStartIdx}; // @[TensorLoadNarrowVME.scala 656:68 657:19 586:26]
  wire [15:0] _GEN_14 = io_start ? _rdCmdStartIdx_T_1 : _GEN_11; // @[TensorLoadNarrowVME.scala 653:19 655:19]
  wire  startIssueCmdRead = blocksReadNb == 22'h0 & rdCmdStartIdxValid; // @[TensorLoadNarrowVME.scala 661:29]
  wire [24:0] _memRow_T = {dec_xstride, 9'h0}; // @[TensorLoadNarrowVME.scala 672:56]
  wire [31:0] _GEN_43 = {{7'd0}, _memRow_T}; // @[TensorLoadNarrowVME.scala 672:41]
  wire [31:0] memRow = rdCmdExtAddrRowBegin + _GEN_43; // @[TensorLoadNarrowVME.scala 672:41]
  wire [7:0] _rdCmdExtAddr_T = {readLen, 3'h0}; // @[TensorLoadNarrowVME.scala 679:47]
  wire [31:0] _GEN_44 = {{24'd0}, _rdCmdExtAddr_T}; // @[TensorLoadNarrowVME.scala 679:36]
  wire [31:0] _rdCmdExtAddr_T_2 = rdCmdExtAddr + _GEN_44; // @[TensorLoadNarrowVME.scala 679:36]
  wire [31:0] _GEN_16 = stride ? memRow : _rdCmdExtAddr_T_2; // @[TensorLoadNarrowVME.scala 671:18 673:20 679:20]
  wire [31:0] _GEN_17 = stride ? memRow : rdCmdExtAddrRowBegin; // @[TensorLoadNarrowVME.scala 671:18 664:24 674:28]
  wire [31:0] _GEN_19 = _T_14 ? _GEN_16 : rdCmdExtAddr; // @[TensorLoadNarrowVME.scala 670:31 682:18]
  wire [31:0] _GEN_20 = _T_14 ? _GEN_17 : rdCmdExtAddrRowBegin; // @[TensorLoadNarrowVME.scala 664:24 670:31]
  wire  _GEN_21 = _T_14 ? stride : newReadRow; // @[TensorLoadNarrowVME.scala 670:31 683:16]
  wire [40:0] _GEN_22 = io_start ? xfer_init_addr : {{9'd0}, _GEN_19}; // @[TensorLoadNarrowVME.scala 666:19 667:18]
  wire [40:0] _GEN_23 = io_start ? xfer_init_addr : {{9'd0}, _GEN_20}; // @[TensorLoadNarrowVME.scala 666:19 668:26]
  reg [11:0] rdCmdDestBlockIdxNext; // @[TensorLoadNarrowVME.scala 700:34]
  wire [11:0] _rdCmdDestBlockIdx_T = {rdCmdStartIdx, 6'h0}; // @[TensorLoadNarrowVME.scala 710:42]
  wire [11:0] _GEN_26 = startIssueCmdRead ? _rdCmdDestBlockIdx_T : rdCmdDestBlockIdxNext; // @[TensorLoadNarrowVME.scala 702:21 709:29 710:25]
  wire [11:0] rdCmdDestBlockIdx = rdCmdStartIdxValid ? _GEN_26 : rdCmdDestBlockIdxNext; // @[TensorLoadNarrowVME.scala 702:21 707:28]
  wire [11:0] _GEN_45 = {{7'd0}, readLen}; // @[TensorLoadNarrowVME.scala 711:49]
  wire [11:0] _rdCmdDestBlockIdxNext_T_1 = rdCmdDestBlockIdx + _GEN_45; // @[TensorLoadNarrowVME.scala 711:49]
  wire [11:0] _rdCmdDestBlockIdxNext_T_3 = rdCmdDestBlockIdxNext + _GEN_45; // @[TensorLoadNarrowVME.scala 714:53]
  wire [4:0] _io_vmeCmd_bits_len_T_1 = readLen - 5'h1; // @[TensorLoadNarrowVME.scala 732:33]
  assign io_vmeCmd_valid = _rdCmdStartIdxValid_T_5 & _rdCmdStartIdxValid_T_6; // @[TensorLoadNarrowVME.scala 651:15]
  assign io_vmeCmd_bits_addr = rdCmdExtAddr; // @[TensorLoadNarrowVME.scala 731:23]
  assign io_vmeCmd_bits_len = _io_vmeCmd_bits_len_T_1[3:0]; // @[TensorLoadNarrowVME.scala 732:22]
  assign io_vmeCmd_bits_tag = {{9'd0}, rdCmdDestBlockIdx}; // @[TensorLoadNarrowVME.scala 737:22]
  assign io_readLen = _GEN_10[4:0]; // @[TensorLoadNarrowVME.scala 587:21]
  assign io_done = commandsDone; // @[TensorLoadNarrowVME.scala 739:11]
  always @(posedge clock) begin
    rdCmdExtAddr <= _GEN_22[31:0];
    rdCmdStartIdx <= _GEN_14[5:0];
    commandsDone <= reset | _GEN_6; // @[TensorLoadNarrowVME.scala 588:{29,29}]
    if (io_start | stride) begin // @[TensorLoadNarrowVME.scala 607:29]
      blocksReadNb <= 22'h0; // @[TensorLoadNarrowVME.scala 608:18]
    end else if (_T_14) begin // @[TensorLoadNarrowVME.scala 610:31]
      blocksReadNb <= nextBlRNb; // @[TensorLoadNarrowVME.scala 612:18]
    end
    rdCmdExtAddrRowBegin <= _GEN_23[31:0];
    newReadRow <= io_start | _GEN_21; // @[TensorLoadNarrowVME.scala 666:19 669:16]
    if (io_start) begin // @[TensorLoadNarrowVME.scala 597:19]
      srcRowIdx <= 16'h0; // @[TensorLoadNarrowVME.scala 598:15]
    end else if (stride) begin // @[TensorLoadNarrowVME.scala 599:23]
      srcRowIdx <= _srcRowIdx_T_1; // @[TensorLoadNarrowVME.scala 600:15]
    end
    if (io_start) begin // @[TensorLoadNarrowVME.scala 653:19]
      currentRowIdx <= 20'h0; // @[TensorLoadNarrowVME.scala 654:19]
    end else if (io_isBusy & (currentRowIdx < _GEN_37 | stride)) begin // @[TensorLoadNarrowVME.scala 656:68]
      currentRowIdx <= _currentRowIdx_T_1; // @[TensorLoadNarrowVME.scala 658:19]
    end
    if (rdCmdStartIdxValid) begin // @[TensorLoadNarrowVME.scala 707:28]
      if (startIssueCmdRead) begin // @[TensorLoadNarrowVME.scala 709:29]
        rdCmdDestBlockIdxNext <= _rdCmdDestBlockIdxNext_T_1; // @[TensorLoadNarrowVME.scala 711:28]
      end else if (_T_14) begin // @[TensorLoadNarrowVME.scala 712:33]
        rdCmdDestBlockIdxNext <= _rdCmdDestBlockIdxNext_T_3; // @[TensorLoadNarrowVME.scala 714:28]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~io_isBusy | blocksReadSize >= blocksReadNb)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorLoadNarrowVME.scala:627 assert(!io.isBusy || blocksReadSize >= blocksReadNb)// define how many block to read at this cycle\n"
            ); // @[TensorLoadNarrowVME.scala 627:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_20 & ~(~io_vmeCmd_valid | _rdCmdExtAddr_T <= _firstMaxTransfer_T_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed: -F- wgt DRAM page alignment failure. DRAM address + len overlaps mp.lenBits*memBlockSize alignment %x %x\n    at TensorLoadNarrowVME.scala:733 assert(!io.vmeCmd.valid || ((readLen << log2Ceil(mp.dataBits/8)) <= (maxTrBytes - rdCmdExtAddr %% maxTrBytes)),\n"
            ,rdCmdExtAddr,readLen); // @[TensorLoadNarrowVME.scala 733:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rdCmdExtAddr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  rdCmdStartIdx = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  commandsDone = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  blocksReadNb = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  rdCmdExtAddrRowBegin = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  newReadRow = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  srcRowIdx = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  currentRowIdx = _RAND_7[19:0];
  _RAND_8 = {1{`RANDOM}};
  rdCmdDestBlockIdxNext = _RAND_8[11:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~io_isBusy | blocksReadSize >= blocksReadNb); // @[TensorLoadNarrowVME.scala 627:9]
    end
    //
    if (_T_20) begin
      assert(~io_vmeCmd_valid | _rdCmdExtAddr_T <= _firstMaxTransfer_T_2); // @[TensorLoadNarrowVME.scala 733:9]
    end
  end
endmodule
module ReadVMEData_1(
  input         clock,
  input         reset,
  input         io_start,
  output        io_vmeData_ready,
  input         io_vmeData_valid,
  input  [20:0] io_vmeData_bits_tag,
  output [5:0]  io_idx,
  output [5:0]  io_col
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [20:0] vmeTagDecodeLast; // @[TensorLoadNarrowVME.scala 502:29]
  wire [14:0] rdDataIdx = io_vmeData_bits_tag[20:6]; // @[TensorLoadNarrowVME.scala 503:31]
  wire [5:0] rdDataCol = io_vmeData_bits_tag[5:0]; // @[TensorLoadNarrowVME.scala 504:65]
  reg [5:0] rdDataDestColNext; // @[TensorLoadNarrowVME.scala 505:30]
  reg [15:0] rdDataDestIdxNext; // @[TensorLoadNarrowVME.scala 506:30]
  reg  vmeTagDecodeLastValidNext; // @[TensorLoadNarrowVME.scala 509:42]
  wire  _T = io_vmeData_ready & io_vmeData_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_0 = _T | vmeTagDecodeLastValidNext; // @[TensorLoadNarrowVME.scala 514:31 515:27 517:27]
  wire  _T_3 = io_vmeData_bits_tag != vmeTagDecodeLast; // @[TensorLoadNarrowVME.scala 525:29]
  wire  _T_4 = vmeTagDecodeLastValidNext & _T_3; // @[TensorLoadNarrowVME.scala 524:34]
  wire  _T_5 = ~vmeTagDecodeLastValidNext | _T_4; // @[TensorLoadNarrowVME.scala 523:34]
  wire [5:0] _rdDataDestColNext_T_1 = rdDataCol + 6'h1; // @[TensorLoadNarrowVME.scala 530:38]
  wire [5:0] _rdDataDestColNext_T_3 = rdDataDestColNext + 6'h1; // @[TensorLoadNarrowVME.scala 534:46]
  wire [5:0] rdDataDestCol = _T_5 ? rdDataCol : rdDataDestColNext; // @[TensorLoadNarrowVME.scala 525:59 528:21 533:21]
  wire [15:0] _rdDataDestIdxNext_T_1 = rdDataDestIdxNext + 16'h1; // @[TensorLoadNarrowVME.scala 537:48]
  wire [15:0] rdDataDestIdx = _T_5 ? {{1'd0}, rdDataIdx} : rdDataDestIdxNext; // @[TensorLoadNarrowVME.scala 525:59 529:21 535:21]
  assign io_vmeData_ready = 1'h1; // @[TensorLoadNarrowVME.scala 498:20]
  assign io_idx = rdDataDestIdx[5:0]; // @[TensorLoadNarrowVME.scala 542:10]
  assign io_col = _T_5 ? rdDataCol : rdDataDestColNext; // @[TensorLoadNarrowVME.scala 525:59 528:21 533:21]
  always @(posedge clock) begin
    if (_T) begin // @[TensorLoadNarrowVME.scala 521:25]
      if (_T_5) begin // @[TensorLoadNarrowVME.scala 525:59]
        vmeTagDecodeLast <= io_vmeData_bits_tag; // @[TensorLoadNarrowVME.scala 527:24]
      end
    end
    if (_T) begin // @[TensorLoadNarrowVME.scala 521:25]
      if (_T_5) begin // @[TensorLoadNarrowVME.scala 525:59]
        rdDataDestColNext <= _rdDataDestColNext_T_1; // @[TensorLoadNarrowVME.scala 530:25]
      end else begin
        rdDataDestColNext <= _rdDataDestColNext_T_3; // @[TensorLoadNarrowVME.scala 534:25]
      end
    end
    if (_T) begin // @[TensorLoadNarrowVME.scala 521:25]
      if (_T_5) begin // @[TensorLoadNarrowVME.scala 525:59]
        rdDataDestIdxNext <= {{1'd0}, rdDataIdx}; // @[TensorLoadNarrowVME.scala 531:25]
      end else if (rdDataDestCol == 6'h3f) begin // @[TensorLoadNarrowVME.scala 536:54]
        rdDataDestIdxNext <= _rdDataDestIdxNext_T_1; // @[TensorLoadNarrowVME.scala 537:27]
      end
    end
    if (reset) begin // @[TensorLoadNarrowVME.scala 509:42]
      vmeTagDecodeLastValidNext <= 1'h0; // @[TensorLoadNarrowVME.scala 509:42]
    end else if (io_start) begin // @[TensorLoadNarrowVME.scala 512:18]
      vmeTagDecodeLastValidNext <= 1'h0; // @[TensorLoadNarrowVME.scala 513:27]
    end else begin
      vmeTagDecodeLastValidNext <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  vmeTagDecodeLast = _RAND_0[20:0];
  _RAND_1 = {1{`RANDOM}};
  rdDataDestColNext = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  rdDataDestIdxNext = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  vmeTagDecodeLastValidNext = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ZeroPadding_1(
  input          clock,
  input          reset,
  input          io_canWriteMem,
  input  [127:0] io_inst,
  output         io_tensorIdx_valid,
  output [5:0]   io_tensorIdx_bits,
  input          io_start,
  output         io_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] dec_sram_offset = io_inst[25:10]; // @[TensorLoadNarrowVME.scala 329:29]
  wire [15:0] dec_ysize = io_inst[79:64]; // @[TensorLoadNarrowVME.scala 329:29]
  wire [15:0] dec_xsize = io_inst[95:80]; // @[TensorLoadNarrowVME.scala 329:29]
  wire [3:0] dec_ypad_0 = io_inst[115:112]; // @[TensorLoadNarrowVME.scala 329:29]
  wire [3:0] dec_ypad_1 = io_inst[119:116]; // @[TensorLoadNarrowVME.scala 329:29]
  wire [3:0] dec_xpad_0 = io_inst[123:120]; // @[TensorLoadNarrowVME.scala 329:29]
  wire [3:0] dec_xpad_1 = io_inst[127:124]; // @[TensorLoadNarrowVME.scala 329:29]
  reg [2:0] zpState; // @[TensorLoadNarrowVME.scala 335:24]
  reg [23:0] zpColIdx; // @[TensorLoadNarrowVME.scala 337:21]
  reg [23:0] zpRowIdx; // @[TensorLoadNarrowVME.scala 340:21]
  reg [15:0] zpDestRowOffset; // @[TensorLoadNarrowVME.scala 342:28]
  wire [15:0] _GEN_35 = {{12'd0}, dec_ypad_0}; // @[TensorLoadNarrowVME.scala 349:47]
  wire [15:0] _zpLastDataRow_T_1 = _GEN_35 + dec_ysize; // @[TensorLoadNarrowVME.scala 349:47]
  wire [15:0] _zpLastDataRow_T_3 = _zpLastDataRow_T_1 - 16'h1; // @[TensorLoadNarrowVME.scala 349:59]
  wire [23:0] _GEN_36 = {{8'd0}, _zpLastDataRow_T_3}; // @[TensorLoadNarrowVME.scala 349:32]
  wire  zpLastDataRow = zpRowIdx == _GEN_36; // @[TensorLoadNarrowVME.scala 349:32]
  wire [15:0] _GEN_37 = {{12'd0}, dec_xpad_0}; // @[TensorLoadNarrowVME.scala 350:33]
  wire [15:0] _zpTopLastIdx_T_1 = _GEN_37 + dec_xsize; // @[TensorLoadNarrowVME.scala 350:33]
  wire [15:0] _GEN_38 = {{12'd0}, dec_xpad_1}; // @[TensorLoadNarrowVME.scala 350:45]
  wire [15:0] _zpTopLastIdx_T_3 = _zpTopLastIdx_T_1 + _GEN_38; // @[TensorLoadNarrowVME.scala 350:45]
  wire [15:0] zpTopLastIdx = _zpTopLastIdx_T_3 - 16'h1; // @[TensorLoadNarrowVME.scala 350:58]
  wire  _zpWideLineEnd_T = zpState == 3'h4; // @[TensorLoadNarrowVME.scala 351:32]
  wire  _zpWideLineEnd_T_1 = zpState == 3'h3; // @[TensorLoadNarrowVME.scala 351:59]
  wire [23:0] _GEN_39 = {{8'd0}, zpTopLastIdx}; // @[TensorLoadNarrowVME.scala 351:89]
  wire  _zpWideLineEnd_T_3 = zpColIdx == _GEN_39; // @[TensorLoadNarrowVME.scala 351:89]
  wire  zpWideLineEnd = (zpState == 3'h4 | zpState == 3'h3) & zpColIdx == _GEN_39; // @[TensorLoadNarrowVME.scala 351:77]
  wire [3:0] _zpNarwLineEnd_T_2 = dec_xpad_0 - 4'h1; // @[TensorLoadNarrowVME.scala 352:74]
  wire [23:0] _GEN_40 = {{20'd0}, _zpNarwLineEnd_T_2}; // @[TensorLoadNarrowVME.scala 352:59]
  wire  _zpNarwLineEnd_T_3 = zpColIdx == _GEN_40; // @[TensorLoadNarrowVME.scala 352:59]
  wire  zpNarwLineEnd = zpState == 3'h2 & zpColIdx == _GEN_40; // @[TensorLoadNarrowVME.scala 352:47]
  wire  zpFillLineEnd = zpWideLineEnd | zpNarwLineEnd; // @[TensorLoadNarrowVME.scala 353:37]
  wire  _T_1 = dec_xpad_1 != 4'h0; // @[TensorLoadNarrowVME.scala 360:43]
  wire  _T_2 = dec_xpad_0 == 4'h0 & dec_xpad_1 != 4'h0; // @[TensorLoadNarrowVME.scala 360:29]
  wire [15:0] _GEN_0 = dec_xpad_0 == 4'h0 & dec_xpad_1 != 4'h0 & dec_ypad_0 == 4'h0 ? _zpTopLastIdx_T_1 : 16'h0; // @[TensorLoadNarrowVME.scala 359:14 360:74 361:16]
  wire  _T_6 = dec_xpad_0 != 4'h0; // @[TensorLoadNarrowVME.scala 365:27]
  wire  _T_15 = dec_ypad_1 != 4'h0; // @[TensorLoadNarrowVME.scala 371:27]
  wire [2:0] _GEN_1 = dec_ypad_1 != 4'h0 ? 3'h5 : 3'h0; // @[TensorLoadNarrowVME.scala 371:36 372:15 374:15]
  wire [2:0] _GEN_2 = _T_6 & _T_1 ? 3'h4 : _GEN_1; // @[TensorLoadNarrowVME.scala 369:58 370:15]
  wire [2:0] _GEN_3 = _T_2 ? 3'h3 : _GEN_2; // @[TensorLoadNarrowVME.scala 367:58 368:15]
  wire [2:0] _GEN_4 = dec_xpad_0 != 4'h0 & dec_xpad_1 == 4'h0 ? 3'h2 : _GEN_3; // @[TensorLoadNarrowVME.scala 365:58 366:15]
  wire  _T_16 = zpState == 3'h1; // @[TensorLoadNarrowVME.scala 378:14]
  wire  _T_17 = io_canWriteMem & _T_16; // @[TensorLoadNarrowVME.scala 377:20]
  wire [3:0] _T_19 = dec_ypad_0 - 4'h1; // @[TensorLoadNarrowVME.scala 379:29]
  wire [23:0] _GEN_42 = {{20'd0}, _T_19}; // @[TensorLoadNarrowVME.scala 379:14]
  wire  _T_20 = zpRowIdx == _GEN_42; // @[TensorLoadNarrowVME.scala 379:14]
  wire  _T_21 = _T_17 & _T_20; // @[TensorLoadNarrowVME.scala 378:25]
  wire  _T_23 = _T_21 & _zpWideLineEnd_T_3; // @[TensorLoadNarrowVME.scala 379:35]
  wire [15:0] _GEN_6 = _T_2 ? _zpTopLastIdx_T_1 : 16'h0; // @[TensorLoadNarrowVME.scala 383:14 384:52 385:16]
  wire  _T_38 = zpState == 3'h5; // @[TensorLoadNarrowVME.scala 401:15]
  wire  _T_39 = zpFillLineEnd & io_canWriteMem | _T_38; // @[TensorLoadNarrowVME.scala 400:40]
  wire  _T_40 = zpLastDataRow & _T_39; // @[TensorLoadNarrowVME.scala 399:19]
  wire [23:0] _GEN_11 = _T_15 ? 24'h0 : zpColIdx; // @[TensorLoadNarrowVME.scala 344:12 405:30 406:16]
  wire [2:0] _GEN_12 = _T_15 ? 3'h6 : 3'h0; // @[TensorLoadNarrowVME.scala 405:30 407:15 409:15]
  wire  _T_42 = zpState == 3'h6; // @[TensorLoadNarrowVME.scala 413:14]
  wire  _T_43 = io_canWriteMem & _T_42; // @[TensorLoadNarrowVME.scala 412:20]
  wire [15:0] _GEN_46 = {{12'd0}, dec_ypad_1}; // @[TensorLoadNarrowVME.scala 414:41]
  wire [15:0] _T_47 = _zpLastDataRow_T_1 + _GEN_46; // @[TensorLoadNarrowVME.scala 414:41]
  wire [15:0] _T_49 = _T_47 - 16'h1; // @[TensorLoadNarrowVME.scala 414:54]
  wire [23:0] _GEN_47 = {{8'd0}, _T_49}; // @[TensorLoadNarrowVME.scala 414:14]
  wire  _T_50 = zpRowIdx == _GEN_47; // @[TensorLoadNarrowVME.scala 414:14]
  wire  _T_51 = _T_43 & _T_50; // @[TensorLoadNarrowVME.scala 413:25]
  wire  _T_53 = _T_51 & _zpWideLineEnd_T_3; // @[TensorLoadNarrowVME.scala 414:60]
  wire [23:0] _GEN_14 = _T_53 ? 24'h0 : zpColIdx; // @[TensorLoadNarrowVME.scala 344:12 415:32 418:14]
  wire [2:0] _GEN_15 = _T_53 ? 3'h0 : zpState; // @[TensorLoadNarrowVME.scala 415:32 419:13 421:13]
  wire  _GEN_16 = _T_40 | _T_53; // @[TensorLoadNarrowVME.scala 401:63 403:20]
  wire [23:0] _GEN_17 = _T_40 ? _GEN_11 : _GEN_14; // @[TensorLoadNarrowVME.scala 401:63]
  wire  _GEN_19 = _T_23 | _GEN_16; // @[TensorLoadNarrowVME.scala 380:32 381:20]
  wire [23:0] _GEN_20 = _T_23 ? {{8'd0}, _GEN_6} : _GEN_17; // @[TensorLoadNarrowVME.scala 380:32]
  wire [23:0] _GEN_24 = io_start ? {{8'd0}, _GEN_0} : _GEN_20; // @[TensorLoadNarrowVME.scala 355:18]
  wire  zpNewFillBlock = io_start ? 1'h0 : _GEN_19; // @[TensorLoadNarrowVME.scala 346:18 355:18]
  wire  isZeroPadWrite = zpState != 3'h0 & zpState != 3'h5 & io_canWriteMem; // @[TensorLoadNarrowVME.scala 424:68]
  wire [23:0] _GEN_49 = {{8'd0}, zpDestRowOffset}; // @[TensorLoadNarrowVME.scala 425:32]
  wire [23:0] _zpDestIdx_T_1 = _GEN_49 + zpColIdx; // @[TensorLoadNarrowVME.scala 425:32]
  wire  _T_62 = (_T_16 | _zpWideLineEnd_T | _zpWideLineEnd_T_1 | _T_42) & _zpWideLineEnd_T_3; // @[TensorLoadNarrowVME.scala 432:106]
  wire  _T_68 = _T_62 | zpNarwLineEnd; // @[TensorLoadNarrowVME.scala 433:34]
  wire  incrementRow = _T_68 & io_canWriteMem | _T_38; // @[TensorLoadNarrowVME.scala 434:84]
  wire [15:0] _zpDestRowOffset_T_1 = zpDestRowOffset + zpTopLastIdx; // @[TensorLoadNarrowVME.scala 437:40]
  wire [15:0] _zpDestRowOffset_T_3 = _zpDestRowOffset_T_1 + 16'h1; // @[TensorLoadNarrowVME.scala 437:55]
  wire [23:0] _zpRowIdx_T_1 = zpRowIdx + 24'h1; // @[TensorLoadNarrowVME.scala 438:26]
  wire  _T_72 = ~zpNewFillBlock; // @[TensorLoadNarrowVME.scala 440:10]
  wire [15:0] _GEN_27 = _zpWideLineEnd_T_1 ? _zpTopLastIdx_T_1 : 16'h0; // @[TensorLoadNarrowVME.scala 441:38 442:18 444:18]
  wire [23:0] _GEN_54 = {{8'd0}, dec_xsize}; // @[TensorLoadNarrowVME.scala 452:28]
  wire [23:0] _zpColIdx_T_7 = zpColIdx + _GEN_54; // @[TensorLoadNarrowVME.scala 452:28]
  wire [23:0] _zpColIdx_T_9 = _zpColIdx_T_7 + 24'h1; // @[TensorLoadNarrowVME.scala 452:40]
  wire [23:0] _zpColIdx_T_11 = zpColIdx + 24'h1; // @[TensorLoadNarrowVME.scala 455:28]
  wire [15:0] zpDestIdx = _zpDestIdx_T_1[15:0]; // @[TensorLoadNarrowVME.scala 332:23 425:13]
  assign io_tensorIdx_valid = zpState != 3'h0 & zpState != 3'h5 & io_canWriteMem; // @[TensorLoadNarrowVME.scala 424:68]
  assign io_tensorIdx_bits = zpDestIdx[5:0]; // @[TensorLoadNarrowVME.scala 460:21]
  assign io_done = zpState == 3'h0; // @[TensorLoadNarrowVME.scala 458:22]
  always @(posedge clock) begin
    if (reset) begin // @[TensorLoadNarrowVME.scala 335:24]
      zpState <= 3'h0; // @[TensorLoadNarrowVME.scala 335:24]
    end else if (io_start) begin // @[TensorLoadNarrowVME.scala 355:18]
      if (dec_ypad_0 != 4'h0) begin // @[TensorLoadNarrowVME.scala 363:30]
        zpState <= 3'h1; // @[TensorLoadNarrowVME.scala 364:15]
      end else begin
        zpState <= _GEN_4;
      end
    end else if (_T_23) begin // @[TensorLoadNarrowVME.scala 380:32]
      zpState <= _GEN_4;
    end else if (_T_40) begin // @[TensorLoadNarrowVME.scala 401:63]
      zpState <= _GEN_12;
    end else begin
      zpState <= _GEN_15;
    end
    if (isZeroPadWrite & _T_72 & ~incrementRow) begin // @[TensorLoadNarrowVME.scala 450:60]
      if (_zpWideLineEnd_T & _zpNarwLineEnd_T_3) begin // @[TensorLoadNarrowVME.scala 451:68]
        zpColIdx <= _zpColIdx_T_9; // @[TensorLoadNarrowVME.scala 452:16]
      end else begin
        zpColIdx <= _zpColIdx_T_11; // @[TensorLoadNarrowVME.scala 455:16]
      end
    end else if (incrementRow) begin // @[TensorLoadNarrowVME.scala 435:30]
      if (~zpNewFillBlock) begin // @[TensorLoadNarrowVME.scala 440:27]
        zpColIdx <= {{8'd0}, _GEN_27};
      end else begin
        zpColIdx <= _GEN_24;
      end
    end else begin
      zpColIdx <= _GEN_24;
    end
    if (incrementRow) begin // @[TensorLoadNarrowVME.scala 435:30]
      zpRowIdx <= _zpRowIdx_T_1; // @[TensorLoadNarrowVME.scala 438:14]
    end else if (io_start) begin // @[TensorLoadNarrowVME.scala 355:18]
      zpRowIdx <= 24'h0; // @[TensorLoadNarrowVME.scala 356:14]
    end
    if (incrementRow) begin // @[TensorLoadNarrowVME.scala 435:30]
      zpDestRowOffset <= _zpDestRowOffset_T_3; // @[TensorLoadNarrowVME.scala 437:21]
    end else if (io_start) begin // @[TensorLoadNarrowVME.scala 355:18]
      zpDestRowOffset <= dec_sram_offset; // @[TensorLoadNarrowVME.scala 357:21]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  zpState = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  zpColIdx = _RAND_1[23:0];
  _RAND_2 = {1{`RANDOM}};
  zpRowIdx = _RAND_2[23:0];
  _RAND_3 = {1{`RANDOM}};
  zpDestRowOffset = _RAND_3[15:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TensorLoadNarrowVME_1(
  input          clock,
  input          reset,
  input          io_start,
  output         io_done,
  input  [127:0] io_inst,
  input  [31:0]  io_baddr,
  input          io_vme_rd_cmd_ready,
  output         io_vme_rd_cmd_valid,
  output [31:0]  io_vme_rd_cmd_bits_addr,
  output [3:0]   io_vme_rd_cmd_bits_len,
  output [20:0]  io_vme_rd_cmd_bits_tag,
  output         io_vme_rd_data_ready,
  input          io_vme_rd_data_valid,
  input  [63:0]  io_vme_rd_data_bits_data,
  input  [20:0]  io_vme_rd_data_bits_tag,
  input          io_tensor_rd_0_idx_valid,
  input  [5:0]   io_tensor_rd_0_idx_bits,
  output         io_tensor_rd_0_data_valid,
  output [7:0]   io_tensor_rd_0_data_bits_0_0,
  output [7:0]   io_tensor_rd_0_data_bits_0_1,
  output [7:0]   io_tensor_rd_0_data_bits_0_2,
  output [7:0]   io_tensor_rd_0_data_bits_0_3,
  output [7:0]   io_tensor_rd_0_data_bits_0_4,
  output [7:0]   io_tensor_rd_0_data_bits_0_5,
  output [7:0]   io_tensor_rd_0_data_bits_0_6,
  output [7:0]   io_tensor_rd_0_data_bits_0_7,
  output [7:0]   io_tensor_rd_0_data_bits_0_8,
  output [7:0]   io_tensor_rd_0_data_bits_0_9,
  output [7:0]   io_tensor_rd_0_data_bits_0_10,
  output [7:0]   io_tensor_rd_0_data_bits_0_11,
  output [7:0]   io_tensor_rd_0_data_bits_0_12,
  output [7:0]   io_tensor_rd_0_data_bits_0_13,
  output [7:0]   io_tensor_rd_0_data_bits_0_14,
  output [7:0]   io_tensor_rd_0_data_bits_0_15,
  output [7:0]   io_tensor_rd_0_data_bits_1_0,
  output [7:0]   io_tensor_rd_0_data_bits_1_1,
  output [7:0]   io_tensor_rd_0_data_bits_1_2,
  output [7:0]   io_tensor_rd_0_data_bits_1_3,
  output [7:0]   io_tensor_rd_0_data_bits_1_4,
  output [7:0]   io_tensor_rd_0_data_bits_1_5,
  output [7:0]   io_tensor_rd_0_data_bits_1_6,
  output [7:0]   io_tensor_rd_0_data_bits_1_7,
  output [7:0]   io_tensor_rd_0_data_bits_1_8,
  output [7:0]   io_tensor_rd_0_data_bits_1_9,
  output [7:0]   io_tensor_rd_0_data_bits_1_10,
  output [7:0]   io_tensor_rd_0_data_bits_1_11,
  output [7:0]   io_tensor_rd_0_data_bits_1_12,
  output [7:0]   io_tensor_rd_0_data_bits_1_13,
  output [7:0]   io_tensor_rd_0_data_bits_1_14,
  output [7:0]   io_tensor_rd_0_data_bits_1_15,
  output [7:0]   io_tensor_rd_0_data_bits_2_0,
  output [7:0]   io_tensor_rd_0_data_bits_2_1,
  output [7:0]   io_tensor_rd_0_data_bits_2_2,
  output [7:0]   io_tensor_rd_0_data_bits_2_3,
  output [7:0]   io_tensor_rd_0_data_bits_2_4,
  output [7:0]   io_tensor_rd_0_data_bits_2_5,
  output [7:0]   io_tensor_rd_0_data_bits_2_6,
  output [7:0]   io_tensor_rd_0_data_bits_2_7,
  output [7:0]   io_tensor_rd_0_data_bits_2_8,
  output [7:0]   io_tensor_rd_0_data_bits_2_9,
  output [7:0]   io_tensor_rd_0_data_bits_2_10,
  output [7:0]   io_tensor_rd_0_data_bits_2_11,
  output [7:0]   io_tensor_rd_0_data_bits_2_12,
  output [7:0]   io_tensor_rd_0_data_bits_2_13,
  output [7:0]   io_tensor_rd_0_data_bits_2_14,
  output [7:0]   io_tensor_rd_0_data_bits_2_15,
  output [7:0]   io_tensor_rd_0_data_bits_3_0,
  output [7:0]   io_tensor_rd_0_data_bits_3_1,
  output [7:0]   io_tensor_rd_0_data_bits_3_2,
  output [7:0]   io_tensor_rd_0_data_bits_3_3,
  output [7:0]   io_tensor_rd_0_data_bits_3_4,
  output [7:0]   io_tensor_rd_0_data_bits_3_5,
  output [7:0]   io_tensor_rd_0_data_bits_3_6,
  output [7:0]   io_tensor_rd_0_data_bits_3_7,
  output [7:0]   io_tensor_rd_0_data_bits_3_8,
  output [7:0]   io_tensor_rd_0_data_bits_3_9,
  output [7:0]   io_tensor_rd_0_data_bits_3_10,
  output [7:0]   io_tensor_rd_0_data_bits_3_11,
  output [7:0]   io_tensor_rd_0_data_bits_3_12,
  output [7:0]   io_tensor_rd_0_data_bits_3_13,
  output [7:0]   io_tensor_rd_0_data_bits_3_14,
  output [7:0]   io_tensor_rd_0_data_bits_3_15,
  output [7:0]   io_tensor_rd_0_data_bits_4_0,
  output [7:0]   io_tensor_rd_0_data_bits_4_1,
  output [7:0]   io_tensor_rd_0_data_bits_4_2,
  output [7:0]   io_tensor_rd_0_data_bits_4_3,
  output [7:0]   io_tensor_rd_0_data_bits_4_4,
  output [7:0]   io_tensor_rd_0_data_bits_4_5,
  output [7:0]   io_tensor_rd_0_data_bits_4_6,
  output [7:0]   io_tensor_rd_0_data_bits_4_7,
  output [7:0]   io_tensor_rd_0_data_bits_4_8,
  output [7:0]   io_tensor_rd_0_data_bits_4_9,
  output [7:0]   io_tensor_rd_0_data_bits_4_10,
  output [7:0]   io_tensor_rd_0_data_bits_4_11,
  output [7:0]   io_tensor_rd_0_data_bits_4_12,
  output [7:0]   io_tensor_rd_0_data_bits_4_13,
  output [7:0]   io_tensor_rd_0_data_bits_4_14,
  output [7:0]   io_tensor_rd_0_data_bits_4_15,
  output [7:0]   io_tensor_rd_0_data_bits_5_0,
  output [7:0]   io_tensor_rd_0_data_bits_5_1,
  output [7:0]   io_tensor_rd_0_data_bits_5_2,
  output [7:0]   io_tensor_rd_0_data_bits_5_3,
  output [7:0]   io_tensor_rd_0_data_bits_5_4,
  output [7:0]   io_tensor_rd_0_data_bits_5_5,
  output [7:0]   io_tensor_rd_0_data_bits_5_6,
  output [7:0]   io_tensor_rd_0_data_bits_5_7,
  output [7:0]   io_tensor_rd_0_data_bits_5_8,
  output [7:0]   io_tensor_rd_0_data_bits_5_9,
  output [7:0]   io_tensor_rd_0_data_bits_5_10,
  output [7:0]   io_tensor_rd_0_data_bits_5_11,
  output [7:0]   io_tensor_rd_0_data_bits_5_12,
  output [7:0]   io_tensor_rd_0_data_bits_5_13,
  output [7:0]   io_tensor_rd_0_data_bits_5_14,
  output [7:0]   io_tensor_rd_0_data_bits_5_15,
  output [7:0]   io_tensor_rd_0_data_bits_6_0,
  output [7:0]   io_tensor_rd_0_data_bits_6_1,
  output [7:0]   io_tensor_rd_0_data_bits_6_2,
  output [7:0]   io_tensor_rd_0_data_bits_6_3,
  output [7:0]   io_tensor_rd_0_data_bits_6_4,
  output [7:0]   io_tensor_rd_0_data_bits_6_5,
  output [7:0]   io_tensor_rd_0_data_bits_6_6,
  output [7:0]   io_tensor_rd_0_data_bits_6_7,
  output [7:0]   io_tensor_rd_0_data_bits_6_8,
  output [7:0]   io_tensor_rd_0_data_bits_6_9,
  output [7:0]   io_tensor_rd_0_data_bits_6_10,
  output [7:0]   io_tensor_rd_0_data_bits_6_11,
  output [7:0]   io_tensor_rd_0_data_bits_6_12,
  output [7:0]   io_tensor_rd_0_data_bits_6_13,
  output [7:0]   io_tensor_rd_0_data_bits_6_14,
  output [7:0]   io_tensor_rd_0_data_bits_6_15,
  output [7:0]   io_tensor_rd_0_data_bits_7_0,
  output [7:0]   io_tensor_rd_0_data_bits_7_1,
  output [7:0]   io_tensor_rd_0_data_bits_7_2,
  output [7:0]   io_tensor_rd_0_data_bits_7_3,
  output [7:0]   io_tensor_rd_0_data_bits_7_4,
  output [7:0]   io_tensor_rd_0_data_bits_7_5,
  output [7:0]   io_tensor_rd_0_data_bits_7_6,
  output [7:0]   io_tensor_rd_0_data_bits_7_7,
  output [7:0]   io_tensor_rd_0_data_bits_7_8,
  output [7:0]   io_tensor_rd_0_data_bits_7_9,
  output [7:0]   io_tensor_rd_0_data_bits_7_10,
  output [7:0]   io_tensor_rd_0_data_bits_7_11,
  output [7:0]   io_tensor_rd_0_data_bits_7_12,
  output [7:0]   io_tensor_rd_0_data_bits_7_13,
  output [7:0]   io_tensor_rd_0_data_bits_7_14,
  output [7:0]   io_tensor_rd_0_data_bits_7_15,
  output [7:0]   io_tensor_rd_0_data_bits_8_0,
  output [7:0]   io_tensor_rd_0_data_bits_8_1,
  output [7:0]   io_tensor_rd_0_data_bits_8_2,
  output [7:0]   io_tensor_rd_0_data_bits_8_3,
  output [7:0]   io_tensor_rd_0_data_bits_8_4,
  output [7:0]   io_tensor_rd_0_data_bits_8_5,
  output [7:0]   io_tensor_rd_0_data_bits_8_6,
  output [7:0]   io_tensor_rd_0_data_bits_8_7,
  output [7:0]   io_tensor_rd_0_data_bits_8_8,
  output [7:0]   io_tensor_rd_0_data_bits_8_9,
  output [7:0]   io_tensor_rd_0_data_bits_8_10,
  output [7:0]   io_tensor_rd_0_data_bits_8_11,
  output [7:0]   io_tensor_rd_0_data_bits_8_12,
  output [7:0]   io_tensor_rd_0_data_bits_8_13,
  output [7:0]   io_tensor_rd_0_data_bits_8_14,
  output [7:0]   io_tensor_rd_0_data_bits_8_15,
  output [7:0]   io_tensor_rd_0_data_bits_9_0,
  output [7:0]   io_tensor_rd_0_data_bits_9_1,
  output [7:0]   io_tensor_rd_0_data_bits_9_2,
  output [7:0]   io_tensor_rd_0_data_bits_9_3,
  output [7:0]   io_tensor_rd_0_data_bits_9_4,
  output [7:0]   io_tensor_rd_0_data_bits_9_5,
  output [7:0]   io_tensor_rd_0_data_bits_9_6,
  output [7:0]   io_tensor_rd_0_data_bits_9_7,
  output [7:0]   io_tensor_rd_0_data_bits_9_8,
  output [7:0]   io_tensor_rd_0_data_bits_9_9,
  output [7:0]   io_tensor_rd_0_data_bits_9_10,
  output [7:0]   io_tensor_rd_0_data_bits_9_11,
  output [7:0]   io_tensor_rd_0_data_bits_9_12,
  output [7:0]   io_tensor_rd_0_data_bits_9_13,
  output [7:0]   io_tensor_rd_0_data_bits_9_14,
  output [7:0]   io_tensor_rd_0_data_bits_9_15,
  output [7:0]   io_tensor_rd_0_data_bits_10_0,
  output [7:0]   io_tensor_rd_0_data_bits_10_1,
  output [7:0]   io_tensor_rd_0_data_bits_10_2,
  output [7:0]   io_tensor_rd_0_data_bits_10_3,
  output [7:0]   io_tensor_rd_0_data_bits_10_4,
  output [7:0]   io_tensor_rd_0_data_bits_10_5,
  output [7:0]   io_tensor_rd_0_data_bits_10_6,
  output [7:0]   io_tensor_rd_0_data_bits_10_7,
  output [7:0]   io_tensor_rd_0_data_bits_10_8,
  output [7:0]   io_tensor_rd_0_data_bits_10_9,
  output [7:0]   io_tensor_rd_0_data_bits_10_10,
  output [7:0]   io_tensor_rd_0_data_bits_10_11,
  output [7:0]   io_tensor_rd_0_data_bits_10_12,
  output [7:0]   io_tensor_rd_0_data_bits_10_13,
  output [7:0]   io_tensor_rd_0_data_bits_10_14,
  output [7:0]   io_tensor_rd_0_data_bits_10_15,
  output [7:0]   io_tensor_rd_0_data_bits_11_0,
  output [7:0]   io_tensor_rd_0_data_bits_11_1,
  output [7:0]   io_tensor_rd_0_data_bits_11_2,
  output [7:0]   io_tensor_rd_0_data_bits_11_3,
  output [7:0]   io_tensor_rd_0_data_bits_11_4,
  output [7:0]   io_tensor_rd_0_data_bits_11_5,
  output [7:0]   io_tensor_rd_0_data_bits_11_6,
  output [7:0]   io_tensor_rd_0_data_bits_11_7,
  output [7:0]   io_tensor_rd_0_data_bits_11_8,
  output [7:0]   io_tensor_rd_0_data_bits_11_9,
  output [7:0]   io_tensor_rd_0_data_bits_11_10,
  output [7:0]   io_tensor_rd_0_data_bits_11_11,
  output [7:0]   io_tensor_rd_0_data_bits_11_12,
  output [7:0]   io_tensor_rd_0_data_bits_11_13,
  output [7:0]   io_tensor_rd_0_data_bits_11_14,
  output [7:0]   io_tensor_rd_0_data_bits_11_15,
  output [7:0]   io_tensor_rd_0_data_bits_12_0,
  output [7:0]   io_tensor_rd_0_data_bits_12_1,
  output [7:0]   io_tensor_rd_0_data_bits_12_2,
  output [7:0]   io_tensor_rd_0_data_bits_12_3,
  output [7:0]   io_tensor_rd_0_data_bits_12_4,
  output [7:0]   io_tensor_rd_0_data_bits_12_5,
  output [7:0]   io_tensor_rd_0_data_bits_12_6,
  output [7:0]   io_tensor_rd_0_data_bits_12_7,
  output [7:0]   io_tensor_rd_0_data_bits_12_8,
  output [7:0]   io_tensor_rd_0_data_bits_12_9,
  output [7:0]   io_tensor_rd_0_data_bits_12_10,
  output [7:0]   io_tensor_rd_0_data_bits_12_11,
  output [7:0]   io_tensor_rd_0_data_bits_12_12,
  output [7:0]   io_tensor_rd_0_data_bits_12_13,
  output [7:0]   io_tensor_rd_0_data_bits_12_14,
  output [7:0]   io_tensor_rd_0_data_bits_12_15,
  output [7:0]   io_tensor_rd_0_data_bits_13_0,
  output [7:0]   io_tensor_rd_0_data_bits_13_1,
  output [7:0]   io_tensor_rd_0_data_bits_13_2,
  output [7:0]   io_tensor_rd_0_data_bits_13_3,
  output [7:0]   io_tensor_rd_0_data_bits_13_4,
  output [7:0]   io_tensor_rd_0_data_bits_13_5,
  output [7:0]   io_tensor_rd_0_data_bits_13_6,
  output [7:0]   io_tensor_rd_0_data_bits_13_7,
  output [7:0]   io_tensor_rd_0_data_bits_13_8,
  output [7:0]   io_tensor_rd_0_data_bits_13_9,
  output [7:0]   io_tensor_rd_0_data_bits_13_10,
  output [7:0]   io_tensor_rd_0_data_bits_13_11,
  output [7:0]   io_tensor_rd_0_data_bits_13_12,
  output [7:0]   io_tensor_rd_0_data_bits_13_13,
  output [7:0]   io_tensor_rd_0_data_bits_13_14,
  output [7:0]   io_tensor_rd_0_data_bits_13_15,
  output [7:0]   io_tensor_rd_0_data_bits_14_0,
  output [7:0]   io_tensor_rd_0_data_bits_14_1,
  output [7:0]   io_tensor_rd_0_data_bits_14_2,
  output [7:0]   io_tensor_rd_0_data_bits_14_3,
  output [7:0]   io_tensor_rd_0_data_bits_14_4,
  output [7:0]   io_tensor_rd_0_data_bits_14_5,
  output [7:0]   io_tensor_rd_0_data_bits_14_6,
  output [7:0]   io_tensor_rd_0_data_bits_14_7,
  output [7:0]   io_tensor_rd_0_data_bits_14_8,
  output [7:0]   io_tensor_rd_0_data_bits_14_9,
  output [7:0]   io_tensor_rd_0_data_bits_14_10,
  output [7:0]   io_tensor_rd_0_data_bits_14_11,
  output [7:0]   io_tensor_rd_0_data_bits_14_12,
  output [7:0]   io_tensor_rd_0_data_bits_14_13,
  output [7:0]   io_tensor_rd_0_data_bits_14_14,
  output [7:0]   io_tensor_rd_0_data_bits_14_15,
  output [7:0]   io_tensor_rd_0_data_bits_15_0,
  output [7:0]   io_tensor_rd_0_data_bits_15_1,
  output [7:0]   io_tensor_rd_0_data_bits_15_2,
  output [7:0]   io_tensor_rd_0_data_bits_15_3,
  output [7:0]   io_tensor_rd_0_data_bits_15_4,
  output [7:0]   io_tensor_rd_0_data_bits_15_5,
  output [7:0]   io_tensor_rd_0_data_bits_15_6,
  output [7:0]   io_tensor_rd_0_data_bits_15_7,
  output [7:0]   io_tensor_rd_0_data_bits_15_8,
  output [7:0]   io_tensor_rd_0_data_bits_15_9,
  output [7:0]   io_tensor_rd_0_data_bits_15_10,
  output [7:0]   io_tensor_rd_0_data_bits_15_11,
  output [7:0]   io_tensor_rd_0_data_bits_15_12,
  output [7:0]   io_tensor_rd_0_data_bits_15_13,
  output [7:0]   io_tensor_rd_0_data_bits_15_14,
  output [7:0]   io_tensor_rd_0_data_bits_15_15,
  output [7:0]   io_tensor_rd_0_data_bits_16_0,
  output [7:0]   io_tensor_rd_0_data_bits_16_1,
  output [7:0]   io_tensor_rd_0_data_bits_16_2,
  output [7:0]   io_tensor_rd_0_data_bits_16_3,
  output [7:0]   io_tensor_rd_0_data_bits_16_4,
  output [7:0]   io_tensor_rd_0_data_bits_16_5,
  output [7:0]   io_tensor_rd_0_data_bits_16_6,
  output [7:0]   io_tensor_rd_0_data_bits_16_7,
  output [7:0]   io_tensor_rd_0_data_bits_16_8,
  output [7:0]   io_tensor_rd_0_data_bits_16_9,
  output [7:0]   io_tensor_rd_0_data_bits_16_10,
  output [7:0]   io_tensor_rd_0_data_bits_16_11,
  output [7:0]   io_tensor_rd_0_data_bits_16_12,
  output [7:0]   io_tensor_rd_0_data_bits_16_13,
  output [7:0]   io_tensor_rd_0_data_bits_16_14,
  output [7:0]   io_tensor_rd_0_data_bits_16_15,
  output [7:0]   io_tensor_rd_0_data_bits_17_0,
  output [7:0]   io_tensor_rd_0_data_bits_17_1,
  output [7:0]   io_tensor_rd_0_data_bits_17_2,
  output [7:0]   io_tensor_rd_0_data_bits_17_3,
  output [7:0]   io_tensor_rd_0_data_bits_17_4,
  output [7:0]   io_tensor_rd_0_data_bits_17_5,
  output [7:0]   io_tensor_rd_0_data_bits_17_6,
  output [7:0]   io_tensor_rd_0_data_bits_17_7,
  output [7:0]   io_tensor_rd_0_data_bits_17_8,
  output [7:0]   io_tensor_rd_0_data_bits_17_9,
  output [7:0]   io_tensor_rd_0_data_bits_17_10,
  output [7:0]   io_tensor_rd_0_data_bits_17_11,
  output [7:0]   io_tensor_rd_0_data_bits_17_12,
  output [7:0]   io_tensor_rd_0_data_bits_17_13,
  output [7:0]   io_tensor_rd_0_data_bits_17_14,
  output [7:0]   io_tensor_rd_0_data_bits_17_15,
  output [7:0]   io_tensor_rd_0_data_bits_18_0,
  output [7:0]   io_tensor_rd_0_data_bits_18_1,
  output [7:0]   io_tensor_rd_0_data_bits_18_2,
  output [7:0]   io_tensor_rd_0_data_bits_18_3,
  output [7:0]   io_tensor_rd_0_data_bits_18_4,
  output [7:0]   io_tensor_rd_0_data_bits_18_5,
  output [7:0]   io_tensor_rd_0_data_bits_18_6,
  output [7:0]   io_tensor_rd_0_data_bits_18_7,
  output [7:0]   io_tensor_rd_0_data_bits_18_8,
  output [7:0]   io_tensor_rd_0_data_bits_18_9,
  output [7:0]   io_tensor_rd_0_data_bits_18_10,
  output [7:0]   io_tensor_rd_0_data_bits_18_11,
  output [7:0]   io_tensor_rd_0_data_bits_18_12,
  output [7:0]   io_tensor_rd_0_data_bits_18_13,
  output [7:0]   io_tensor_rd_0_data_bits_18_14,
  output [7:0]   io_tensor_rd_0_data_bits_18_15,
  output [7:0]   io_tensor_rd_0_data_bits_19_0,
  output [7:0]   io_tensor_rd_0_data_bits_19_1,
  output [7:0]   io_tensor_rd_0_data_bits_19_2,
  output [7:0]   io_tensor_rd_0_data_bits_19_3,
  output [7:0]   io_tensor_rd_0_data_bits_19_4,
  output [7:0]   io_tensor_rd_0_data_bits_19_5,
  output [7:0]   io_tensor_rd_0_data_bits_19_6,
  output [7:0]   io_tensor_rd_0_data_bits_19_7,
  output [7:0]   io_tensor_rd_0_data_bits_19_8,
  output [7:0]   io_tensor_rd_0_data_bits_19_9,
  output [7:0]   io_tensor_rd_0_data_bits_19_10,
  output [7:0]   io_tensor_rd_0_data_bits_19_11,
  output [7:0]   io_tensor_rd_0_data_bits_19_12,
  output [7:0]   io_tensor_rd_0_data_bits_19_13,
  output [7:0]   io_tensor_rd_0_data_bits_19_14,
  output [7:0]   io_tensor_rd_0_data_bits_19_15,
  output [7:0]   io_tensor_rd_0_data_bits_20_0,
  output [7:0]   io_tensor_rd_0_data_bits_20_1,
  output [7:0]   io_tensor_rd_0_data_bits_20_2,
  output [7:0]   io_tensor_rd_0_data_bits_20_3,
  output [7:0]   io_tensor_rd_0_data_bits_20_4,
  output [7:0]   io_tensor_rd_0_data_bits_20_5,
  output [7:0]   io_tensor_rd_0_data_bits_20_6,
  output [7:0]   io_tensor_rd_0_data_bits_20_7,
  output [7:0]   io_tensor_rd_0_data_bits_20_8,
  output [7:0]   io_tensor_rd_0_data_bits_20_9,
  output [7:0]   io_tensor_rd_0_data_bits_20_10,
  output [7:0]   io_tensor_rd_0_data_bits_20_11,
  output [7:0]   io_tensor_rd_0_data_bits_20_12,
  output [7:0]   io_tensor_rd_0_data_bits_20_13,
  output [7:0]   io_tensor_rd_0_data_bits_20_14,
  output [7:0]   io_tensor_rd_0_data_bits_20_15,
  output [7:0]   io_tensor_rd_0_data_bits_21_0,
  output [7:0]   io_tensor_rd_0_data_bits_21_1,
  output [7:0]   io_tensor_rd_0_data_bits_21_2,
  output [7:0]   io_tensor_rd_0_data_bits_21_3,
  output [7:0]   io_tensor_rd_0_data_bits_21_4,
  output [7:0]   io_tensor_rd_0_data_bits_21_5,
  output [7:0]   io_tensor_rd_0_data_bits_21_6,
  output [7:0]   io_tensor_rd_0_data_bits_21_7,
  output [7:0]   io_tensor_rd_0_data_bits_21_8,
  output [7:0]   io_tensor_rd_0_data_bits_21_9,
  output [7:0]   io_tensor_rd_0_data_bits_21_10,
  output [7:0]   io_tensor_rd_0_data_bits_21_11,
  output [7:0]   io_tensor_rd_0_data_bits_21_12,
  output [7:0]   io_tensor_rd_0_data_bits_21_13,
  output [7:0]   io_tensor_rd_0_data_bits_21_14,
  output [7:0]   io_tensor_rd_0_data_bits_21_15,
  output [7:0]   io_tensor_rd_0_data_bits_22_0,
  output [7:0]   io_tensor_rd_0_data_bits_22_1,
  output [7:0]   io_tensor_rd_0_data_bits_22_2,
  output [7:0]   io_tensor_rd_0_data_bits_22_3,
  output [7:0]   io_tensor_rd_0_data_bits_22_4,
  output [7:0]   io_tensor_rd_0_data_bits_22_5,
  output [7:0]   io_tensor_rd_0_data_bits_22_6,
  output [7:0]   io_tensor_rd_0_data_bits_22_7,
  output [7:0]   io_tensor_rd_0_data_bits_22_8,
  output [7:0]   io_tensor_rd_0_data_bits_22_9,
  output [7:0]   io_tensor_rd_0_data_bits_22_10,
  output [7:0]   io_tensor_rd_0_data_bits_22_11,
  output [7:0]   io_tensor_rd_0_data_bits_22_12,
  output [7:0]   io_tensor_rd_0_data_bits_22_13,
  output [7:0]   io_tensor_rd_0_data_bits_22_14,
  output [7:0]   io_tensor_rd_0_data_bits_22_15,
  output [7:0]   io_tensor_rd_0_data_bits_23_0,
  output [7:0]   io_tensor_rd_0_data_bits_23_1,
  output [7:0]   io_tensor_rd_0_data_bits_23_2,
  output [7:0]   io_tensor_rd_0_data_bits_23_3,
  output [7:0]   io_tensor_rd_0_data_bits_23_4,
  output [7:0]   io_tensor_rd_0_data_bits_23_5,
  output [7:0]   io_tensor_rd_0_data_bits_23_6,
  output [7:0]   io_tensor_rd_0_data_bits_23_7,
  output [7:0]   io_tensor_rd_0_data_bits_23_8,
  output [7:0]   io_tensor_rd_0_data_bits_23_9,
  output [7:0]   io_tensor_rd_0_data_bits_23_10,
  output [7:0]   io_tensor_rd_0_data_bits_23_11,
  output [7:0]   io_tensor_rd_0_data_bits_23_12,
  output [7:0]   io_tensor_rd_0_data_bits_23_13,
  output [7:0]   io_tensor_rd_0_data_bits_23_14,
  output [7:0]   io_tensor_rd_0_data_bits_23_15,
  output [7:0]   io_tensor_rd_0_data_bits_24_0,
  output [7:0]   io_tensor_rd_0_data_bits_24_1,
  output [7:0]   io_tensor_rd_0_data_bits_24_2,
  output [7:0]   io_tensor_rd_0_data_bits_24_3,
  output [7:0]   io_tensor_rd_0_data_bits_24_4,
  output [7:0]   io_tensor_rd_0_data_bits_24_5,
  output [7:0]   io_tensor_rd_0_data_bits_24_6,
  output [7:0]   io_tensor_rd_0_data_bits_24_7,
  output [7:0]   io_tensor_rd_0_data_bits_24_8,
  output [7:0]   io_tensor_rd_0_data_bits_24_9,
  output [7:0]   io_tensor_rd_0_data_bits_24_10,
  output [7:0]   io_tensor_rd_0_data_bits_24_11,
  output [7:0]   io_tensor_rd_0_data_bits_24_12,
  output [7:0]   io_tensor_rd_0_data_bits_24_13,
  output [7:0]   io_tensor_rd_0_data_bits_24_14,
  output [7:0]   io_tensor_rd_0_data_bits_24_15,
  output [7:0]   io_tensor_rd_0_data_bits_25_0,
  output [7:0]   io_tensor_rd_0_data_bits_25_1,
  output [7:0]   io_tensor_rd_0_data_bits_25_2,
  output [7:0]   io_tensor_rd_0_data_bits_25_3,
  output [7:0]   io_tensor_rd_0_data_bits_25_4,
  output [7:0]   io_tensor_rd_0_data_bits_25_5,
  output [7:0]   io_tensor_rd_0_data_bits_25_6,
  output [7:0]   io_tensor_rd_0_data_bits_25_7,
  output [7:0]   io_tensor_rd_0_data_bits_25_8,
  output [7:0]   io_tensor_rd_0_data_bits_25_9,
  output [7:0]   io_tensor_rd_0_data_bits_25_10,
  output [7:0]   io_tensor_rd_0_data_bits_25_11,
  output [7:0]   io_tensor_rd_0_data_bits_25_12,
  output [7:0]   io_tensor_rd_0_data_bits_25_13,
  output [7:0]   io_tensor_rd_0_data_bits_25_14,
  output [7:0]   io_tensor_rd_0_data_bits_25_15,
  output [7:0]   io_tensor_rd_0_data_bits_26_0,
  output [7:0]   io_tensor_rd_0_data_bits_26_1,
  output [7:0]   io_tensor_rd_0_data_bits_26_2,
  output [7:0]   io_tensor_rd_0_data_bits_26_3,
  output [7:0]   io_tensor_rd_0_data_bits_26_4,
  output [7:0]   io_tensor_rd_0_data_bits_26_5,
  output [7:0]   io_tensor_rd_0_data_bits_26_6,
  output [7:0]   io_tensor_rd_0_data_bits_26_7,
  output [7:0]   io_tensor_rd_0_data_bits_26_8,
  output [7:0]   io_tensor_rd_0_data_bits_26_9,
  output [7:0]   io_tensor_rd_0_data_bits_26_10,
  output [7:0]   io_tensor_rd_0_data_bits_26_11,
  output [7:0]   io_tensor_rd_0_data_bits_26_12,
  output [7:0]   io_tensor_rd_0_data_bits_26_13,
  output [7:0]   io_tensor_rd_0_data_bits_26_14,
  output [7:0]   io_tensor_rd_0_data_bits_26_15,
  output [7:0]   io_tensor_rd_0_data_bits_27_0,
  output [7:0]   io_tensor_rd_0_data_bits_27_1,
  output [7:0]   io_tensor_rd_0_data_bits_27_2,
  output [7:0]   io_tensor_rd_0_data_bits_27_3,
  output [7:0]   io_tensor_rd_0_data_bits_27_4,
  output [7:0]   io_tensor_rd_0_data_bits_27_5,
  output [7:0]   io_tensor_rd_0_data_bits_27_6,
  output [7:0]   io_tensor_rd_0_data_bits_27_7,
  output [7:0]   io_tensor_rd_0_data_bits_27_8,
  output [7:0]   io_tensor_rd_0_data_bits_27_9,
  output [7:0]   io_tensor_rd_0_data_bits_27_10,
  output [7:0]   io_tensor_rd_0_data_bits_27_11,
  output [7:0]   io_tensor_rd_0_data_bits_27_12,
  output [7:0]   io_tensor_rd_0_data_bits_27_13,
  output [7:0]   io_tensor_rd_0_data_bits_27_14,
  output [7:0]   io_tensor_rd_0_data_bits_27_15,
  output [7:0]   io_tensor_rd_0_data_bits_28_0,
  output [7:0]   io_tensor_rd_0_data_bits_28_1,
  output [7:0]   io_tensor_rd_0_data_bits_28_2,
  output [7:0]   io_tensor_rd_0_data_bits_28_3,
  output [7:0]   io_tensor_rd_0_data_bits_28_4,
  output [7:0]   io_tensor_rd_0_data_bits_28_5,
  output [7:0]   io_tensor_rd_0_data_bits_28_6,
  output [7:0]   io_tensor_rd_0_data_bits_28_7,
  output [7:0]   io_tensor_rd_0_data_bits_28_8,
  output [7:0]   io_tensor_rd_0_data_bits_28_9,
  output [7:0]   io_tensor_rd_0_data_bits_28_10,
  output [7:0]   io_tensor_rd_0_data_bits_28_11,
  output [7:0]   io_tensor_rd_0_data_bits_28_12,
  output [7:0]   io_tensor_rd_0_data_bits_28_13,
  output [7:0]   io_tensor_rd_0_data_bits_28_14,
  output [7:0]   io_tensor_rd_0_data_bits_28_15,
  output [7:0]   io_tensor_rd_0_data_bits_29_0,
  output [7:0]   io_tensor_rd_0_data_bits_29_1,
  output [7:0]   io_tensor_rd_0_data_bits_29_2,
  output [7:0]   io_tensor_rd_0_data_bits_29_3,
  output [7:0]   io_tensor_rd_0_data_bits_29_4,
  output [7:0]   io_tensor_rd_0_data_bits_29_5,
  output [7:0]   io_tensor_rd_0_data_bits_29_6,
  output [7:0]   io_tensor_rd_0_data_bits_29_7,
  output [7:0]   io_tensor_rd_0_data_bits_29_8,
  output [7:0]   io_tensor_rd_0_data_bits_29_9,
  output [7:0]   io_tensor_rd_0_data_bits_29_10,
  output [7:0]   io_tensor_rd_0_data_bits_29_11,
  output [7:0]   io_tensor_rd_0_data_bits_29_12,
  output [7:0]   io_tensor_rd_0_data_bits_29_13,
  output [7:0]   io_tensor_rd_0_data_bits_29_14,
  output [7:0]   io_tensor_rd_0_data_bits_29_15,
  output [7:0]   io_tensor_rd_0_data_bits_30_0,
  output [7:0]   io_tensor_rd_0_data_bits_30_1,
  output [7:0]   io_tensor_rd_0_data_bits_30_2,
  output [7:0]   io_tensor_rd_0_data_bits_30_3,
  output [7:0]   io_tensor_rd_0_data_bits_30_4,
  output [7:0]   io_tensor_rd_0_data_bits_30_5,
  output [7:0]   io_tensor_rd_0_data_bits_30_6,
  output [7:0]   io_tensor_rd_0_data_bits_30_7,
  output [7:0]   io_tensor_rd_0_data_bits_30_8,
  output [7:0]   io_tensor_rd_0_data_bits_30_9,
  output [7:0]   io_tensor_rd_0_data_bits_30_10,
  output [7:0]   io_tensor_rd_0_data_bits_30_11,
  output [7:0]   io_tensor_rd_0_data_bits_30_12,
  output [7:0]   io_tensor_rd_0_data_bits_30_13,
  output [7:0]   io_tensor_rd_0_data_bits_30_14,
  output [7:0]   io_tensor_rd_0_data_bits_30_15,
  output [7:0]   io_tensor_rd_0_data_bits_31_0,
  output [7:0]   io_tensor_rd_0_data_bits_31_1,
  output [7:0]   io_tensor_rd_0_data_bits_31_2,
  output [7:0]   io_tensor_rd_0_data_bits_31_3,
  output [7:0]   io_tensor_rd_0_data_bits_31_4,
  output [7:0]   io_tensor_rd_0_data_bits_31_5,
  output [7:0]   io_tensor_rd_0_data_bits_31_6,
  output [7:0]   io_tensor_rd_0_data_bits_31_7,
  output [7:0]   io_tensor_rd_0_data_bits_31_8,
  output [7:0]   io_tensor_rd_0_data_bits_31_9,
  output [7:0]   io_tensor_rd_0_data_bits_31_10,
  output [7:0]   io_tensor_rd_0_data_bits_31_11,
  output [7:0]   io_tensor_rd_0_data_bits_31_12,
  output [7:0]   io_tensor_rd_0_data_bits_31_13,
  output [7:0]   io_tensor_rd_0_data_bits_31_14,
  output [7:0]   io_tensor_rd_0_data_bits_31_15
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_45;
  reg [63:0] _RAND_48;
  reg [63:0] _RAND_51;
  reg [63:0] _RAND_54;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_60;
  reg [63:0] _RAND_63;
  reg [63:0] _RAND_66;
  reg [63:0] _RAND_69;
  reg [63:0] _RAND_72;
  reg [63:0] _RAND_75;
  reg [63:0] _RAND_78;
  reg [63:0] _RAND_81;
  reg [63:0] _RAND_84;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_90;
  reg [63:0] _RAND_93;
  reg [63:0] _RAND_96;
  reg [63:0] _RAND_99;
  reg [63:0] _RAND_102;
  reg [63:0] _RAND_105;
  reg [63:0] _RAND_108;
  reg [63:0] _RAND_111;
  reg [63:0] _RAND_114;
  reg [63:0] _RAND_117;
  reg [63:0] _RAND_120;
  reg [63:0] _RAND_123;
  reg [63:0] _RAND_126;
  reg [63:0] _RAND_129;
  reg [63:0] _RAND_132;
  reg [63:0] _RAND_135;
  reg [63:0] _RAND_138;
  reg [63:0] _RAND_141;
  reg [63:0] _RAND_144;
  reg [63:0] _RAND_147;
  reg [63:0] _RAND_150;
  reg [63:0] _RAND_153;
  reg [63:0] _RAND_156;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_180;
  reg [63:0] _RAND_183;
  reg [63:0] _RAND_186;
  reg [63:0] _RAND_189;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [63:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [127:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
`endif // RANDOMIZE_REG_INIT
  wire  vmeCmd_clock; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_reset; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_start; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_isBusy; // @[TensorLoadNarrowVME.scala 75:23]
  wire [127:0] vmeCmd_io_inst; // @[TensorLoadNarrowVME.scala 75:23]
  wire [31:0] vmeCmd_io_baddr; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_vmeCmd_ready; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_vmeCmd_valid; // @[TensorLoadNarrowVME.scala 75:23]
  wire [31:0] vmeCmd_io_vmeCmd_bits_addr; // @[TensorLoadNarrowVME.scala 75:23]
  wire [3:0] vmeCmd_io_vmeCmd_bits_len; // @[TensorLoadNarrowVME.scala 75:23]
  wire [20:0] vmeCmd_io_vmeCmd_bits_tag; // @[TensorLoadNarrowVME.scala 75:23]
  wire [4:0] vmeCmd_io_readLen; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_done; // @[TensorLoadNarrowVME.scala 75:23]
  wire  readData_clock; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_reset; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_io_start; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_io_vmeData_ready; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_io_vmeData_valid; // @[TensorLoadNarrowVME.scala 105:24]
  wire [20:0] readData_io_vmeData_bits_tag; // @[TensorLoadNarrowVME.scala 105:24]
  wire [5:0] readData_io_idx; // @[TensorLoadNarrowVME.scala 105:24]
  wire [5:0] readData_io_col; // @[TensorLoadNarrowVME.scala 105:24]
  wire  fillPadding_clock; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_reset; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_io_canWriteMem; // @[TensorLoadNarrowVME.scala 119:27]
  wire [127:0] fillPadding_io_inst; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_io_tensorIdx_valid; // @[TensorLoadNarrowVME.scala 119:27]
  wire [5:0] fillPadding_io_tensorIdx_bits; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_io_start; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_io_done; // @[TensorLoadNarrowVME.scala 119:27]
  reg [63:0] tensorFile_0 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_0_MPORT_64_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_0_MPORT_64_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_0_MPORT_64_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_0_MPORT_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_0_MPORT_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_0_MPORT_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_0_MPORT_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_0_MPORT_64_en_pipe_0;
  reg [5:0] tensorFile_0_MPORT_64_addr_pipe_0;
  reg [63:0] tensorFile_1 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_1_MPORT_65_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_1_MPORT_65_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_1_MPORT_65_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_1_MPORT_1_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_1_MPORT_1_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_1_MPORT_1_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_1_MPORT_1_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_1_MPORT_65_en_pipe_0;
  reg [5:0] tensorFile_1_MPORT_65_addr_pipe_0;
  reg [63:0] tensorFile_2 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_2_MPORT_66_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_2_MPORT_66_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_2_MPORT_66_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_2_MPORT_2_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_2_MPORT_2_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_2_MPORT_2_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_2_MPORT_2_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_2_MPORT_66_en_pipe_0;
  reg [5:0] tensorFile_2_MPORT_66_addr_pipe_0;
  reg [63:0] tensorFile_3 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_3_MPORT_67_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_3_MPORT_67_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_3_MPORT_67_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_3_MPORT_3_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_3_MPORT_3_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_3_MPORT_3_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_3_MPORT_3_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_3_MPORT_67_en_pipe_0;
  reg [5:0] tensorFile_3_MPORT_67_addr_pipe_0;
  reg [63:0] tensorFile_4 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_4_MPORT_68_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_4_MPORT_68_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_4_MPORT_68_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_4_MPORT_4_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_4_MPORT_4_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_4_MPORT_4_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_4_MPORT_4_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_4_MPORT_68_en_pipe_0;
  reg [5:0] tensorFile_4_MPORT_68_addr_pipe_0;
  reg [63:0] tensorFile_5 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_5_MPORT_69_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_5_MPORT_69_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_5_MPORT_69_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_5_MPORT_5_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_5_MPORT_5_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_5_MPORT_5_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_5_MPORT_5_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_5_MPORT_69_en_pipe_0;
  reg [5:0] tensorFile_5_MPORT_69_addr_pipe_0;
  reg [63:0] tensorFile_6 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_6_MPORT_70_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_6_MPORT_70_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_6_MPORT_70_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_6_MPORT_6_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_6_MPORT_6_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_6_MPORT_6_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_6_MPORT_6_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_6_MPORT_70_en_pipe_0;
  reg [5:0] tensorFile_6_MPORT_70_addr_pipe_0;
  reg [63:0] tensorFile_7 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_7_MPORT_71_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_7_MPORT_71_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_7_MPORT_71_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_7_MPORT_7_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_7_MPORT_7_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_7_MPORT_7_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_7_MPORT_7_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_7_MPORT_71_en_pipe_0;
  reg [5:0] tensorFile_7_MPORT_71_addr_pipe_0;
  reg [63:0] tensorFile_8 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_8_MPORT_72_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_8_MPORT_72_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_8_MPORT_72_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_8_MPORT_8_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_8_MPORT_8_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_8_MPORT_8_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_8_MPORT_8_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_8_MPORT_72_en_pipe_0;
  reg [5:0] tensorFile_8_MPORT_72_addr_pipe_0;
  reg [63:0] tensorFile_9 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_9_MPORT_73_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_9_MPORT_73_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_9_MPORT_73_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_9_MPORT_9_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_9_MPORT_9_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_9_MPORT_9_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_9_MPORT_9_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_9_MPORT_73_en_pipe_0;
  reg [5:0] tensorFile_9_MPORT_73_addr_pipe_0;
  reg [63:0] tensorFile_10 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_10_MPORT_74_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_10_MPORT_74_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_10_MPORT_74_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_10_MPORT_10_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_10_MPORT_10_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_10_MPORT_10_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_10_MPORT_10_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_10_MPORT_74_en_pipe_0;
  reg [5:0] tensorFile_10_MPORT_74_addr_pipe_0;
  reg [63:0] tensorFile_11 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_11_MPORT_75_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_11_MPORT_75_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_11_MPORT_75_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_11_MPORT_11_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_11_MPORT_11_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_11_MPORT_11_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_11_MPORT_11_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_11_MPORT_75_en_pipe_0;
  reg [5:0] tensorFile_11_MPORT_75_addr_pipe_0;
  reg [63:0] tensorFile_12 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_12_MPORT_76_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_12_MPORT_76_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_12_MPORT_76_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_12_MPORT_12_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_12_MPORT_12_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_12_MPORT_12_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_12_MPORT_12_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_12_MPORT_76_en_pipe_0;
  reg [5:0] tensorFile_12_MPORT_76_addr_pipe_0;
  reg [63:0] tensorFile_13 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_13_MPORT_77_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_13_MPORT_77_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_13_MPORT_77_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_13_MPORT_13_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_13_MPORT_13_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_13_MPORT_13_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_13_MPORT_13_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_13_MPORT_77_en_pipe_0;
  reg [5:0] tensorFile_13_MPORT_77_addr_pipe_0;
  reg [63:0] tensorFile_14 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_14_MPORT_78_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_14_MPORT_78_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_14_MPORT_78_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_14_MPORT_14_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_14_MPORT_14_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_14_MPORT_14_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_14_MPORT_14_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_14_MPORT_78_en_pipe_0;
  reg [5:0] tensorFile_14_MPORT_78_addr_pipe_0;
  reg [63:0] tensorFile_15 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_15_MPORT_79_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_15_MPORT_79_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_15_MPORT_79_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_15_MPORT_15_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_15_MPORT_15_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_15_MPORT_15_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_15_MPORT_15_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_15_MPORT_79_en_pipe_0;
  reg [5:0] tensorFile_15_MPORT_79_addr_pipe_0;
  reg [63:0] tensorFile_16 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_16_MPORT_80_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_16_MPORT_80_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_16_MPORT_80_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_16_MPORT_16_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_16_MPORT_16_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_16_MPORT_16_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_16_MPORT_16_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_16_MPORT_80_en_pipe_0;
  reg [5:0] tensorFile_16_MPORT_80_addr_pipe_0;
  reg [63:0] tensorFile_17 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_17_MPORT_81_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_17_MPORT_81_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_17_MPORT_81_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_17_MPORT_17_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_17_MPORT_17_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_17_MPORT_17_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_17_MPORT_17_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_17_MPORT_81_en_pipe_0;
  reg [5:0] tensorFile_17_MPORT_81_addr_pipe_0;
  reg [63:0] tensorFile_18 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_18_MPORT_82_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_18_MPORT_82_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_18_MPORT_82_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_18_MPORT_18_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_18_MPORT_18_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_18_MPORT_18_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_18_MPORT_18_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_18_MPORT_82_en_pipe_0;
  reg [5:0] tensorFile_18_MPORT_82_addr_pipe_0;
  reg [63:0] tensorFile_19 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_19_MPORT_83_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_19_MPORT_83_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_19_MPORT_83_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_19_MPORT_19_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_19_MPORT_19_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_19_MPORT_19_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_19_MPORT_19_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_19_MPORT_83_en_pipe_0;
  reg [5:0] tensorFile_19_MPORT_83_addr_pipe_0;
  reg [63:0] tensorFile_20 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_20_MPORT_84_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_20_MPORT_84_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_20_MPORT_84_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_20_MPORT_20_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_20_MPORT_20_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_20_MPORT_20_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_20_MPORT_20_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_20_MPORT_84_en_pipe_0;
  reg [5:0] tensorFile_20_MPORT_84_addr_pipe_0;
  reg [63:0] tensorFile_21 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_21_MPORT_85_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_21_MPORT_85_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_21_MPORT_85_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_21_MPORT_21_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_21_MPORT_21_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_21_MPORT_21_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_21_MPORT_21_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_21_MPORT_85_en_pipe_0;
  reg [5:0] tensorFile_21_MPORT_85_addr_pipe_0;
  reg [63:0] tensorFile_22 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_22_MPORT_86_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_22_MPORT_86_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_22_MPORT_86_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_22_MPORT_22_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_22_MPORT_22_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_22_MPORT_22_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_22_MPORT_22_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_22_MPORT_86_en_pipe_0;
  reg [5:0] tensorFile_22_MPORT_86_addr_pipe_0;
  reg [63:0] tensorFile_23 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_23_MPORT_87_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_23_MPORT_87_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_23_MPORT_87_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_23_MPORT_23_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_23_MPORT_23_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_23_MPORT_23_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_23_MPORT_23_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_23_MPORT_87_en_pipe_0;
  reg [5:0] tensorFile_23_MPORT_87_addr_pipe_0;
  reg [63:0] tensorFile_24 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_24_MPORT_88_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_24_MPORT_88_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_24_MPORT_88_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_24_MPORT_24_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_24_MPORT_24_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_24_MPORT_24_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_24_MPORT_24_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_24_MPORT_88_en_pipe_0;
  reg [5:0] tensorFile_24_MPORT_88_addr_pipe_0;
  reg [63:0] tensorFile_25 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_25_MPORT_89_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_25_MPORT_89_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_25_MPORT_89_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_25_MPORT_25_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_25_MPORT_25_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_25_MPORT_25_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_25_MPORT_25_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_25_MPORT_89_en_pipe_0;
  reg [5:0] tensorFile_25_MPORT_89_addr_pipe_0;
  reg [63:0] tensorFile_26 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_26_MPORT_90_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_26_MPORT_90_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_26_MPORT_90_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_26_MPORT_26_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_26_MPORT_26_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_26_MPORT_26_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_26_MPORT_26_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_26_MPORT_90_en_pipe_0;
  reg [5:0] tensorFile_26_MPORT_90_addr_pipe_0;
  reg [63:0] tensorFile_27 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_27_MPORT_91_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_27_MPORT_91_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_27_MPORT_91_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_27_MPORT_27_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_27_MPORT_27_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_27_MPORT_27_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_27_MPORT_27_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_27_MPORT_91_en_pipe_0;
  reg [5:0] tensorFile_27_MPORT_91_addr_pipe_0;
  reg [63:0] tensorFile_28 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_28_MPORT_92_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_28_MPORT_92_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_28_MPORT_92_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_28_MPORT_28_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_28_MPORT_28_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_28_MPORT_28_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_28_MPORT_28_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_28_MPORT_92_en_pipe_0;
  reg [5:0] tensorFile_28_MPORT_92_addr_pipe_0;
  reg [63:0] tensorFile_29 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_29_MPORT_93_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_29_MPORT_93_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_29_MPORT_93_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_29_MPORT_29_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_29_MPORT_29_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_29_MPORT_29_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_29_MPORT_29_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_29_MPORT_93_en_pipe_0;
  reg [5:0] tensorFile_29_MPORT_93_addr_pipe_0;
  reg [63:0] tensorFile_30 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_30_MPORT_94_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_30_MPORT_94_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_30_MPORT_94_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_30_MPORT_30_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_30_MPORT_30_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_30_MPORT_30_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_30_MPORT_30_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_30_MPORT_94_en_pipe_0;
  reg [5:0] tensorFile_30_MPORT_94_addr_pipe_0;
  reg [63:0] tensorFile_31 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_31_MPORT_95_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_31_MPORT_95_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_31_MPORT_95_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_31_MPORT_31_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_31_MPORT_31_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_31_MPORT_31_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_31_MPORT_31_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_31_MPORT_95_en_pipe_0;
  reg [5:0] tensorFile_31_MPORT_95_addr_pipe_0;
  reg [63:0] tensorFile_32 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_32_MPORT_96_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_32_MPORT_96_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_32_MPORT_96_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_32_MPORT_32_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_32_MPORT_32_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_32_MPORT_32_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_32_MPORT_32_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_32_MPORT_96_en_pipe_0;
  reg [5:0] tensorFile_32_MPORT_96_addr_pipe_0;
  reg [63:0] tensorFile_33 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_33_MPORT_97_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_33_MPORT_97_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_33_MPORT_97_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_33_MPORT_33_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_33_MPORT_33_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_33_MPORT_33_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_33_MPORT_33_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_33_MPORT_97_en_pipe_0;
  reg [5:0] tensorFile_33_MPORT_97_addr_pipe_0;
  reg [63:0] tensorFile_34 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_34_MPORT_98_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_34_MPORT_98_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_34_MPORT_98_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_34_MPORT_34_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_34_MPORT_34_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_34_MPORT_34_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_34_MPORT_34_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_34_MPORT_98_en_pipe_0;
  reg [5:0] tensorFile_34_MPORT_98_addr_pipe_0;
  reg [63:0] tensorFile_35 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_35_MPORT_99_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_35_MPORT_99_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_35_MPORT_99_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_35_MPORT_35_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_35_MPORT_35_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_35_MPORT_35_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_35_MPORT_35_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_35_MPORT_99_en_pipe_0;
  reg [5:0] tensorFile_35_MPORT_99_addr_pipe_0;
  reg [63:0] tensorFile_36 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_36_MPORT_100_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_36_MPORT_100_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_36_MPORT_100_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_36_MPORT_36_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_36_MPORT_36_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_36_MPORT_36_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_36_MPORT_36_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_36_MPORT_100_en_pipe_0;
  reg [5:0] tensorFile_36_MPORT_100_addr_pipe_0;
  reg [63:0] tensorFile_37 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_37_MPORT_101_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_37_MPORT_101_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_37_MPORT_101_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_37_MPORT_37_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_37_MPORT_37_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_37_MPORT_37_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_37_MPORT_37_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_37_MPORT_101_en_pipe_0;
  reg [5:0] tensorFile_37_MPORT_101_addr_pipe_0;
  reg [63:0] tensorFile_38 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_38_MPORT_102_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_38_MPORT_102_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_38_MPORT_102_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_38_MPORT_38_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_38_MPORT_38_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_38_MPORT_38_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_38_MPORT_38_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_38_MPORT_102_en_pipe_0;
  reg [5:0] tensorFile_38_MPORT_102_addr_pipe_0;
  reg [63:0] tensorFile_39 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_39_MPORT_103_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_39_MPORT_103_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_39_MPORT_103_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_39_MPORT_39_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_39_MPORT_39_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_39_MPORT_39_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_39_MPORT_39_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_39_MPORT_103_en_pipe_0;
  reg [5:0] tensorFile_39_MPORT_103_addr_pipe_0;
  reg [63:0] tensorFile_40 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_40_MPORT_104_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_40_MPORT_104_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_40_MPORT_104_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_40_MPORT_40_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_40_MPORT_40_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_40_MPORT_40_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_40_MPORT_40_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_40_MPORT_104_en_pipe_0;
  reg [5:0] tensorFile_40_MPORT_104_addr_pipe_0;
  reg [63:0] tensorFile_41 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_41_MPORT_105_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_41_MPORT_105_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_41_MPORT_105_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_41_MPORT_41_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_41_MPORT_41_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_41_MPORT_41_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_41_MPORT_41_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_41_MPORT_105_en_pipe_0;
  reg [5:0] tensorFile_41_MPORT_105_addr_pipe_0;
  reg [63:0] tensorFile_42 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_42_MPORT_106_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_42_MPORT_106_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_42_MPORT_106_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_42_MPORT_42_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_42_MPORT_42_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_42_MPORT_42_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_42_MPORT_42_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_42_MPORT_106_en_pipe_0;
  reg [5:0] tensorFile_42_MPORT_106_addr_pipe_0;
  reg [63:0] tensorFile_43 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_43_MPORT_107_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_43_MPORT_107_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_43_MPORT_107_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_43_MPORT_43_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_43_MPORT_43_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_43_MPORT_43_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_43_MPORT_43_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_43_MPORT_107_en_pipe_0;
  reg [5:0] tensorFile_43_MPORT_107_addr_pipe_0;
  reg [63:0] tensorFile_44 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_44_MPORT_108_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_44_MPORT_108_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_44_MPORT_108_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_44_MPORT_44_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_44_MPORT_44_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_44_MPORT_44_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_44_MPORT_44_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_44_MPORT_108_en_pipe_0;
  reg [5:0] tensorFile_44_MPORT_108_addr_pipe_0;
  reg [63:0] tensorFile_45 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_45_MPORT_109_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_45_MPORT_109_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_45_MPORT_109_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_45_MPORT_45_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_45_MPORT_45_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_45_MPORT_45_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_45_MPORT_45_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_45_MPORT_109_en_pipe_0;
  reg [5:0] tensorFile_45_MPORT_109_addr_pipe_0;
  reg [63:0] tensorFile_46 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_46_MPORT_110_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_46_MPORT_110_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_46_MPORT_110_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_46_MPORT_46_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_46_MPORT_46_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_46_MPORT_46_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_46_MPORT_46_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_46_MPORT_110_en_pipe_0;
  reg [5:0] tensorFile_46_MPORT_110_addr_pipe_0;
  reg [63:0] tensorFile_47 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_47_MPORT_111_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_47_MPORT_111_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_47_MPORT_111_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_47_MPORT_47_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_47_MPORT_47_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_47_MPORT_47_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_47_MPORT_47_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_47_MPORT_111_en_pipe_0;
  reg [5:0] tensorFile_47_MPORT_111_addr_pipe_0;
  reg [63:0] tensorFile_48 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_48_MPORT_112_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_48_MPORT_112_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_48_MPORT_112_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_48_MPORT_48_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_48_MPORT_48_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_48_MPORT_48_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_48_MPORT_48_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_48_MPORT_112_en_pipe_0;
  reg [5:0] tensorFile_48_MPORT_112_addr_pipe_0;
  reg [63:0] tensorFile_49 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_49_MPORT_113_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_49_MPORT_113_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_49_MPORT_113_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_49_MPORT_49_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_49_MPORT_49_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_49_MPORT_49_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_49_MPORT_49_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_49_MPORT_113_en_pipe_0;
  reg [5:0] tensorFile_49_MPORT_113_addr_pipe_0;
  reg [63:0] tensorFile_50 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_50_MPORT_114_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_50_MPORT_114_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_50_MPORT_114_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_50_MPORT_50_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_50_MPORT_50_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_50_MPORT_50_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_50_MPORT_50_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_50_MPORT_114_en_pipe_0;
  reg [5:0] tensorFile_50_MPORT_114_addr_pipe_0;
  reg [63:0] tensorFile_51 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_51_MPORT_115_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_51_MPORT_115_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_51_MPORT_115_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_51_MPORT_51_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_51_MPORT_51_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_51_MPORT_51_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_51_MPORT_51_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_51_MPORT_115_en_pipe_0;
  reg [5:0] tensorFile_51_MPORT_115_addr_pipe_0;
  reg [63:0] tensorFile_52 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_52_MPORT_116_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_52_MPORT_116_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_52_MPORT_116_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_52_MPORT_52_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_52_MPORT_52_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_52_MPORT_52_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_52_MPORT_52_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_52_MPORT_116_en_pipe_0;
  reg [5:0] tensorFile_52_MPORT_116_addr_pipe_0;
  reg [63:0] tensorFile_53 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_53_MPORT_117_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_53_MPORT_117_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_53_MPORT_117_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_53_MPORT_53_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_53_MPORT_53_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_53_MPORT_53_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_53_MPORT_53_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_53_MPORT_117_en_pipe_0;
  reg [5:0] tensorFile_53_MPORT_117_addr_pipe_0;
  reg [63:0] tensorFile_54 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_54_MPORT_118_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_54_MPORT_118_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_54_MPORT_118_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_54_MPORT_54_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_54_MPORT_54_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_54_MPORT_54_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_54_MPORT_54_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_54_MPORT_118_en_pipe_0;
  reg [5:0] tensorFile_54_MPORT_118_addr_pipe_0;
  reg [63:0] tensorFile_55 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_55_MPORT_119_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_55_MPORT_119_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_55_MPORT_119_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_55_MPORT_55_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_55_MPORT_55_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_55_MPORT_55_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_55_MPORT_55_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_55_MPORT_119_en_pipe_0;
  reg [5:0] tensorFile_55_MPORT_119_addr_pipe_0;
  reg [63:0] tensorFile_56 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_56_MPORT_120_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_56_MPORT_120_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_56_MPORT_120_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_56_MPORT_56_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_56_MPORT_56_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_56_MPORT_56_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_56_MPORT_56_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_56_MPORT_120_en_pipe_0;
  reg [5:0] tensorFile_56_MPORT_120_addr_pipe_0;
  reg [63:0] tensorFile_57 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_57_MPORT_121_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_57_MPORT_121_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_57_MPORT_121_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_57_MPORT_57_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_57_MPORT_57_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_57_MPORT_57_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_57_MPORT_57_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_57_MPORT_121_en_pipe_0;
  reg [5:0] tensorFile_57_MPORT_121_addr_pipe_0;
  reg [63:0] tensorFile_58 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_58_MPORT_122_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_58_MPORT_122_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_58_MPORT_122_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_58_MPORT_58_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_58_MPORT_58_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_58_MPORT_58_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_58_MPORT_58_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_58_MPORT_122_en_pipe_0;
  reg [5:0] tensorFile_58_MPORT_122_addr_pipe_0;
  reg [63:0] tensorFile_59 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_59_MPORT_123_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_59_MPORT_123_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_59_MPORT_123_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_59_MPORT_59_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_59_MPORT_59_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_59_MPORT_59_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_59_MPORT_59_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_59_MPORT_123_en_pipe_0;
  reg [5:0] tensorFile_59_MPORT_123_addr_pipe_0;
  reg [63:0] tensorFile_60 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_60_MPORT_124_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_60_MPORT_124_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_60_MPORT_124_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_60_MPORT_60_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_60_MPORT_60_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_60_MPORT_60_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_60_MPORT_60_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_60_MPORT_124_en_pipe_0;
  reg [5:0] tensorFile_60_MPORT_124_addr_pipe_0;
  reg [63:0] tensorFile_61 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_61_MPORT_125_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_61_MPORT_125_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_61_MPORT_125_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_61_MPORT_61_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_61_MPORT_61_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_61_MPORT_61_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_61_MPORT_61_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_61_MPORT_125_en_pipe_0;
  reg [5:0] tensorFile_61_MPORT_125_addr_pipe_0;
  reg [63:0] tensorFile_62 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_62_MPORT_126_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_62_MPORT_126_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_62_MPORT_126_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_62_MPORT_62_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_62_MPORT_62_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_62_MPORT_62_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_62_MPORT_62_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_62_MPORT_126_en_pipe_0;
  reg [5:0] tensorFile_62_MPORT_126_addr_pipe_0;
  reg [63:0] tensorFile_63 [0:63]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_63_MPORT_127_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_63_MPORT_127_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_63_MPORT_127_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_63_MPORT_63_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [5:0] tensorFile_63_MPORT_63_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_63_MPORT_63_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_63_MPORT_63_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_63_MPORT_127_en_pipe_0;
  reg [5:0] tensorFile_63_MPORT_127_addr_pipe_0;
  reg  state; // @[TensorLoadNarrowVME.scala 54:22]
  reg [11:0] blocksInFlight; // @[TensorLoadNarrowVME.scala 87:27]
  wire  loadDone = blocksInFlight == 12'h0 & vmeCmd_io_done & state; // @[TensorLoadNarrowVME.scala 292:57]
  wire  localDone = loadDone & fillPadding_io_done; // @[TensorLoadNarrowVME.scala 293:25]
  wire  _GEN_0 = localDone ? 1'h0 : state; // @[TensorLoadNarrowVME.scala 61:25 62:11 54:22]
  wire  _GEN_1 = io_start | _GEN_0; // @[TensorLoadNarrowVME.scala 59:18 60:11]
  reg [63:0] vmeDataBitsPipe_data; // @[TensorLoadNarrowVME.scala 67:32]
  reg [20:0] vmeDataBitsPipe_tag; // @[TensorLoadNarrowVME.scala 67:32]
  reg  vmeDataValidPipe; // @[TensorLoadNarrowVME.scala 68:33]
  reg  vmeDataReadyPipe; // @[TensorLoadNarrowVME.scala 69:33]
  wire  vmeDataFirePipe = vmeDataValidPipe & vmeDataReadyPipe; // @[TensorLoadNarrowVME.scala 70:42]
  wire  _T = io_vme_rd_cmd_ready & io_vme_rd_cmd_valid; // @[Decoupled.scala 50:35]
  wire  _T_1 = state & _T; // @[TensorLoadNarrowVME.scala 90:21]
  wire  _T_3 = state & _T & ~vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 90:43]
  wire [11:0] _GEN_394 = {{7'd0}, vmeCmd_io_readLen}; // @[TensorLoadNarrowVME.scala 91:38]
  wire [11:0] _blocksInFlight_T_1 = blocksInFlight + _GEN_394; // @[TensorLoadNarrowVME.scala 91:38]
  wire  _T_6 = _T_1 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 92:43]
  wire [11:0] _blocksInFlight_T_5 = _blocksInFlight_T_1 - 12'h1; // @[TensorLoadNarrowVME.scala 93:48]
  wire  _T_10 = state & ~_T & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 94:44]
  wire  _T_13 = ~reset; // @[TensorLoadNarrowVME.scala 95:11]
  wire [11:0] _blocksInFlight_T_7 = blocksInFlight - 12'h1; // @[TensorLoadNarrowVME.scala 96:38]
  reg [127:0] fillPadding_io_inst_REG; // @[TensorLoadNarrowVME.scala 121:33]
  reg  fillPadding_io_start_REG; // @[TensorLoadNarrowVME.scala 122:34]
  wire [5:0] waddrTensInstrTmp = fillPadding_io_tensorIdx_valid ? fillPadding_io_tensorIdx_bits : readData_io_idx; // @[TensorLoadNarrowVME.scala 166:30]
  wire  _waddr_0_T = ~state; // @[TensorLoadNarrowVME.scala 186:27]
  wire  wenTensInstr_0 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h0 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_1 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h1 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_2 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h2 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_3 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h3 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_4 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h4 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_5 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h5 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_6 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h6 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_7 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h7 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_8 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h8 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_9 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h9 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_10 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'ha & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_11 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'hb & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_12 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'hc & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_13 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'hd & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_14 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'he & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_15 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'hf & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_16 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h10 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_17 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h11 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_18 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h12 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_19 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h13 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_20 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h14 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_21 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h15 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_22 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h16 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_23 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h17 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_24 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h18 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_25 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h19 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_26 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h1a & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_27 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h1b & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_28 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h1c & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_29 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h1d & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_30 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h1e & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_31 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h1f & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_32 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h20 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_33 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h21 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_34 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h22 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_35 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h23 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_36 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h24 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_37 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h25 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_38 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h26 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_39 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h27 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_40 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h28 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_41 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h29 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_42 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h2a & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_43 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h2b & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_44 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h2c & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_45 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h2d & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_46 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h2e & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_47 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h2f & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_48 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h30 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_49 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h31 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_50 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h32 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_51 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h33 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_52 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h34 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_53 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h35 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_54 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h36 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_55 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h37 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_56 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h38 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_57 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h39 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_58 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h3a & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_59 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h3b & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_60 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h3c & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_61 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h3d & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_62 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h3e & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_63 = fillPadding_io_tensorIdx_valid | readData_io_col == 6'h3f & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire [63:0] wdataTensInstr_0 = fillPadding_io_tensorIdx_valid ? 64'h0 : vmeDataBitsPipe_data; // @[TensorLoadNarrowVME.scala 234:29]
  reg  rvalid; // @[Reg.scala 28:20]
  wire [63:0] _WIRE_64_1 = tensorFile_1_MPORT_65_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_0 = tensorFile_0_MPORT_64_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_3 = tensorFile_3_MPORT_67_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_2 = tensorFile_2_MPORT_66_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_5 = tensorFile_5_MPORT_69_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_4 = tensorFile_4_MPORT_68_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_7 = tensorFile_7_MPORT_71_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_6 = tensorFile_6_MPORT_70_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [511:0] lo_lo_lo = {_WIRE_64_7,_WIRE_64_6,_WIRE_64_5,_WIRE_64_4,_WIRE_64_3,_WIRE_64_2,_WIRE_64_1,_WIRE_64_0}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_64_9 = tensorFile_9_MPORT_73_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_8 = tensorFile_8_MPORT_72_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_11 = tensorFile_11_MPORT_75_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_10 = tensorFile_10_MPORT_74_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_13 = tensorFile_13_MPORT_77_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_12 = tensorFile_12_MPORT_76_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_15 = tensorFile_15_MPORT_79_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_14 = tensorFile_14_MPORT_78_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [1023:0] lo_lo = {_WIRE_64_15,_WIRE_64_14,_WIRE_64_13,_WIRE_64_12,_WIRE_64_11,_WIRE_64_10,_WIRE_64_9,_WIRE_64_8,
    lo_lo_lo}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_64_17 = tensorFile_17_MPORT_81_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_16 = tensorFile_16_MPORT_80_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_19 = tensorFile_19_MPORT_83_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_18 = tensorFile_18_MPORT_82_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_21 = tensorFile_21_MPORT_85_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_20 = tensorFile_20_MPORT_84_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_23 = tensorFile_23_MPORT_87_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_22 = tensorFile_22_MPORT_86_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [511:0] lo_hi_lo = {_WIRE_64_23,_WIRE_64_22,_WIRE_64_21,_WIRE_64_20,_WIRE_64_19,_WIRE_64_18,_WIRE_64_17,
    _WIRE_64_16}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_64_25 = tensorFile_25_MPORT_89_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_24 = tensorFile_24_MPORT_88_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_27 = tensorFile_27_MPORT_91_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_26 = tensorFile_26_MPORT_90_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_29 = tensorFile_29_MPORT_93_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_28 = tensorFile_28_MPORT_92_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_31 = tensorFile_31_MPORT_95_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_30 = tensorFile_30_MPORT_94_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [2047:0] lo = {_WIRE_64_31,_WIRE_64_30,_WIRE_64_29,_WIRE_64_28,_WIRE_64_27,_WIRE_64_26,_WIRE_64_25,_WIRE_64_24,
    lo_hi_lo,lo_lo}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_64_33 = tensorFile_33_MPORT_97_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_32 = tensorFile_32_MPORT_96_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_35 = tensorFile_35_MPORT_99_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_34 = tensorFile_34_MPORT_98_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_37 = tensorFile_37_MPORT_101_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_36 = tensorFile_36_MPORT_100_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_39 = tensorFile_39_MPORT_103_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_38 = tensorFile_38_MPORT_102_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [511:0] hi_lo_lo = {_WIRE_64_39,_WIRE_64_38,_WIRE_64_37,_WIRE_64_36,_WIRE_64_35,_WIRE_64_34,_WIRE_64_33,
    _WIRE_64_32}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_64_41 = tensorFile_41_MPORT_105_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_40 = tensorFile_40_MPORT_104_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_43 = tensorFile_43_MPORT_107_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_42 = tensorFile_42_MPORT_106_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_45 = tensorFile_45_MPORT_109_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_44 = tensorFile_44_MPORT_108_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_47 = tensorFile_47_MPORT_111_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_46 = tensorFile_46_MPORT_110_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [1023:0] hi_lo = {_WIRE_64_47,_WIRE_64_46,_WIRE_64_45,_WIRE_64_44,_WIRE_64_43,_WIRE_64_42,_WIRE_64_41,_WIRE_64_40
    ,hi_lo_lo}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_64_49 = tensorFile_49_MPORT_113_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_48 = tensorFile_48_MPORT_112_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_51 = tensorFile_51_MPORT_115_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_50 = tensorFile_50_MPORT_114_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_53 = tensorFile_53_MPORT_117_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_52 = tensorFile_52_MPORT_116_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_55 = tensorFile_55_MPORT_119_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_54 = tensorFile_54_MPORT_118_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [511:0] hi_hi_lo = {_WIRE_64_55,_WIRE_64_54,_WIRE_64_53,_WIRE_64_52,_WIRE_64_51,_WIRE_64_50,_WIRE_64_49,
    _WIRE_64_48}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_64_57 = tensorFile_57_MPORT_121_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_56 = tensorFile_56_MPORT_120_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_59 = tensorFile_59_MPORT_123_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_58 = tensorFile_58_MPORT_122_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_61 = tensorFile_61_MPORT_125_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_60 = tensorFile_60_MPORT_124_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_63 = tensorFile_63_MPORT_127_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_64_62 = tensorFile_62_MPORT_126_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [2047:0] hi = {_WIRE_64_63,_WIRE_64_62,_WIRE_64_61,_WIRE_64_60,_WIRE_64_59,_WIRE_64_58,_WIRE_64_57,_WIRE_64_56,
    hi_hi_lo,hi_lo}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [4095:0] _T_148 = {hi,lo}; // @[TensorLoadNarrowVME.scala 288:18]
  GenVMECmd_1 vmeCmd ( // @[TensorLoadNarrowVME.scala 75:23]
    .clock(vmeCmd_clock),
    .reset(vmeCmd_reset),
    .io_start(vmeCmd_io_start),
    .io_isBusy(vmeCmd_io_isBusy),
    .io_inst(vmeCmd_io_inst),
    .io_baddr(vmeCmd_io_baddr),
    .io_vmeCmd_ready(vmeCmd_io_vmeCmd_ready),
    .io_vmeCmd_valid(vmeCmd_io_vmeCmd_valid),
    .io_vmeCmd_bits_addr(vmeCmd_io_vmeCmd_bits_addr),
    .io_vmeCmd_bits_len(vmeCmd_io_vmeCmd_bits_len),
    .io_vmeCmd_bits_tag(vmeCmd_io_vmeCmd_bits_tag),
    .io_readLen(vmeCmd_io_readLen),
    .io_done(vmeCmd_io_done)
  );
  ReadVMEData_1 readData ( // @[TensorLoadNarrowVME.scala 105:24]
    .clock(readData_clock),
    .reset(readData_reset),
    .io_start(readData_io_start),
    .io_vmeData_ready(readData_io_vmeData_ready),
    .io_vmeData_valid(readData_io_vmeData_valid),
    .io_vmeData_bits_tag(readData_io_vmeData_bits_tag),
    .io_idx(readData_io_idx),
    .io_col(readData_io_col)
  );
  ZeroPadding_1 fillPadding ( // @[TensorLoadNarrowVME.scala 119:27]
    .clock(fillPadding_clock),
    .reset(fillPadding_reset),
    .io_canWriteMem(fillPadding_io_canWriteMem),
    .io_inst(fillPadding_io_inst),
    .io_tensorIdx_valid(fillPadding_io_tensorIdx_valid),
    .io_tensorIdx_bits(fillPadding_io_tensorIdx_bits),
    .io_start(fillPadding_io_start),
    .io_done(fillPadding_io_done)
  );
  assign tensorFile_0_MPORT_64_en = tensorFile_0_MPORT_64_en_pipe_0;
  assign tensorFile_0_MPORT_64_addr = tensorFile_0_MPORT_64_addr_pipe_0;
  assign tensorFile_0_MPORT_64_data = tensorFile_0[tensorFile_0_MPORT_64_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_0_MPORT_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_0_MPORT_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_0_MPORT_mask = 1'h1;
  assign tensorFile_0_MPORT_en = _waddr_0_T ? 1'h0 : wenTensInstr_0;
  assign tensorFile_1_MPORT_65_en = tensorFile_1_MPORT_65_en_pipe_0;
  assign tensorFile_1_MPORT_65_addr = tensorFile_1_MPORT_65_addr_pipe_0;
  assign tensorFile_1_MPORT_65_data = tensorFile_1[tensorFile_1_MPORT_65_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_1_MPORT_1_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_1_MPORT_1_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_1_MPORT_1_mask = 1'h1;
  assign tensorFile_1_MPORT_1_en = _waddr_0_T ? 1'h0 : wenTensInstr_1;
  assign tensorFile_2_MPORT_66_en = tensorFile_2_MPORT_66_en_pipe_0;
  assign tensorFile_2_MPORT_66_addr = tensorFile_2_MPORT_66_addr_pipe_0;
  assign tensorFile_2_MPORT_66_data = tensorFile_2[tensorFile_2_MPORT_66_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_2_MPORT_2_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_2_MPORT_2_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_2_MPORT_2_mask = 1'h1;
  assign tensorFile_2_MPORT_2_en = _waddr_0_T ? 1'h0 : wenTensInstr_2;
  assign tensorFile_3_MPORT_67_en = tensorFile_3_MPORT_67_en_pipe_0;
  assign tensorFile_3_MPORT_67_addr = tensorFile_3_MPORT_67_addr_pipe_0;
  assign tensorFile_3_MPORT_67_data = tensorFile_3[tensorFile_3_MPORT_67_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_3_MPORT_3_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_3_MPORT_3_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_3_MPORT_3_mask = 1'h1;
  assign tensorFile_3_MPORT_3_en = _waddr_0_T ? 1'h0 : wenTensInstr_3;
  assign tensorFile_4_MPORT_68_en = tensorFile_4_MPORT_68_en_pipe_0;
  assign tensorFile_4_MPORT_68_addr = tensorFile_4_MPORT_68_addr_pipe_0;
  assign tensorFile_4_MPORT_68_data = tensorFile_4[tensorFile_4_MPORT_68_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_4_MPORT_4_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_4_MPORT_4_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_4_MPORT_4_mask = 1'h1;
  assign tensorFile_4_MPORT_4_en = _waddr_0_T ? 1'h0 : wenTensInstr_4;
  assign tensorFile_5_MPORT_69_en = tensorFile_5_MPORT_69_en_pipe_0;
  assign tensorFile_5_MPORT_69_addr = tensorFile_5_MPORT_69_addr_pipe_0;
  assign tensorFile_5_MPORT_69_data = tensorFile_5[tensorFile_5_MPORT_69_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_5_MPORT_5_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_5_MPORT_5_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_5_MPORT_5_mask = 1'h1;
  assign tensorFile_5_MPORT_5_en = _waddr_0_T ? 1'h0 : wenTensInstr_5;
  assign tensorFile_6_MPORT_70_en = tensorFile_6_MPORT_70_en_pipe_0;
  assign tensorFile_6_MPORT_70_addr = tensorFile_6_MPORT_70_addr_pipe_0;
  assign tensorFile_6_MPORT_70_data = tensorFile_6[tensorFile_6_MPORT_70_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_6_MPORT_6_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_6_MPORT_6_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_6_MPORT_6_mask = 1'h1;
  assign tensorFile_6_MPORT_6_en = _waddr_0_T ? 1'h0 : wenTensInstr_6;
  assign tensorFile_7_MPORT_71_en = tensorFile_7_MPORT_71_en_pipe_0;
  assign tensorFile_7_MPORT_71_addr = tensorFile_7_MPORT_71_addr_pipe_0;
  assign tensorFile_7_MPORT_71_data = tensorFile_7[tensorFile_7_MPORT_71_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_7_MPORT_7_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_7_MPORT_7_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_7_MPORT_7_mask = 1'h1;
  assign tensorFile_7_MPORT_7_en = _waddr_0_T ? 1'h0 : wenTensInstr_7;
  assign tensorFile_8_MPORT_72_en = tensorFile_8_MPORT_72_en_pipe_0;
  assign tensorFile_8_MPORT_72_addr = tensorFile_8_MPORT_72_addr_pipe_0;
  assign tensorFile_8_MPORT_72_data = tensorFile_8[tensorFile_8_MPORT_72_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_8_MPORT_8_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_8_MPORT_8_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_8_MPORT_8_mask = 1'h1;
  assign tensorFile_8_MPORT_8_en = _waddr_0_T ? 1'h0 : wenTensInstr_8;
  assign tensorFile_9_MPORT_73_en = tensorFile_9_MPORT_73_en_pipe_0;
  assign tensorFile_9_MPORT_73_addr = tensorFile_9_MPORT_73_addr_pipe_0;
  assign tensorFile_9_MPORT_73_data = tensorFile_9[tensorFile_9_MPORT_73_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_9_MPORT_9_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_9_MPORT_9_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_9_MPORT_9_mask = 1'h1;
  assign tensorFile_9_MPORT_9_en = _waddr_0_T ? 1'h0 : wenTensInstr_9;
  assign tensorFile_10_MPORT_74_en = tensorFile_10_MPORT_74_en_pipe_0;
  assign tensorFile_10_MPORT_74_addr = tensorFile_10_MPORT_74_addr_pipe_0;
  assign tensorFile_10_MPORT_74_data = tensorFile_10[tensorFile_10_MPORT_74_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_10_MPORT_10_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_10_MPORT_10_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_10_MPORT_10_mask = 1'h1;
  assign tensorFile_10_MPORT_10_en = _waddr_0_T ? 1'h0 : wenTensInstr_10;
  assign tensorFile_11_MPORT_75_en = tensorFile_11_MPORT_75_en_pipe_0;
  assign tensorFile_11_MPORT_75_addr = tensorFile_11_MPORT_75_addr_pipe_0;
  assign tensorFile_11_MPORT_75_data = tensorFile_11[tensorFile_11_MPORT_75_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_11_MPORT_11_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_11_MPORT_11_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_11_MPORT_11_mask = 1'h1;
  assign tensorFile_11_MPORT_11_en = _waddr_0_T ? 1'h0 : wenTensInstr_11;
  assign tensorFile_12_MPORT_76_en = tensorFile_12_MPORT_76_en_pipe_0;
  assign tensorFile_12_MPORT_76_addr = tensorFile_12_MPORT_76_addr_pipe_0;
  assign tensorFile_12_MPORT_76_data = tensorFile_12[tensorFile_12_MPORT_76_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_12_MPORT_12_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_12_MPORT_12_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_12_MPORT_12_mask = 1'h1;
  assign tensorFile_12_MPORT_12_en = _waddr_0_T ? 1'h0 : wenTensInstr_12;
  assign tensorFile_13_MPORT_77_en = tensorFile_13_MPORT_77_en_pipe_0;
  assign tensorFile_13_MPORT_77_addr = tensorFile_13_MPORT_77_addr_pipe_0;
  assign tensorFile_13_MPORT_77_data = tensorFile_13[tensorFile_13_MPORT_77_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_13_MPORT_13_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_13_MPORT_13_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_13_MPORT_13_mask = 1'h1;
  assign tensorFile_13_MPORT_13_en = _waddr_0_T ? 1'h0 : wenTensInstr_13;
  assign tensorFile_14_MPORT_78_en = tensorFile_14_MPORT_78_en_pipe_0;
  assign tensorFile_14_MPORT_78_addr = tensorFile_14_MPORT_78_addr_pipe_0;
  assign tensorFile_14_MPORT_78_data = tensorFile_14[tensorFile_14_MPORT_78_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_14_MPORT_14_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_14_MPORT_14_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_14_MPORT_14_mask = 1'h1;
  assign tensorFile_14_MPORT_14_en = _waddr_0_T ? 1'h0 : wenTensInstr_14;
  assign tensorFile_15_MPORT_79_en = tensorFile_15_MPORT_79_en_pipe_0;
  assign tensorFile_15_MPORT_79_addr = tensorFile_15_MPORT_79_addr_pipe_0;
  assign tensorFile_15_MPORT_79_data = tensorFile_15[tensorFile_15_MPORT_79_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_15_MPORT_15_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_15_MPORT_15_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_15_MPORT_15_mask = 1'h1;
  assign tensorFile_15_MPORT_15_en = _waddr_0_T ? 1'h0 : wenTensInstr_15;
  assign tensorFile_16_MPORT_80_en = tensorFile_16_MPORT_80_en_pipe_0;
  assign tensorFile_16_MPORT_80_addr = tensorFile_16_MPORT_80_addr_pipe_0;
  assign tensorFile_16_MPORT_80_data = tensorFile_16[tensorFile_16_MPORT_80_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_16_MPORT_16_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_16_MPORT_16_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_16_MPORT_16_mask = 1'h1;
  assign tensorFile_16_MPORT_16_en = _waddr_0_T ? 1'h0 : wenTensInstr_16;
  assign tensorFile_17_MPORT_81_en = tensorFile_17_MPORT_81_en_pipe_0;
  assign tensorFile_17_MPORT_81_addr = tensorFile_17_MPORT_81_addr_pipe_0;
  assign tensorFile_17_MPORT_81_data = tensorFile_17[tensorFile_17_MPORT_81_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_17_MPORT_17_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_17_MPORT_17_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_17_MPORT_17_mask = 1'h1;
  assign tensorFile_17_MPORT_17_en = _waddr_0_T ? 1'h0 : wenTensInstr_17;
  assign tensorFile_18_MPORT_82_en = tensorFile_18_MPORT_82_en_pipe_0;
  assign tensorFile_18_MPORT_82_addr = tensorFile_18_MPORT_82_addr_pipe_0;
  assign tensorFile_18_MPORT_82_data = tensorFile_18[tensorFile_18_MPORT_82_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_18_MPORT_18_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_18_MPORT_18_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_18_MPORT_18_mask = 1'h1;
  assign tensorFile_18_MPORT_18_en = _waddr_0_T ? 1'h0 : wenTensInstr_18;
  assign tensorFile_19_MPORT_83_en = tensorFile_19_MPORT_83_en_pipe_0;
  assign tensorFile_19_MPORT_83_addr = tensorFile_19_MPORT_83_addr_pipe_0;
  assign tensorFile_19_MPORT_83_data = tensorFile_19[tensorFile_19_MPORT_83_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_19_MPORT_19_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_19_MPORT_19_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_19_MPORT_19_mask = 1'h1;
  assign tensorFile_19_MPORT_19_en = _waddr_0_T ? 1'h0 : wenTensInstr_19;
  assign tensorFile_20_MPORT_84_en = tensorFile_20_MPORT_84_en_pipe_0;
  assign tensorFile_20_MPORT_84_addr = tensorFile_20_MPORT_84_addr_pipe_0;
  assign tensorFile_20_MPORT_84_data = tensorFile_20[tensorFile_20_MPORT_84_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_20_MPORT_20_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_20_MPORT_20_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_20_MPORT_20_mask = 1'h1;
  assign tensorFile_20_MPORT_20_en = _waddr_0_T ? 1'h0 : wenTensInstr_20;
  assign tensorFile_21_MPORT_85_en = tensorFile_21_MPORT_85_en_pipe_0;
  assign tensorFile_21_MPORT_85_addr = tensorFile_21_MPORT_85_addr_pipe_0;
  assign tensorFile_21_MPORT_85_data = tensorFile_21[tensorFile_21_MPORT_85_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_21_MPORT_21_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_21_MPORT_21_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_21_MPORT_21_mask = 1'h1;
  assign tensorFile_21_MPORT_21_en = _waddr_0_T ? 1'h0 : wenTensInstr_21;
  assign tensorFile_22_MPORT_86_en = tensorFile_22_MPORT_86_en_pipe_0;
  assign tensorFile_22_MPORT_86_addr = tensorFile_22_MPORT_86_addr_pipe_0;
  assign tensorFile_22_MPORT_86_data = tensorFile_22[tensorFile_22_MPORT_86_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_22_MPORT_22_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_22_MPORT_22_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_22_MPORT_22_mask = 1'h1;
  assign tensorFile_22_MPORT_22_en = _waddr_0_T ? 1'h0 : wenTensInstr_22;
  assign tensorFile_23_MPORT_87_en = tensorFile_23_MPORT_87_en_pipe_0;
  assign tensorFile_23_MPORT_87_addr = tensorFile_23_MPORT_87_addr_pipe_0;
  assign tensorFile_23_MPORT_87_data = tensorFile_23[tensorFile_23_MPORT_87_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_23_MPORT_23_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_23_MPORT_23_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_23_MPORT_23_mask = 1'h1;
  assign tensorFile_23_MPORT_23_en = _waddr_0_T ? 1'h0 : wenTensInstr_23;
  assign tensorFile_24_MPORT_88_en = tensorFile_24_MPORT_88_en_pipe_0;
  assign tensorFile_24_MPORT_88_addr = tensorFile_24_MPORT_88_addr_pipe_0;
  assign tensorFile_24_MPORT_88_data = tensorFile_24[tensorFile_24_MPORT_88_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_24_MPORT_24_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_24_MPORT_24_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_24_MPORT_24_mask = 1'h1;
  assign tensorFile_24_MPORT_24_en = _waddr_0_T ? 1'h0 : wenTensInstr_24;
  assign tensorFile_25_MPORT_89_en = tensorFile_25_MPORT_89_en_pipe_0;
  assign tensorFile_25_MPORT_89_addr = tensorFile_25_MPORT_89_addr_pipe_0;
  assign tensorFile_25_MPORT_89_data = tensorFile_25[tensorFile_25_MPORT_89_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_25_MPORT_25_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_25_MPORT_25_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_25_MPORT_25_mask = 1'h1;
  assign tensorFile_25_MPORT_25_en = _waddr_0_T ? 1'h0 : wenTensInstr_25;
  assign tensorFile_26_MPORT_90_en = tensorFile_26_MPORT_90_en_pipe_0;
  assign tensorFile_26_MPORT_90_addr = tensorFile_26_MPORT_90_addr_pipe_0;
  assign tensorFile_26_MPORT_90_data = tensorFile_26[tensorFile_26_MPORT_90_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_26_MPORT_26_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_26_MPORT_26_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_26_MPORT_26_mask = 1'h1;
  assign tensorFile_26_MPORT_26_en = _waddr_0_T ? 1'h0 : wenTensInstr_26;
  assign tensorFile_27_MPORT_91_en = tensorFile_27_MPORT_91_en_pipe_0;
  assign tensorFile_27_MPORT_91_addr = tensorFile_27_MPORT_91_addr_pipe_0;
  assign tensorFile_27_MPORT_91_data = tensorFile_27[tensorFile_27_MPORT_91_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_27_MPORT_27_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_27_MPORT_27_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_27_MPORT_27_mask = 1'h1;
  assign tensorFile_27_MPORT_27_en = _waddr_0_T ? 1'h0 : wenTensInstr_27;
  assign tensorFile_28_MPORT_92_en = tensorFile_28_MPORT_92_en_pipe_0;
  assign tensorFile_28_MPORT_92_addr = tensorFile_28_MPORT_92_addr_pipe_0;
  assign tensorFile_28_MPORT_92_data = tensorFile_28[tensorFile_28_MPORT_92_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_28_MPORT_28_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_28_MPORT_28_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_28_MPORT_28_mask = 1'h1;
  assign tensorFile_28_MPORT_28_en = _waddr_0_T ? 1'h0 : wenTensInstr_28;
  assign tensorFile_29_MPORT_93_en = tensorFile_29_MPORT_93_en_pipe_0;
  assign tensorFile_29_MPORT_93_addr = tensorFile_29_MPORT_93_addr_pipe_0;
  assign tensorFile_29_MPORT_93_data = tensorFile_29[tensorFile_29_MPORT_93_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_29_MPORT_29_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_29_MPORT_29_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_29_MPORT_29_mask = 1'h1;
  assign tensorFile_29_MPORT_29_en = _waddr_0_T ? 1'h0 : wenTensInstr_29;
  assign tensorFile_30_MPORT_94_en = tensorFile_30_MPORT_94_en_pipe_0;
  assign tensorFile_30_MPORT_94_addr = tensorFile_30_MPORT_94_addr_pipe_0;
  assign tensorFile_30_MPORT_94_data = tensorFile_30[tensorFile_30_MPORT_94_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_30_MPORT_30_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_30_MPORT_30_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_30_MPORT_30_mask = 1'h1;
  assign tensorFile_30_MPORT_30_en = _waddr_0_T ? 1'h0 : wenTensInstr_30;
  assign tensorFile_31_MPORT_95_en = tensorFile_31_MPORT_95_en_pipe_0;
  assign tensorFile_31_MPORT_95_addr = tensorFile_31_MPORT_95_addr_pipe_0;
  assign tensorFile_31_MPORT_95_data = tensorFile_31[tensorFile_31_MPORT_95_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_31_MPORT_31_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_31_MPORT_31_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_31_MPORT_31_mask = 1'h1;
  assign tensorFile_31_MPORT_31_en = _waddr_0_T ? 1'h0 : wenTensInstr_31;
  assign tensorFile_32_MPORT_96_en = tensorFile_32_MPORT_96_en_pipe_0;
  assign tensorFile_32_MPORT_96_addr = tensorFile_32_MPORT_96_addr_pipe_0;
  assign tensorFile_32_MPORT_96_data = tensorFile_32[tensorFile_32_MPORT_96_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_32_MPORT_32_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_32_MPORT_32_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_32_MPORT_32_mask = 1'h1;
  assign tensorFile_32_MPORT_32_en = _waddr_0_T ? 1'h0 : wenTensInstr_32;
  assign tensorFile_33_MPORT_97_en = tensorFile_33_MPORT_97_en_pipe_0;
  assign tensorFile_33_MPORT_97_addr = tensorFile_33_MPORT_97_addr_pipe_0;
  assign tensorFile_33_MPORT_97_data = tensorFile_33[tensorFile_33_MPORT_97_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_33_MPORT_33_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_33_MPORT_33_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_33_MPORT_33_mask = 1'h1;
  assign tensorFile_33_MPORT_33_en = _waddr_0_T ? 1'h0 : wenTensInstr_33;
  assign tensorFile_34_MPORT_98_en = tensorFile_34_MPORT_98_en_pipe_0;
  assign tensorFile_34_MPORT_98_addr = tensorFile_34_MPORT_98_addr_pipe_0;
  assign tensorFile_34_MPORT_98_data = tensorFile_34[tensorFile_34_MPORT_98_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_34_MPORT_34_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_34_MPORT_34_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_34_MPORT_34_mask = 1'h1;
  assign tensorFile_34_MPORT_34_en = _waddr_0_T ? 1'h0 : wenTensInstr_34;
  assign tensorFile_35_MPORT_99_en = tensorFile_35_MPORT_99_en_pipe_0;
  assign tensorFile_35_MPORT_99_addr = tensorFile_35_MPORT_99_addr_pipe_0;
  assign tensorFile_35_MPORT_99_data = tensorFile_35[tensorFile_35_MPORT_99_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_35_MPORT_35_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_35_MPORT_35_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_35_MPORT_35_mask = 1'h1;
  assign tensorFile_35_MPORT_35_en = _waddr_0_T ? 1'h0 : wenTensInstr_35;
  assign tensorFile_36_MPORT_100_en = tensorFile_36_MPORT_100_en_pipe_0;
  assign tensorFile_36_MPORT_100_addr = tensorFile_36_MPORT_100_addr_pipe_0;
  assign tensorFile_36_MPORT_100_data = tensorFile_36[tensorFile_36_MPORT_100_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_36_MPORT_36_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_36_MPORT_36_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_36_MPORT_36_mask = 1'h1;
  assign tensorFile_36_MPORT_36_en = _waddr_0_T ? 1'h0 : wenTensInstr_36;
  assign tensorFile_37_MPORT_101_en = tensorFile_37_MPORT_101_en_pipe_0;
  assign tensorFile_37_MPORT_101_addr = tensorFile_37_MPORT_101_addr_pipe_0;
  assign tensorFile_37_MPORT_101_data = tensorFile_37[tensorFile_37_MPORT_101_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_37_MPORT_37_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_37_MPORT_37_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_37_MPORT_37_mask = 1'h1;
  assign tensorFile_37_MPORT_37_en = _waddr_0_T ? 1'h0 : wenTensInstr_37;
  assign tensorFile_38_MPORT_102_en = tensorFile_38_MPORT_102_en_pipe_0;
  assign tensorFile_38_MPORT_102_addr = tensorFile_38_MPORT_102_addr_pipe_0;
  assign tensorFile_38_MPORT_102_data = tensorFile_38[tensorFile_38_MPORT_102_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_38_MPORT_38_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_38_MPORT_38_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_38_MPORT_38_mask = 1'h1;
  assign tensorFile_38_MPORT_38_en = _waddr_0_T ? 1'h0 : wenTensInstr_38;
  assign tensorFile_39_MPORT_103_en = tensorFile_39_MPORT_103_en_pipe_0;
  assign tensorFile_39_MPORT_103_addr = tensorFile_39_MPORT_103_addr_pipe_0;
  assign tensorFile_39_MPORT_103_data = tensorFile_39[tensorFile_39_MPORT_103_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_39_MPORT_39_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_39_MPORT_39_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_39_MPORT_39_mask = 1'h1;
  assign tensorFile_39_MPORT_39_en = _waddr_0_T ? 1'h0 : wenTensInstr_39;
  assign tensorFile_40_MPORT_104_en = tensorFile_40_MPORT_104_en_pipe_0;
  assign tensorFile_40_MPORT_104_addr = tensorFile_40_MPORT_104_addr_pipe_0;
  assign tensorFile_40_MPORT_104_data = tensorFile_40[tensorFile_40_MPORT_104_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_40_MPORT_40_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_40_MPORT_40_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_40_MPORT_40_mask = 1'h1;
  assign tensorFile_40_MPORT_40_en = _waddr_0_T ? 1'h0 : wenTensInstr_40;
  assign tensorFile_41_MPORT_105_en = tensorFile_41_MPORT_105_en_pipe_0;
  assign tensorFile_41_MPORT_105_addr = tensorFile_41_MPORT_105_addr_pipe_0;
  assign tensorFile_41_MPORT_105_data = tensorFile_41[tensorFile_41_MPORT_105_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_41_MPORT_41_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_41_MPORT_41_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_41_MPORT_41_mask = 1'h1;
  assign tensorFile_41_MPORT_41_en = _waddr_0_T ? 1'h0 : wenTensInstr_41;
  assign tensorFile_42_MPORT_106_en = tensorFile_42_MPORT_106_en_pipe_0;
  assign tensorFile_42_MPORT_106_addr = tensorFile_42_MPORT_106_addr_pipe_0;
  assign tensorFile_42_MPORT_106_data = tensorFile_42[tensorFile_42_MPORT_106_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_42_MPORT_42_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_42_MPORT_42_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_42_MPORT_42_mask = 1'h1;
  assign tensorFile_42_MPORT_42_en = _waddr_0_T ? 1'h0 : wenTensInstr_42;
  assign tensorFile_43_MPORT_107_en = tensorFile_43_MPORT_107_en_pipe_0;
  assign tensorFile_43_MPORT_107_addr = tensorFile_43_MPORT_107_addr_pipe_0;
  assign tensorFile_43_MPORT_107_data = tensorFile_43[tensorFile_43_MPORT_107_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_43_MPORT_43_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_43_MPORT_43_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_43_MPORT_43_mask = 1'h1;
  assign tensorFile_43_MPORT_43_en = _waddr_0_T ? 1'h0 : wenTensInstr_43;
  assign tensorFile_44_MPORT_108_en = tensorFile_44_MPORT_108_en_pipe_0;
  assign tensorFile_44_MPORT_108_addr = tensorFile_44_MPORT_108_addr_pipe_0;
  assign tensorFile_44_MPORT_108_data = tensorFile_44[tensorFile_44_MPORT_108_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_44_MPORT_44_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_44_MPORT_44_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_44_MPORT_44_mask = 1'h1;
  assign tensorFile_44_MPORT_44_en = _waddr_0_T ? 1'h0 : wenTensInstr_44;
  assign tensorFile_45_MPORT_109_en = tensorFile_45_MPORT_109_en_pipe_0;
  assign tensorFile_45_MPORT_109_addr = tensorFile_45_MPORT_109_addr_pipe_0;
  assign tensorFile_45_MPORT_109_data = tensorFile_45[tensorFile_45_MPORT_109_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_45_MPORT_45_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_45_MPORT_45_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_45_MPORT_45_mask = 1'h1;
  assign tensorFile_45_MPORT_45_en = _waddr_0_T ? 1'h0 : wenTensInstr_45;
  assign tensorFile_46_MPORT_110_en = tensorFile_46_MPORT_110_en_pipe_0;
  assign tensorFile_46_MPORT_110_addr = tensorFile_46_MPORT_110_addr_pipe_0;
  assign tensorFile_46_MPORT_110_data = tensorFile_46[tensorFile_46_MPORT_110_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_46_MPORT_46_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_46_MPORT_46_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_46_MPORT_46_mask = 1'h1;
  assign tensorFile_46_MPORT_46_en = _waddr_0_T ? 1'h0 : wenTensInstr_46;
  assign tensorFile_47_MPORT_111_en = tensorFile_47_MPORT_111_en_pipe_0;
  assign tensorFile_47_MPORT_111_addr = tensorFile_47_MPORT_111_addr_pipe_0;
  assign tensorFile_47_MPORT_111_data = tensorFile_47[tensorFile_47_MPORT_111_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_47_MPORT_47_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_47_MPORT_47_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_47_MPORT_47_mask = 1'h1;
  assign tensorFile_47_MPORT_47_en = _waddr_0_T ? 1'h0 : wenTensInstr_47;
  assign tensorFile_48_MPORT_112_en = tensorFile_48_MPORT_112_en_pipe_0;
  assign tensorFile_48_MPORT_112_addr = tensorFile_48_MPORT_112_addr_pipe_0;
  assign tensorFile_48_MPORT_112_data = tensorFile_48[tensorFile_48_MPORT_112_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_48_MPORT_48_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_48_MPORT_48_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_48_MPORT_48_mask = 1'h1;
  assign tensorFile_48_MPORT_48_en = _waddr_0_T ? 1'h0 : wenTensInstr_48;
  assign tensorFile_49_MPORT_113_en = tensorFile_49_MPORT_113_en_pipe_0;
  assign tensorFile_49_MPORT_113_addr = tensorFile_49_MPORT_113_addr_pipe_0;
  assign tensorFile_49_MPORT_113_data = tensorFile_49[tensorFile_49_MPORT_113_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_49_MPORT_49_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_49_MPORT_49_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_49_MPORT_49_mask = 1'h1;
  assign tensorFile_49_MPORT_49_en = _waddr_0_T ? 1'h0 : wenTensInstr_49;
  assign tensorFile_50_MPORT_114_en = tensorFile_50_MPORT_114_en_pipe_0;
  assign tensorFile_50_MPORT_114_addr = tensorFile_50_MPORT_114_addr_pipe_0;
  assign tensorFile_50_MPORT_114_data = tensorFile_50[tensorFile_50_MPORT_114_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_50_MPORT_50_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_50_MPORT_50_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_50_MPORT_50_mask = 1'h1;
  assign tensorFile_50_MPORT_50_en = _waddr_0_T ? 1'h0 : wenTensInstr_50;
  assign tensorFile_51_MPORT_115_en = tensorFile_51_MPORT_115_en_pipe_0;
  assign tensorFile_51_MPORT_115_addr = tensorFile_51_MPORT_115_addr_pipe_0;
  assign tensorFile_51_MPORT_115_data = tensorFile_51[tensorFile_51_MPORT_115_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_51_MPORT_51_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_51_MPORT_51_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_51_MPORT_51_mask = 1'h1;
  assign tensorFile_51_MPORT_51_en = _waddr_0_T ? 1'h0 : wenTensInstr_51;
  assign tensorFile_52_MPORT_116_en = tensorFile_52_MPORT_116_en_pipe_0;
  assign tensorFile_52_MPORT_116_addr = tensorFile_52_MPORT_116_addr_pipe_0;
  assign tensorFile_52_MPORT_116_data = tensorFile_52[tensorFile_52_MPORT_116_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_52_MPORT_52_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_52_MPORT_52_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_52_MPORT_52_mask = 1'h1;
  assign tensorFile_52_MPORT_52_en = _waddr_0_T ? 1'h0 : wenTensInstr_52;
  assign tensorFile_53_MPORT_117_en = tensorFile_53_MPORT_117_en_pipe_0;
  assign tensorFile_53_MPORT_117_addr = tensorFile_53_MPORT_117_addr_pipe_0;
  assign tensorFile_53_MPORT_117_data = tensorFile_53[tensorFile_53_MPORT_117_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_53_MPORT_53_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_53_MPORT_53_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_53_MPORT_53_mask = 1'h1;
  assign tensorFile_53_MPORT_53_en = _waddr_0_T ? 1'h0 : wenTensInstr_53;
  assign tensorFile_54_MPORT_118_en = tensorFile_54_MPORT_118_en_pipe_0;
  assign tensorFile_54_MPORT_118_addr = tensorFile_54_MPORT_118_addr_pipe_0;
  assign tensorFile_54_MPORT_118_data = tensorFile_54[tensorFile_54_MPORT_118_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_54_MPORT_54_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_54_MPORT_54_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_54_MPORT_54_mask = 1'h1;
  assign tensorFile_54_MPORT_54_en = _waddr_0_T ? 1'h0 : wenTensInstr_54;
  assign tensorFile_55_MPORT_119_en = tensorFile_55_MPORT_119_en_pipe_0;
  assign tensorFile_55_MPORT_119_addr = tensorFile_55_MPORT_119_addr_pipe_0;
  assign tensorFile_55_MPORT_119_data = tensorFile_55[tensorFile_55_MPORT_119_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_55_MPORT_55_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_55_MPORT_55_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_55_MPORT_55_mask = 1'h1;
  assign tensorFile_55_MPORT_55_en = _waddr_0_T ? 1'h0 : wenTensInstr_55;
  assign tensorFile_56_MPORT_120_en = tensorFile_56_MPORT_120_en_pipe_0;
  assign tensorFile_56_MPORT_120_addr = tensorFile_56_MPORT_120_addr_pipe_0;
  assign tensorFile_56_MPORT_120_data = tensorFile_56[tensorFile_56_MPORT_120_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_56_MPORT_56_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_56_MPORT_56_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_56_MPORT_56_mask = 1'h1;
  assign tensorFile_56_MPORT_56_en = _waddr_0_T ? 1'h0 : wenTensInstr_56;
  assign tensorFile_57_MPORT_121_en = tensorFile_57_MPORT_121_en_pipe_0;
  assign tensorFile_57_MPORT_121_addr = tensorFile_57_MPORT_121_addr_pipe_0;
  assign tensorFile_57_MPORT_121_data = tensorFile_57[tensorFile_57_MPORT_121_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_57_MPORT_57_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_57_MPORT_57_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_57_MPORT_57_mask = 1'h1;
  assign tensorFile_57_MPORT_57_en = _waddr_0_T ? 1'h0 : wenTensInstr_57;
  assign tensorFile_58_MPORT_122_en = tensorFile_58_MPORT_122_en_pipe_0;
  assign tensorFile_58_MPORT_122_addr = tensorFile_58_MPORT_122_addr_pipe_0;
  assign tensorFile_58_MPORT_122_data = tensorFile_58[tensorFile_58_MPORT_122_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_58_MPORT_58_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_58_MPORT_58_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_58_MPORT_58_mask = 1'h1;
  assign tensorFile_58_MPORT_58_en = _waddr_0_T ? 1'h0 : wenTensInstr_58;
  assign tensorFile_59_MPORT_123_en = tensorFile_59_MPORT_123_en_pipe_0;
  assign tensorFile_59_MPORT_123_addr = tensorFile_59_MPORT_123_addr_pipe_0;
  assign tensorFile_59_MPORT_123_data = tensorFile_59[tensorFile_59_MPORT_123_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_59_MPORT_59_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_59_MPORT_59_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_59_MPORT_59_mask = 1'h1;
  assign tensorFile_59_MPORT_59_en = _waddr_0_T ? 1'h0 : wenTensInstr_59;
  assign tensorFile_60_MPORT_124_en = tensorFile_60_MPORT_124_en_pipe_0;
  assign tensorFile_60_MPORT_124_addr = tensorFile_60_MPORT_124_addr_pipe_0;
  assign tensorFile_60_MPORT_124_data = tensorFile_60[tensorFile_60_MPORT_124_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_60_MPORT_60_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_60_MPORT_60_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_60_MPORT_60_mask = 1'h1;
  assign tensorFile_60_MPORT_60_en = _waddr_0_T ? 1'h0 : wenTensInstr_60;
  assign tensorFile_61_MPORT_125_en = tensorFile_61_MPORT_125_en_pipe_0;
  assign tensorFile_61_MPORT_125_addr = tensorFile_61_MPORT_125_addr_pipe_0;
  assign tensorFile_61_MPORT_125_data = tensorFile_61[tensorFile_61_MPORT_125_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_61_MPORT_61_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_61_MPORT_61_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_61_MPORT_61_mask = 1'h1;
  assign tensorFile_61_MPORT_61_en = _waddr_0_T ? 1'h0 : wenTensInstr_61;
  assign tensorFile_62_MPORT_126_en = tensorFile_62_MPORT_126_en_pipe_0;
  assign tensorFile_62_MPORT_126_addr = tensorFile_62_MPORT_126_addr_pipe_0;
  assign tensorFile_62_MPORT_126_data = tensorFile_62[tensorFile_62_MPORT_126_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_62_MPORT_62_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_62_MPORT_62_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_62_MPORT_62_mask = 1'h1;
  assign tensorFile_62_MPORT_62_en = _waddr_0_T ? 1'h0 : wenTensInstr_62;
  assign tensorFile_63_MPORT_127_en = tensorFile_63_MPORT_127_en_pipe_0;
  assign tensorFile_63_MPORT_127_addr = tensorFile_63_MPORT_127_addr_pipe_0;
  assign tensorFile_63_MPORT_127_data = tensorFile_63[tensorFile_63_MPORT_127_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_63_MPORT_63_data = _waddr_0_T ? 64'h0 : wdataTensInstr_0;
  assign tensorFile_63_MPORT_63_addr = _waddr_0_T ? 6'h0 : waddrTensInstrTmp;
  assign tensorFile_63_MPORT_63_mask = 1'h1;
  assign tensorFile_63_MPORT_63_en = _waddr_0_T ? 1'h0 : wenTensInstr_63;
  assign io_done = loadDone & fillPadding_io_done; // @[TensorLoadNarrowVME.scala 293:25]
  assign io_vme_rd_cmd_valid = vmeCmd_io_vmeCmd_valid; // @[TensorLoadNarrowVME.scala 80:20]
  assign io_vme_rd_cmd_bits_addr = vmeCmd_io_vmeCmd_bits_addr; // @[TensorLoadNarrowVME.scala 80:20]
  assign io_vme_rd_cmd_bits_len = vmeCmd_io_vmeCmd_bits_len; // @[TensorLoadNarrowVME.scala 80:20]
  assign io_vme_rd_cmd_bits_tag = vmeCmd_io_vmeCmd_bits_tag; // @[TensorLoadNarrowVME.scala 80:20]
  assign io_vme_rd_data_ready = 1'h1; // @[TensorLoadNarrowVME.scala 111:24]
  assign io_tensor_rd_0_data_valid = rvalid; // @[TensorLoadNarrowVME.scala 278:36]
  assign io_tensor_rd_0_data_bits_0_0 = _T_148[7:0]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_1 = _T_148[15:8]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_2 = _T_148[23:16]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_3 = _T_148[31:24]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_4 = _T_148[39:32]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_5 = _T_148[47:40]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_6 = _T_148[55:48]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_7 = _T_148[63:56]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_8 = _T_148[71:64]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_9 = _T_148[79:72]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_10 = _T_148[87:80]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_11 = _T_148[95:88]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_12 = _T_148[103:96]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_13 = _T_148[111:104]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_14 = _T_148[119:112]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_15 = _T_148[127:120]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_0 = _T_148[135:128]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_1 = _T_148[143:136]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_2 = _T_148[151:144]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_3 = _T_148[159:152]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_4 = _T_148[167:160]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_5 = _T_148[175:168]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_6 = _T_148[183:176]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_7 = _T_148[191:184]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_8 = _T_148[199:192]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_9 = _T_148[207:200]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_10 = _T_148[215:208]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_11 = _T_148[223:216]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_12 = _T_148[231:224]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_13 = _T_148[239:232]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_14 = _T_148[247:240]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_1_15 = _T_148[255:248]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_0 = _T_148[263:256]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_1 = _T_148[271:264]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_2 = _T_148[279:272]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_3 = _T_148[287:280]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_4 = _T_148[295:288]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_5 = _T_148[303:296]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_6 = _T_148[311:304]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_7 = _T_148[319:312]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_8 = _T_148[327:320]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_9 = _T_148[335:328]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_10 = _T_148[343:336]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_11 = _T_148[351:344]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_12 = _T_148[359:352]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_13 = _T_148[367:360]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_14 = _T_148[375:368]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_2_15 = _T_148[383:376]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_0 = _T_148[391:384]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_1 = _T_148[399:392]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_2 = _T_148[407:400]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_3 = _T_148[415:408]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_4 = _T_148[423:416]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_5 = _T_148[431:424]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_6 = _T_148[439:432]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_7 = _T_148[447:440]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_8 = _T_148[455:448]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_9 = _T_148[463:456]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_10 = _T_148[471:464]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_11 = _T_148[479:472]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_12 = _T_148[487:480]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_13 = _T_148[495:488]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_14 = _T_148[503:496]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_3_15 = _T_148[511:504]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_0 = _T_148[519:512]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_1 = _T_148[527:520]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_2 = _T_148[535:528]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_3 = _T_148[543:536]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_4 = _T_148[551:544]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_5 = _T_148[559:552]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_6 = _T_148[567:560]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_7 = _T_148[575:568]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_8 = _T_148[583:576]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_9 = _T_148[591:584]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_10 = _T_148[599:592]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_11 = _T_148[607:600]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_12 = _T_148[615:608]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_13 = _T_148[623:616]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_14 = _T_148[631:624]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_4_15 = _T_148[639:632]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_0 = _T_148[647:640]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_1 = _T_148[655:648]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_2 = _T_148[663:656]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_3 = _T_148[671:664]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_4 = _T_148[679:672]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_5 = _T_148[687:680]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_6 = _T_148[695:688]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_7 = _T_148[703:696]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_8 = _T_148[711:704]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_9 = _T_148[719:712]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_10 = _T_148[727:720]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_11 = _T_148[735:728]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_12 = _T_148[743:736]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_13 = _T_148[751:744]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_14 = _T_148[759:752]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_5_15 = _T_148[767:760]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_0 = _T_148[775:768]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_1 = _T_148[783:776]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_2 = _T_148[791:784]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_3 = _T_148[799:792]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_4 = _T_148[807:800]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_5 = _T_148[815:808]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_6 = _T_148[823:816]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_7 = _T_148[831:824]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_8 = _T_148[839:832]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_9 = _T_148[847:840]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_10 = _T_148[855:848]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_11 = _T_148[863:856]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_12 = _T_148[871:864]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_13 = _T_148[879:872]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_14 = _T_148[887:880]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_6_15 = _T_148[895:888]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_0 = _T_148[903:896]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_1 = _T_148[911:904]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_2 = _T_148[919:912]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_3 = _T_148[927:920]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_4 = _T_148[935:928]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_5 = _T_148[943:936]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_6 = _T_148[951:944]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_7 = _T_148[959:952]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_8 = _T_148[967:960]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_9 = _T_148[975:968]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_10 = _T_148[983:976]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_11 = _T_148[991:984]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_12 = _T_148[999:992]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_13 = _T_148[1007:1000]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_14 = _T_148[1015:1008]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_7_15 = _T_148[1023:1016]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_0 = _T_148[1031:1024]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_1 = _T_148[1039:1032]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_2 = _T_148[1047:1040]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_3 = _T_148[1055:1048]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_4 = _T_148[1063:1056]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_5 = _T_148[1071:1064]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_6 = _T_148[1079:1072]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_7 = _T_148[1087:1080]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_8 = _T_148[1095:1088]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_9 = _T_148[1103:1096]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_10 = _T_148[1111:1104]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_11 = _T_148[1119:1112]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_12 = _T_148[1127:1120]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_13 = _T_148[1135:1128]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_14 = _T_148[1143:1136]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_8_15 = _T_148[1151:1144]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_0 = _T_148[1159:1152]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_1 = _T_148[1167:1160]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_2 = _T_148[1175:1168]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_3 = _T_148[1183:1176]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_4 = _T_148[1191:1184]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_5 = _T_148[1199:1192]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_6 = _T_148[1207:1200]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_7 = _T_148[1215:1208]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_8 = _T_148[1223:1216]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_9 = _T_148[1231:1224]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_10 = _T_148[1239:1232]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_11 = _T_148[1247:1240]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_12 = _T_148[1255:1248]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_13 = _T_148[1263:1256]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_14 = _T_148[1271:1264]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_9_15 = _T_148[1279:1272]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_0 = _T_148[1287:1280]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_1 = _T_148[1295:1288]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_2 = _T_148[1303:1296]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_3 = _T_148[1311:1304]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_4 = _T_148[1319:1312]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_5 = _T_148[1327:1320]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_6 = _T_148[1335:1328]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_7 = _T_148[1343:1336]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_8 = _T_148[1351:1344]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_9 = _T_148[1359:1352]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_10 = _T_148[1367:1360]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_11 = _T_148[1375:1368]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_12 = _T_148[1383:1376]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_13 = _T_148[1391:1384]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_14 = _T_148[1399:1392]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_10_15 = _T_148[1407:1400]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_0 = _T_148[1415:1408]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_1 = _T_148[1423:1416]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_2 = _T_148[1431:1424]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_3 = _T_148[1439:1432]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_4 = _T_148[1447:1440]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_5 = _T_148[1455:1448]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_6 = _T_148[1463:1456]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_7 = _T_148[1471:1464]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_8 = _T_148[1479:1472]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_9 = _T_148[1487:1480]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_10 = _T_148[1495:1488]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_11 = _T_148[1503:1496]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_12 = _T_148[1511:1504]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_13 = _T_148[1519:1512]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_14 = _T_148[1527:1520]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_11_15 = _T_148[1535:1528]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_0 = _T_148[1543:1536]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_1 = _T_148[1551:1544]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_2 = _T_148[1559:1552]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_3 = _T_148[1567:1560]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_4 = _T_148[1575:1568]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_5 = _T_148[1583:1576]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_6 = _T_148[1591:1584]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_7 = _T_148[1599:1592]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_8 = _T_148[1607:1600]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_9 = _T_148[1615:1608]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_10 = _T_148[1623:1616]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_11 = _T_148[1631:1624]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_12 = _T_148[1639:1632]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_13 = _T_148[1647:1640]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_14 = _T_148[1655:1648]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_12_15 = _T_148[1663:1656]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_0 = _T_148[1671:1664]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_1 = _T_148[1679:1672]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_2 = _T_148[1687:1680]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_3 = _T_148[1695:1688]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_4 = _T_148[1703:1696]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_5 = _T_148[1711:1704]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_6 = _T_148[1719:1712]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_7 = _T_148[1727:1720]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_8 = _T_148[1735:1728]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_9 = _T_148[1743:1736]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_10 = _T_148[1751:1744]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_11 = _T_148[1759:1752]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_12 = _T_148[1767:1760]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_13 = _T_148[1775:1768]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_14 = _T_148[1783:1776]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_13_15 = _T_148[1791:1784]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_0 = _T_148[1799:1792]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_1 = _T_148[1807:1800]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_2 = _T_148[1815:1808]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_3 = _T_148[1823:1816]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_4 = _T_148[1831:1824]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_5 = _T_148[1839:1832]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_6 = _T_148[1847:1840]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_7 = _T_148[1855:1848]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_8 = _T_148[1863:1856]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_9 = _T_148[1871:1864]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_10 = _T_148[1879:1872]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_11 = _T_148[1887:1880]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_12 = _T_148[1895:1888]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_13 = _T_148[1903:1896]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_14 = _T_148[1911:1904]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_14_15 = _T_148[1919:1912]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_0 = _T_148[1927:1920]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_1 = _T_148[1935:1928]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_2 = _T_148[1943:1936]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_3 = _T_148[1951:1944]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_4 = _T_148[1959:1952]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_5 = _T_148[1967:1960]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_6 = _T_148[1975:1968]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_7 = _T_148[1983:1976]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_8 = _T_148[1991:1984]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_9 = _T_148[1999:1992]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_10 = _T_148[2007:2000]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_11 = _T_148[2015:2008]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_12 = _T_148[2023:2016]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_13 = _T_148[2031:2024]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_14 = _T_148[2039:2032]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_15_15 = _T_148[2047:2040]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_16_0 = _T_148[2055:2048]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_16_1 = _T_148[2063:2056]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_16_2 = _T_148[2071:2064]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_16_3 = _T_148[2079:2072]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_16_4 = _T_148[2087:2080]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_16_5 = _T_148[2095:2088]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_16_6 = _T_148[2103:2096]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_16_7 = _T_148[2111:2104]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_16_8 = _T_148[2119:2112]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_16_9 = _T_148[2127:2120]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_16_10 = _T_148[2135:2128]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_16_11 = _T_148[2143:2136]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_16_12 = _T_148[2151:2144]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_16_13 = _T_148[2159:2152]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_16_14 = _T_148[2167:2160]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_16_15 = _T_148[2175:2168]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_17_0 = _T_148[2183:2176]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_17_1 = _T_148[2191:2184]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_17_2 = _T_148[2199:2192]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_17_3 = _T_148[2207:2200]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_17_4 = _T_148[2215:2208]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_17_5 = _T_148[2223:2216]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_17_6 = _T_148[2231:2224]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_17_7 = _T_148[2239:2232]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_17_8 = _T_148[2247:2240]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_17_9 = _T_148[2255:2248]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_17_10 = _T_148[2263:2256]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_17_11 = _T_148[2271:2264]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_17_12 = _T_148[2279:2272]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_17_13 = _T_148[2287:2280]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_17_14 = _T_148[2295:2288]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_17_15 = _T_148[2303:2296]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_18_0 = _T_148[2311:2304]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_18_1 = _T_148[2319:2312]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_18_2 = _T_148[2327:2320]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_18_3 = _T_148[2335:2328]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_18_4 = _T_148[2343:2336]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_18_5 = _T_148[2351:2344]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_18_6 = _T_148[2359:2352]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_18_7 = _T_148[2367:2360]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_18_8 = _T_148[2375:2368]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_18_9 = _T_148[2383:2376]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_18_10 = _T_148[2391:2384]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_18_11 = _T_148[2399:2392]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_18_12 = _T_148[2407:2400]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_18_13 = _T_148[2415:2408]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_18_14 = _T_148[2423:2416]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_18_15 = _T_148[2431:2424]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_19_0 = _T_148[2439:2432]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_19_1 = _T_148[2447:2440]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_19_2 = _T_148[2455:2448]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_19_3 = _T_148[2463:2456]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_19_4 = _T_148[2471:2464]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_19_5 = _T_148[2479:2472]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_19_6 = _T_148[2487:2480]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_19_7 = _T_148[2495:2488]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_19_8 = _T_148[2503:2496]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_19_9 = _T_148[2511:2504]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_19_10 = _T_148[2519:2512]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_19_11 = _T_148[2527:2520]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_19_12 = _T_148[2535:2528]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_19_13 = _T_148[2543:2536]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_19_14 = _T_148[2551:2544]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_19_15 = _T_148[2559:2552]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_20_0 = _T_148[2567:2560]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_20_1 = _T_148[2575:2568]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_20_2 = _T_148[2583:2576]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_20_3 = _T_148[2591:2584]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_20_4 = _T_148[2599:2592]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_20_5 = _T_148[2607:2600]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_20_6 = _T_148[2615:2608]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_20_7 = _T_148[2623:2616]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_20_8 = _T_148[2631:2624]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_20_9 = _T_148[2639:2632]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_20_10 = _T_148[2647:2640]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_20_11 = _T_148[2655:2648]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_20_12 = _T_148[2663:2656]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_20_13 = _T_148[2671:2664]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_20_14 = _T_148[2679:2672]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_20_15 = _T_148[2687:2680]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_21_0 = _T_148[2695:2688]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_21_1 = _T_148[2703:2696]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_21_2 = _T_148[2711:2704]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_21_3 = _T_148[2719:2712]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_21_4 = _T_148[2727:2720]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_21_5 = _T_148[2735:2728]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_21_6 = _T_148[2743:2736]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_21_7 = _T_148[2751:2744]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_21_8 = _T_148[2759:2752]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_21_9 = _T_148[2767:2760]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_21_10 = _T_148[2775:2768]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_21_11 = _T_148[2783:2776]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_21_12 = _T_148[2791:2784]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_21_13 = _T_148[2799:2792]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_21_14 = _T_148[2807:2800]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_21_15 = _T_148[2815:2808]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_22_0 = _T_148[2823:2816]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_22_1 = _T_148[2831:2824]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_22_2 = _T_148[2839:2832]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_22_3 = _T_148[2847:2840]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_22_4 = _T_148[2855:2848]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_22_5 = _T_148[2863:2856]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_22_6 = _T_148[2871:2864]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_22_7 = _T_148[2879:2872]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_22_8 = _T_148[2887:2880]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_22_9 = _T_148[2895:2888]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_22_10 = _T_148[2903:2896]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_22_11 = _T_148[2911:2904]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_22_12 = _T_148[2919:2912]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_22_13 = _T_148[2927:2920]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_22_14 = _T_148[2935:2928]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_22_15 = _T_148[2943:2936]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_23_0 = _T_148[2951:2944]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_23_1 = _T_148[2959:2952]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_23_2 = _T_148[2967:2960]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_23_3 = _T_148[2975:2968]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_23_4 = _T_148[2983:2976]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_23_5 = _T_148[2991:2984]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_23_6 = _T_148[2999:2992]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_23_7 = _T_148[3007:3000]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_23_8 = _T_148[3015:3008]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_23_9 = _T_148[3023:3016]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_23_10 = _T_148[3031:3024]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_23_11 = _T_148[3039:3032]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_23_12 = _T_148[3047:3040]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_23_13 = _T_148[3055:3048]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_23_14 = _T_148[3063:3056]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_23_15 = _T_148[3071:3064]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_24_0 = _T_148[3079:3072]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_24_1 = _T_148[3087:3080]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_24_2 = _T_148[3095:3088]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_24_3 = _T_148[3103:3096]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_24_4 = _T_148[3111:3104]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_24_5 = _T_148[3119:3112]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_24_6 = _T_148[3127:3120]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_24_7 = _T_148[3135:3128]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_24_8 = _T_148[3143:3136]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_24_9 = _T_148[3151:3144]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_24_10 = _T_148[3159:3152]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_24_11 = _T_148[3167:3160]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_24_12 = _T_148[3175:3168]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_24_13 = _T_148[3183:3176]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_24_14 = _T_148[3191:3184]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_24_15 = _T_148[3199:3192]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_25_0 = _T_148[3207:3200]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_25_1 = _T_148[3215:3208]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_25_2 = _T_148[3223:3216]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_25_3 = _T_148[3231:3224]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_25_4 = _T_148[3239:3232]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_25_5 = _T_148[3247:3240]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_25_6 = _T_148[3255:3248]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_25_7 = _T_148[3263:3256]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_25_8 = _T_148[3271:3264]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_25_9 = _T_148[3279:3272]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_25_10 = _T_148[3287:3280]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_25_11 = _T_148[3295:3288]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_25_12 = _T_148[3303:3296]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_25_13 = _T_148[3311:3304]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_25_14 = _T_148[3319:3312]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_25_15 = _T_148[3327:3320]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_26_0 = _T_148[3335:3328]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_26_1 = _T_148[3343:3336]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_26_2 = _T_148[3351:3344]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_26_3 = _T_148[3359:3352]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_26_4 = _T_148[3367:3360]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_26_5 = _T_148[3375:3368]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_26_6 = _T_148[3383:3376]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_26_7 = _T_148[3391:3384]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_26_8 = _T_148[3399:3392]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_26_9 = _T_148[3407:3400]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_26_10 = _T_148[3415:3408]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_26_11 = _T_148[3423:3416]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_26_12 = _T_148[3431:3424]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_26_13 = _T_148[3439:3432]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_26_14 = _T_148[3447:3440]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_26_15 = _T_148[3455:3448]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_27_0 = _T_148[3463:3456]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_27_1 = _T_148[3471:3464]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_27_2 = _T_148[3479:3472]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_27_3 = _T_148[3487:3480]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_27_4 = _T_148[3495:3488]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_27_5 = _T_148[3503:3496]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_27_6 = _T_148[3511:3504]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_27_7 = _T_148[3519:3512]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_27_8 = _T_148[3527:3520]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_27_9 = _T_148[3535:3528]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_27_10 = _T_148[3543:3536]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_27_11 = _T_148[3551:3544]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_27_12 = _T_148[3559:3552]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_27_13 = _T_148[3567:3560]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_27_14 = _T_148[3575:3568]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_27_15 = _T_148[3583:3576]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_28_0 = _T_148[3591:3584]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_28_1 = _T_148[3599:3592]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_28_2 = _T_148[3607:3600]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_28_3 = _T_148[3615:3608]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_28_4 = _T_148[3623:3616]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_28_5 = _T_148[3631:3624]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_28_6 = _T_148[3639:3632]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_28_7 = _T_148[3647:3640]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_28_8 = _T_148[3655:3648]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_28_9 = _T_148[3663:3656]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_28_10 = _T_148[3671:3664]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_28_11 = _T_148[3679:3672]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_28_12 = _T_148[3687:3680]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_28_13 = _T_148[3695:3688]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_28_14 = _T_148[3703:3696]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_28_15 = _T_148[3711:3704]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_29_0 = _T_148[3719:3712]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_29_1 = _T_148[3727:3720]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_29_2 = _T_148[3735:3728]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_29_3 = _T_148[3743:3736]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_29_4 = _T_148[3751:3744]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_29_5 = _T_148[3759:3752]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_29_6 = _T_148[3767:3760]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_29_7 = _T_148[3775:3768]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_29_8 = _T_148[3783:3776]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_29_9 = _T_148[3791:3784]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_29_10 = _T_148[3799:3792]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_29_11 = _T_148[3807:3800]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_29_12 = _T_148[3815:3808]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_29_13 = _T_148[3823:3816]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_29_14 = _T_148[3831:3824]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_29_15 = _T_148[3839:3832]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_30_0 = _T_148[3847:3840]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_30_1 = _T_148[3855:3848]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_30_2 = _T_148[3863:3856]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_30_3 = _T_148[3871:3864]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_30_4 = _T_148[3879:3872]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_30_5 = _T_148[3887:3880]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_30_6 = _T_148[3895:3888]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_30_7 = _T_148[3903:3896]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_30_8 = _T_148[3911:3904]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_30_9 = _T_148[3919:3912]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_30_10 = _T_148[3927:3920]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_30_11 = _T_148[3935:3928]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_30_12 = _T_148[3943:3936]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_30_13 = _T_148[3951:3944]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_30_14 = _T_148[3959:3952]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_30_15 = _T_148[3967:3960]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_31_0 = _T_148[3975:3968]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_31_1 = _T_148[3983:3976]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_31_2 = _T_148[3991:3984]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_31_3 = _T_148[3999:3992]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_31_4 = _T_148[4007:4000]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_31_5 = _T_148[4015:4008]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_31_6 = _T_148[4023:4016]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_31_7 = _T_148[4031:4024]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_31_8 = _T_148[4039:4032]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_31_9 = _T_148[4047:4040]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_31_10 = _T_148[4055:4048]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_31_11 = _T_148[4063:4056]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_31_12 = _T_148[4071:4064]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_31_13 = _T_148[4079:4072]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_31_14 = _T_148[4087:4080]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_31_15 = _T_148[4095:4088]; // @[TensorLoadNarrowVME.scala 288:18]
  assign vmeCmd_clock = clock;
  assign vmeCmd_reset = reset;
  assign vmeCmd_io_start = io_start; // @[TensorLoadNarrowVME.scala 76:19]
  assign vmeCmd_io_isBusy = state; // @[TensorLoadNarrowVME.scala 56:22]
  assign vmeCmd_io_inst = io_inst; // @[TensorLoadNarrowVME.scala 78:18]
  assign vmeCmd_io_baddr = io_baddr; // @[TensorLoadNarrowVME.scala 79:19]
  assign vmeCmd_io_vmeCmd_ready = io_vme_rd_cmd_ready; // @[TensorLoadNarrowVME.scala 80:20]
  assign readData_clock = clock;
  assign readData_reset = reset;
  assign readData_io_start = io_start; // @[TensorLoadNarrowVME.scala 106:21]
  assign readData_io_vmeData_valid = vmeDataValidPipe; // @[TensorLoadNarrowVME.scala 107:29]
  assign readData_io_vmeData_bits_tag = vmeDataBitsPipe_tag; // @[TensorLoadNarrowVME.scala 108:28]
  assign fillPadding_clock = clock;
  assign fillPadding_reset = reset;
  assign fillPadding_io_canWriteMem = ~vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 120:33]
  assign fillPadding_io_inst = fillPadding_io_inst_REG; // @[TensorLoadNarrowVME.scala 121:23]
  assign fillPadding_io_start = fillPadding_io_start_REG; // @[TensorLoadNarrowVME.scala 122:24]
  always @(posedge clock) begin
    if (tensorFile_0_MPORT_en & tensorFile_0_MPORT_mask) begin
      tensorFile_0[tensorFile_0_MPORT_addr] <= tensorFile_0_MPORT_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_0_MPORT_64_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_0_MPORT_64_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_1_MPORT_1_en & tensorFile_1_MPORT_1_mask) begin
      tensorFile_1[tensorFile_1_MPORT_1_addr] <= tensorFile_1_MPORT_1_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_1_MPORT_65_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_1_MPORT_65_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_2_MPORT_2_en & tensorFile_2_MPORT_2_mask) begin
      tensorFile_2[tensorFile_2_MPORT_2_addr] <= tensorFile_2_MPORT_2_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_2_MPORT_66_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_2_MPORT_66_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_3_MPORT_3_en & tensorFile_3_MPORT_3_mask) begin
      tensorFile_3[tensorFile_3_MPORT_3_addr] <= tensorFile_3_MPORT_3_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_3_MPORT_67_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_3_MPORT_67_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_4_MPORT_4_en & tensorFile_4_MPORT_4_mask) begin
      tensorFile_4[tensorFile_4_MPORT_4_addr] <= tensorFile_4_MPORT_4_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_4_MPORT_68_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_4_MPORT_68_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_5_MPORT_5_en & tensorFile_5_MPORT_5_mask) begin
      tensorFile_5[tensorFile_5_MPORT_5_addr] <= tensorFile_5_MPORT_5_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_5_MPORT_69_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_5_MPORT_69_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_6_MPORT_6_en & tensorFile_6_MPORT_6_mask) begin
      tensorFile_6[tensorFile_6_MPORT_6_addr] <= tensorFile_6_MPORT_6_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_6_MPORT_70_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_6_MPORT_70_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_7_MPORT_7_en & tensorFile_7_MPORT_7_mask) begin
      tensorFile_7[tensorFile_7_MPORT_7_addr] <= tensorFile_7_MPORT_7_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_7_MPORT_71_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_7_MPORT_71_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_8_MPORT_8_en & tensorFile_8_MPORT_8_mask) begin
      tensorFile_8[tensorFile_8_MPORT_8_addr] <= tensorFile_8_MPORT_8_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_8_MPORT_72_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_8_MPORT_72_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_9_MPORT_9_en & tensorFile_9_MPORT_9_mask) begin
      tensorFile_9[tensorFile_9_MPORT_9_addr] <= tensorFile_9_MPORT_9_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_9_MPORT_73_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_9_MPORT_73_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_10_MPORT_10_en & tensorFile_10_MPORT_10_mask) begin
      tensorFile_10[tensorFile_10_MPORT_10_addr] <= tensorFile_10_MPORT_10_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_10_MPORT_74_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_10_MPORT_74_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_11_MPORT_11_en & tensorFile_11_MPORT_11_mask) begin
      tensorFile_11[tensorFile_11_MPORT_11_addr] <= tensorFile_11_MPORT_11_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_11_MPORT_75_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_11_MPORT_75_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_12_MPORT_12_en & tensorFile_12_MPORT_12_mask) begin
      tensorFile_12[tensorFile_12_MPORT_12_addr] <= tensorFile_12_MPORT_12_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_12_MPORT_76_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_12_MPORT_76_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_13_MPORT_13_en & tensorFile_13_MPORT_13_mask) begin
      tensorFile_13[tensorFile_13_MPORT_13_addr] <= tensorFile_13_MPORT_13_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_13_MPORT_77_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_13_MPORT_77_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_14_MPORT_14_en & tensorFile_14_MPORT_14_mask) begin
      tensorFile_14[tensorFile_14_MPORT_14_addr] <= tensorFile_14_MPORT_14_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_14_MPORT_78_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_14_MPORT_78_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_15_MPORT_15_en & tensorFile_15_MPORT_15_mask) begin
      tensorFile_15[tensorFile_15_MPORT_15_addr] <= tensorFile_15_MPORT_15_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_15_MPORT_79_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_15_MPORT_79_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_16_MPORT_16_en & tensorFile_16_MPORT_16_mask) begin
      tensorFile_16[tensorFile_16_MPORT_16_addr] <= tensorFile_16_MPORT_16_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_16_MPORT_80_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_16_MPORT_80_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_17_MPORT_17_en & tensorFile_17_MPORT_17_mask) begin
      tensorFile_17[tensorFile_17_MPORT_17_addr] <= tensorFile_17_MPORT_17_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_17_MPORT_81_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_17_MPORT_81_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_18_MPORT_18_en & tensorFile_18_MPORT_18_mask) begin
      tensorFile_18[tensorFile_18_MPORT_18_addr] <= tensorFile_18_MPORT_18_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_18_MPORT_82_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_18_MPORT_82_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_19_MPORT_19_en & tensorFile_19_MPORT_19_mask) begin
      tensorFile_19[tensorFile_19_MPORT_19_addr] <= tensorFile_19_MPORT_19_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_19_MPORT_83_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_19_MPORT_83_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_20_MPORT_20_en & tensorFile_20_MPORT_20_mask) begin
      tensorFile_20[tensorFile_20_MPORT_20_addr] <= tensorFile_20_MPORT_20_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_20_MPORT_84_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_20_MPORT_84_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_21_MPORT_21_en & tensorFile_21_MPORT_21_mask) begin
      tensorFile_21[tensorFile_21_MPORT_21_addr] <= tensorFile_21_MPORT_21_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_21_MPORT_85_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_21_MPORT_85_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_22_MPORT_22_en & tensorFile_22_MPORT_22_mask) begin
      tensorFile_22[tensorFile_22_MPORT_22_addr] <= tensorFile_22_MPORT_22_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_22_MPORT_86_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_22_MPORT_86_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_23_MPORT_23_en & tensorFile_23_MPORT_23_mask) begin
      tensorFile_23[tensorFile_23_MPORT_23_addr] <= tensorFile_23_MPORT_23_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_23_MPORT_87_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_23_MPORT_87_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_24_MPORT_24_en & tensorFile_24_MPORT_24_mask) begin
      tensorFile_24[tensorFile_24_MPORT_24_addr] <= tensorFile_24_MPORT_24_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_24_MPORT_88_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_24_MPORT_88_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_25_MPORT_25_en & tensorFile_25_MPORT_25_mask) begin
      tensorFile_25[tensorFile_25_MPORT_25_addr] <= tensorFile_25_MPORT_25_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_25_MPORT_89_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_25_MPORT_89_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_26_MPORT_26_en & tensorFile_26_MPORT_26_mask) begin
      tensorFile_26[tensorFile_26_MPORT_26_addr] <= tensorFile_26_MPORT_26_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_26_MPORT_90_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_26_MPORT_90_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_27_MPORT_27_en & tensorFile_27_MPORT_27_mask) begin
      tensorFile_27[tensorFile_27_MPORT_27_addr] <= tensorFile_27_MPORT_27_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_27_MPORT_91_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_27_MPORT_91_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_28_MPORT_28_en & tensorFile_28_MPORT_28_mask) begin
      tensorFile_28[tensorFile_28_MPORT_28_addr] <= tensorFile_28_MPORT_28_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_28_MPORT_92_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_28_MPORT_92_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_29_MPORT_29_en & tensorFile_29_MPORT_29_mask) begin
      tensorFile_29[tensorFile_29_MPORT_29_addr] <= tensorFile_29_MPORT_29_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_29_MPORT_93_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_29_MPORT_93_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_30_MPORT_30_en & tensorFile_30_MPORT_30_mask) begin
      tensorFile_30[tensorFile_30_MPORT_30_addr] <= tensorFile_30_MPORT_30_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_30_MPORT_94_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_30_MPORT_94_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_31_MPORT_31_en & tensorFile_31_MPORT_31_mask) begin
      tensorFile_31[tensorFile_31_MPORT_31_addr] <= tensorFile_31_MPORT_31_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_31_MPORT_95_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_31_MPORT_95_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_32_MPORT_32_en & tensorFile_32_MPORT_32_mask) begin
      tensorFile_32[tensorFile_32_MPORT_32_addr] <= tensorFile_32_MPORT_32_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_32_MPORT_96_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_32_MPORT_96_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_33_MPORT_33_en & tensorFile_33_MPORT_33_mask) begin
      tensorFile_33[tensorFile_33_MPORT_33_addr] <= tensorFile_33_MPORT_33_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_33_MPORT_97_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_33_MPORT_97_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_34_MPORT_34_en & tensorFile_34_MPORT_34_mask) begin
      tensorFile_34[tensorFile_34_MPORT_34_addr] <= tensorFile_34_MPORT_34_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_34_MPORT_98_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_34_MPORT_98_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_35_MPORT_35_en & tensorFile_35_MPORT_35_mask) begin
      tensorFile_35[tensorFile_35_MPORT_35_addr] <= tensorFile_35_MPORT_35_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_35_MPORT_99_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_35_MPORT_99_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_36_MPORT_36_en & tensorFile_36_MPORT_36_mask) begin
      tensorFile_36[tensorFile_36_MPORT_36_addr] <= tensorFile_36_MPORT_36_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_36_MPORT_100_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_36_MPORT_100_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_37_MPORT_37_en & tensorFile_37_MPORT_37_mask) begin
      tensorFile_37[tensorFile_37_MPORT_37_addr] <= tensorFile_37_MPORT_37_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_37_MPORT_101_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_37_MPORT_101_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_38_MPORT_38_en & tensorFile_38_MPORT_38_mask) begin
      tensorFile_38[tensorFile_38_MPORT_38_addr] <= tensorFile_38_MPORT_38_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_38_MPORT_102_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_38_MPORT_102_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_39_MPORT_39_en & tensorFile_39_MPORT_39_mask) begin
      tensorFile_39[tensorFile_39_MPORT_39_addr] <= tensorFile_39_MPORT_39_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_39_MPORT_103_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_39_MPORT_103_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_40_MPORT_40_en & tensorFile_40_MPORT_40_mask) begin
      tensorFile_40[tensorFile_40_MPORT_40_addr] <= tensorFile_40_MPORT_40_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_40_MPORT_104_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_40_MPORT_104_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_41_MPORT_41_en & tensorFile_41_MPORT_41_mask) begin
      tensorFile_41[tensorFile_41_MPORT_41_addr] <= tensorFile_41_MPORT_41_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_41_MPORT_105_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_41_MPORT_105_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_42_MPORT_42_en & tensorFile_42_MPORT_42_mask) begin
      tensorFile_42[tensorFile_42_MPORT_42_addr] <= tensorFile_42_MPORT_42_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_42_MPORT_106_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_42_MPORT_106_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_43_MPORT_43_en & tensorFile_43_MPORT_43_mask) begin
      tensorFile_43[tensorFile_43_MPORT_43_addr] <= tensorFile_43_MPORT_43_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_43_MPORT_107_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_43_MPORT_107_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_44_MPORT_44_en & tensorFile_44_MPORT_44_mask) begin
      tensorFile_44[tensorFile_44_MPORT_44_addr] <= tensorFile_44_MPORT_44_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_44_MPORT_108_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_44_MPORT_108_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_45_MPORT_45_en & tensorFile_45_MPORT_45_mask) begin
      tensorFile_45[tensorFile_45_MPORT_45_addr] <= tensorFile_45_MPORT_45_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_45_MPORT_109_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_45_MPORT_109_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_46_MPORT_46_en & tensorFile_46_MPORT_46_mask) begin
      tensorFile_46[tensorFile_46_MPORT_46_addr] <= tensorFile_46_MPORT_46_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_46_MPORT_110_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_46_MPORT_110_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_47_MPORT_47_en & tensorFile_47_MPORT_47_mask) begin
      tensorFile_47[tensorFile_47_MPORT_47_addr] <= tensorFile_47_MPORT_47_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_47_MPORT_111_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_47_MPORT_111_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_48_MPORT_48_en & tensorFile_48_MPORT_48_mask) begin
      tensorFile_48[tensorFile_48_MPORT_48_addr] <= tensorFile_48_MPORT_48_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_48_MPORT_112_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_48_MPORT_112_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_49_MPORT_49_en & tensorFile_49_MPORT_49_mask) begin
      tensorFile_49[tensorFile_49_MPORT_49_addr] <= tensorFile_49_MPORT_49_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_49_MPORT_113_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_49_MPORT_113_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_50_MPORT_50_en & tensorFile_50_MPORT_50_mask) begin
      tensorFile_50[tensorFile_50_MPORT_50_addr] <= tensorFile_50_MPORT_50_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_50_MPORT_114_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_50_MPORT_114_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_51_MPORT_51_en & tensorFile_51_MPORT_51_mask) begin
      tensorFile_51[tensorFile_51_MPORT_51_addr] <= tensorFile_51_MPORT_51_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_51_MPORT_115_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_51_MPORT_115_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_52_MPORT_52_en & tensorFile_52_MPORT_52_mask) begin
      tensorFile_52[tensorFile_52_MPORT_52_addr] <= tensorFile_52_MPORT_52_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_52_MPORT_116_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_52_MPORT_116_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_53_MPORT_53_en & tensorFile_53_MPORT_53_mask) begin
      tensorFile_53[tensorFile_53_MPORT_53_addr] <= tensorFile_53_MPORT_53_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_53_MPORT_117_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_53_MPORT_117_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_54_MPORT_54_en & tensorFile_54_MPORT_54_mask) begin
      tensorFile_54[tensorFile_54_MPORT_54_addr] <= tensorFile_54_MPORT_54_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_54_MPORT_118_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_54_MPORT_118_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_55_MPORT_55_en & tensorFile_55_MPORT_55_mask) begin
      tensorFile_55[tensorFile_55_MPORT_55_addr] <= tensorFile_55_MPORT_55_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_55_MPORT_119_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_55_MPORT_119_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_56_MPORT_56_en & tensorFile_56_MPORT_56_mask) begin
      tensorFile_56[tensorFile_56_MPORT_56_addr] <= tensorFile_56_MPORT_56_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_56_MPORT_120_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_56_MPORT_120_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_57_MPORT_57_en & tensorFile_57_MPORT_57_mask) begin
      tensorFile_57[tensorFile_57_MPORT_57_addr] <= tensorFile_57_MPORT_57_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_57_MPORT_121_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_57_MPORT_121_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_58_MPORT_58_en & tensorFile_58_MPORT_58_mask) begin
      tensorFile_58[tensorFile_58_MPORT_58_addr] <= tensorFile_58_MPORT_58_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_58_MPORT_122_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_58_MPORT_122_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_59_MPORT_59_en & tensorFile_59_MPORT_59_mask) begin
      tensorFile_59[tensorFile_59_MPORT_59_addr] <= tensorFile_59_MPORT_59_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_59_MPORT_123_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_59_MPORT_123_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_60_MPORT_60_en & tensorFile_60_MPORT_60_mask) begin
      tensorFile_60[tensorFile_60_MPORT_60_addr] <= tensorFile_60_MPORT_60_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_60_MPORT_124_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_60_MPORT_124_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_61_MPORT_61_en & tensorFile_61_MPORT_61_mask) begin
      tensorFile_61[tensorFile_61_MPORT_61_addr] <= tensorFile_61_MPORT_61_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_61_MPORT_125_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_61_MPORT_125_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_62_MPORT_62_en & tensorFile_62_MPORT_62_mask) begin
      tensorFile_62[tensorFile_62_MPORT_62_addr] <= tensorFile_62_MPORT_62_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_62_MPORT_126_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_62_MPORT_126_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_63_MPORT_63_en & tensorFile_63_MPORT_63_mask) begin
      tensorFile_63[tensorFile_63_MPORT_63_addr] <= tensorFile_63_MPORT_63_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_63_MPORT_127_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_63_MPORT_127_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (reset) begin // @[TensorLoadNarrowVME.scala 54:22]
      state <= 1'h0; // @[TensorLoadNarrowVME.scala 54:22]
    end else begin
      state <= _GEN_1;
    end
    if (io_start) begin // @[TensorLoadNarrowVME.scala 88:18]
      blocksInFlight <= 12'h0; // @[TensorLoadNarrowVME.scala 89:20]
    end else if (state & _T & ~vmeDataFirePipe) begin // @[TensorLoadNarrowVME.scala 90:64]
      blocksInFlight <= _blocksInFlight_T_1; // @[TensorLoadNarrowVME.scala 91:20]
    end else if (_T_1 & vmeDataFirePipe) begin // @[TensorLoadNarrowVME.scala 92:63]
      blocksInFlight <= _blocksInFlight_T_5; // @[TensorLoadNarrowVME.scala 93:20]
    end else if (state & ~_T & vmeDataFirePipe) begin // @[TensorLoadNarrowVME.scala 94:64]
      blocksInFlight <= _blocksInFlight_T_7; // @[TensorLoadNarrowVME.scala 96:20]
    end
    vmeDataBitsPipe_data <= io_vme_rd_data_bits_data; // @[TensorLoadNarrowVME.scala 67:32]
    vmeDataBitsPipe_tag <= io_vme_rd_data_bits_tag; // @[TensorLoadNarrowVME.scala 67:32]
    if (reset) begin // @[TensorLoadNarrowVME.scala 68:33]
      vmeDataValidPipe <= 1'h0; // @[TensorLoadNarrowVME.scala 68:33]
    end else begin
      vmeDataValidPipe <= io_vme_rd_data_valid; // @[TensorLoadNarrowVME.scala 68:33]
    end
    if (reset) begin // @[TensorLoadNarrowVME.scala 69:33]
      vmeDataReadyPipe <= 1'h0; // @[TensorLoadNarrowVME.scala 69:33]
    end else begin
      vmeDataReadyPipe <= io_vme_rd_data_ready; // @[TensorLoadNarrowVME.scala 69:33]
    end
    fillPadding_io_inst_REG <= io_inst; // @[TensorLoadNarrowVME.scala 121:33]
    if (reset) begin // @[TensorLoadNarrowVME.scala 122:34]
      fillPadding_io_start_REG <= 1'h0; // @[TensorLoadNarrowVME.scala 122:34]
    end else begin
      fillPadding_io_start_REG <= io_start; // @[TensorLoadNarrowVME.scala 122:34]
    end
    if (reset) begin // @[Reg.scala 28:20]
      rvalid <= 1'h0; // @[Reg.scala 28:20]
    end else begin
      rvalid <= io_tensor_rd_0_idx_valid;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~io_start & ~_T_3 & ~_T_6 & _T_10 & ~reset & ~(blocksInFlight > 12'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TensorLoadNarrowVME.scala:95 assert(blocksInFlight > 0.U)\n"); // @[TensorLoadNarrowVME.scala 95:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_0[initvar] = _RAND_0[63:0];
  _RAND_3 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_1[initvar] = _RAND_3[63:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_2[initvar] = _RAND_6[63:0];
  _RAND_9 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_3[initvar] = _RAND_9[63:0];
  _RAND_12 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_4[initvar] = _RAND_12[63:0];
  _RAND_15 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_5[initvar] = _RAND_15[63:0];
  _RAND_18 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_6[initvar] = _RAND_18[63:0];
  _RAND_21 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_7[initvar] = _RAND_21[63:0];
  _RAND_24 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_8[initvar] = _RAND_24[63:0];
  _RAND_27 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_9[initvar] = _RAND_27[63:0];
  _RAND_30 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_10[initvar] = _RAND_30[63:0];
  _RAND_33 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_11[initvar] = _RAND_33[63:0];
  _RAND_36 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_12[initvar] = _RAND_36[63:0];
  _RAND_39 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_13[initvar] = _RAND_39[63:0];
  _RAND_42 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_14[initvar] = _RAND_42[63:0];
  _RAND_45 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_15[initvar] = _RAND_45[63:0];
  _RAND_48 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_16[initvar] = _RAND_48[63:0];
  _RAND_51 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_17[initvar] = _RAND_51[63:0];
  _RAND_54 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_18[initvar] = _RAND_54[63:0];
  _RAND_57 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_19[initvar] = _RAND_57[63:0];
  _RAND_60 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_20[initvar] = _RAND_60[63:0];
  _RAND_63 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_21[initvar] = _RAND_63[63:0];
  _RAND_66 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_22[initvar] = _RAND_66[63:0];
  _RAND_69 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_23[initvar] = _RAND_69[63:0];
  _RAND_72 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_24[initvar] = _RAND_72[63:0];
  _RAND_75 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_25[initvar] = _RAND_75[63:0];
  _RAND_78 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_26[initvar] = _RAND_78[63:0];
  _RAND_81 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_27[initvar] = _RAND_81[63:0];
  _RAND_84 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_28[initvar] = _RAND_84[63:0];
  _RAND_87 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_29[initvar] = _RAND_87[63:0];
  _RAND_90 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_30[initvar] = _RAND_90[63:0];
  _RAND_93 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_31[initvar] = _RAND_93[63:0];
  _RAND_96 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_32[initvar] = _RAND_96[63:0];
  _RAND_99 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_33[initvar] = _RAND_99[63:0];
  _RAND_102 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_34[initvar] = _RAND_102[63:0];
  _RAND_105 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_35[initvar] = _RAND_105[63:0];
  _RAND_108 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_36[initvar] = _RAND_108[63:0];
  _RAND_111 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_37[initvar] = _RAND_111[63:0];
  _RAND_114 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_38[initvar] = _RAND_114[63:0];
  _RAND_117 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_39[initvar] = _RAND_117[63:0];
  _RAND_120 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_40[initvar] = _RAND_120[63:0];
  _RAND_123 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_41[initvar] = _RAND_123[63:0];
  _RAND_126 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_42[initvar] = _RAND_126[63:0];
  _RAND_129 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_43[initvar] = _RAND_129[63:0];
  _RAND_132 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_44[initvar] = _RAND_132[63:0];
  _RAND_135 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_45[initvar] = _RAND_135[63:0];
  _RAND_138 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_46[initvar] = _RAND_138[63:0];
  _RAND_141 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_47[initvar] = _RAND_141[63:0];
  _RAND_144 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_48[initvar] = _RAND_144[63:0];
  _RAND_147 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_49[initvar] = _RAND_147[63:0];
  _RAND_150 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_50[initvar] = _RAND_150[63:0];
  _RAND_153 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_51[initvar] = _RAND_153[63:0];
  _RAND_156 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_52[initvar] = _RAND_156[63:0];
  _RAND_159 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_53[initvar] = _RAND_159[63:0];
  _RAND_162 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_54[initvar] = _RAND_162[63:0];
  _RAND_165 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_55[initvar] = _RAND_165[63:0];
  _RAND_168 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_56[initvar] = _RAND_168[63:0];
  _RAND_171 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_57[initvar] = _RAND_171[63:0];
  _RAND_174 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_58[initvar] = _RAND_174[63:0];
  _RAND_177 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_59[initvar] = _RAND_177[63:0];
  _RAND_180 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_60[initvar] = _RAND_180[63:0];
  _RAND_183 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_61[initvar] = _RAND_183[63:0];
  _RAND_186 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_62[initvar] = _RAND_186[63:0];
  _RAND_189 = {2{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_63[initvar] = _RAND_189[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tensorFile_0_MPORT_64_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  tensorFile_0_MPORT_64_addr_pipe_0 = _RAND_2[5:0];
  _RAND_4 = {1{`RANDOM}};
  tensorFile_1_MPORT_65_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  tensorFile_1_MPORT_65_addr_pipe_0 = _RAND_5[5:0];
  _RAND_7 = {1{`RANDOM}};
  tensorFile_2_MPORT_66_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  tensorFile_2_MPORT_66_addr_pipe_0 = _RAND_8[5:0];
  _RAND_10 = {1{`RANDOM}};
  tensorFile_3_MPORT_67_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  tensorFile_3_MPORT_67_addr_pipe_0 = _RAND_11[5:0];
  _RAND_13 = {1{`RANDOM}};
  tensorFile_4_MPORT_68_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  tensorFile_4_MPORT_68_addr_pipe_0 = _RAND_14[5:0];
  _RAND_16 = {1{`RANDOM}};
  tensorFile_5_MPORT_69_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  tensorFile_5_MPORT_69_addr_pipe_0 = _RAND_17[5:0];
  _RAND_19 = {1{`RANDOM}};
  tensorFile_6_MPORT_70_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  tensorFile_6_MPORT_70_addr_pipe_0 = _RAND_20[5:0];
  _RAND_22 = {1{`RANDOM}};
  tensorFile_7_MPORT_71_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  tensorFile_7_MPORT_71_addr_pipe_0 = _RAND_23[5:0];
  _RAND_25 = {1{`RANDOM}};
  tensorFile_8_MPORT_72_en_pipe_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  tensorFile_8_MPORT_72_addr_pipe_0 = _RAND_26[5:0];
  _RAND_28 = {1{`RANDOM}};
  tensorFile_9_MPORT_73_en_pipe_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  tensorFile_9_MPORT_73_addr_pipe_0 = _RAND_29[5:0];
  _RAND_31 = {1{`RANDOM}};
  tensorFile_10_MPORT_74_en_pipe_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  tensorFile_10_MPORT_74_addr_pipe_0 = _RAND_32[5:0];
  _RAND_34 = {1{`RANDOM}};
  tensorFile_11_MPORT_75_en_pipe_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  tensorFile_11_MPORT_75_addr_pipe_0 = _RAND_35[5:0];
  _RAND_37 = {1{`RANDOM}};
  tensorFile_12_MPORT_76_en_pipe_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  tensorFile_12_MPORT_76_addr_pipe_0 = _RAND_38[5:0];
  _RAND_40 = {1{`RANDOM}};
  tensorFile_13_MPORT_77_en_pipe_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  tensorFile_13_MPORT_77_addr_pipe_0 = _RAND_41[5:0];
  _RAND_43 = {1{`RANDOM}};
  tensorFile_14_MPORT_78_en_pipe_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  tensorFile_14_MPORT_78_addr_pipe_0 = _RAND_44[5:0];
  _RAND_46 = {1{`RANDOM}};
  tensorFile_15_MPORT_79_en_pipe_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  tensorFile_15_MPORT_79_addr_pipe_0 = _RAND_47[5:0];
  _RAND_49 = {1{`RANDOM}};
  tensorFile_16_MPORT_80_en_pipe_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  tensorFile_16_MPORT_80_addr_pipe_0 = _RAND_50[5:0];
  _RAND_52 = {1{`RANDOM}};
  tensorFile_17_MPORT_81_en_pipe_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  tensorFile_17_MPORT_81_addr_pipe_0 = _RAND_53[5:0];
  _RAND_55 = {1{`RANDOM}};
  tensorFile_18_MPORT_82_en_pipe_0 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  tensorFile_18_MPORT_82_addr_pipe_0 = _RAND_56[5:0];
  _RAND_58 = {1{`RANDOM}};
  tensorFile_19_MPORT_83_en_pipe_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  tensorFile_19_MPORT_83_addr_pipe_0 = _RAND_59[5:0];
  _RAND_61 = {1{`RANDOM}};
  tensorFile_20_MPORT_84_en_pipe_0 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  tensorFile_20_MPORT_84_addr_pipe_0 = _RAND_62[5:0];
  _RAND_64 = {1{`RANDOM}};
  tensorFile_21_MPORT_85_en_pipe_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  tensorFile_21_MPORT_85_addr_pipe_0 = _RAND_65[5:0];
  _RAND_67 = {1{`RANDOM}};
  tensorFile_22_MPORT_86_en_pipe_0 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  tensorFile_22_MPORT_86_addr_pipe_0 = _RAND_68[5:0];
  _RAND_70 = {1{`RANDOM}};
  tensorFile_23_MPORT_87_en_pipe_0 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  tensorFile_23_MPORT_87_addr_pipe_0 = _RAND_71[5:0];
  _RAND_73 = {1{`RANDOM}};
  tensorFile_24_MPORT_88_en_pipe_0 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  tensorFile_24_MPORT_88_addr_pipe_0 = _RAND_74[5:0];
  _RAND_76 = {1{`RANDOM}};
  tensorFile_25_MPORT_89_en_pipe_0 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  tensorFile_25_MPORT_89_addr_pipe_0 = _RAND_77[5:0];
  _RAND_79 = {1{`RANDOM}};
  tensorFile_26_MPORT_90_en_pipe_0 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  tensorFile_26_MPORT_90_addr_pipe_0 = _RAND_80[5:0];
  _RAND_82 = {1{`RANDOM}};
  tensorFile_27_MPORT_91_en_pipe_0 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  tensorFile_27_MPORT_91_addr_pipe_0 = _RAND_83[5:0];
  _RAND_85 = {1{`RANDOM}};
  tensorFile_28_MPORT_92_en_pipe_0 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  tensorFile_28_MPORT_92_addr_pipe_0 = _RAND_86[5:0];
  _RAND_88 = {1{`RANDOM}};
  tensorFile_29_MPORT_93_en_pipe_0 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  tensorFile_29_MPORT_93_addr_pipe_0 = _RAND_89[5:0];
  _RAND_91 = {1{`RANDOM}};
  tensorFile_30_MPORT_94_en_pipe_0 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  tensorFile_30_MPORT_94_addr_pipe_0 = _RAND_92[5:0];
  _RAND_94 = {1{`RANDOM}};
  tensorFile_31_MPORT_95_en_pipe_0 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  tensorFile_31_MPORT_95_addr_pipe_0 = _RAND_95[5:0];
  _RAND_97 = {1{`RANDOM}};
  tensorFile_32_MPORT_96_en_pipe_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  tensorFile_32_MPORT_96_addr_pipe_0 = _RAND_98[5:0];
  _RAND_100 = {1{`RANDOM}};
  tensorFile_33_MPORT_97_en_pipe_0 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  tensorFile_33_MPORT_97_addr_pipe_0 = _RAND_101[5:0];
  _RAND_103 = {1{`RANDOM}};
  tensorFile_34_MPORT_98_en_pipe_0 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  tensorFile_34_MPORT_98_addr_pipe_0 = _RAND_104[5:0];
  _RAND_106 = {1{`RANDOM}};
  tensorFile_35_MPORT_99_en_pipe_0 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  tensorFile_35_MPORT_99_addr_pipe_0 = _RAND_107[5:0];
  _RAND_109 = {1{`RANDOM}};
  tensorFile_36_MPORT_100_en_pipe_0 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  tensorFile_36_MPORT_100_addr_pipe_0 = _RAND_110[5:0];
  _RAND_112 = {1{`RANDOM}};
  tensorFile_37_MPORT_101_en_pipe_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  tensorFile_37_MPORT_101_addr_pipe_0 = _RAND_113[5:0];
  _RAND_115 = {1{`RANDOM}};
  tensorFile_38_MPORT_102_en_pipe_0 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  tensorFile_38_MPORT_102_addr_pipe_0 = _RAND_116[5:0];
  _RAND_118 = {1{`RANDOM}};
  tensorFile_39_MPORT_103_en_pipe_0 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  tensorFile_39_MPORT_103_addr_pipe_0 = _RAND_119[5:0];
  _RAND_121 = {1{`RANDOM}};
  tensorFile_40_MPORT_104_en_pipe_0 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  tensorFile_40_MPORT_104_addr_pipe_0 = _RAND_122[5:0];
  _RAND_124 = {1{`RANDOM}};
  tensorFile_41_MPORT_105_en_pipe_0 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  tensorFile_41_MPORT_105_addr_pipe_0 = _RAND_125[5:0];
  _RAND_127 = {1{`RANDOM}};
  tensorFile_42_MPORT_106_en_pipe_0 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  tensorFile_42_MPORT_106_addr_pipe_0 = _RAND_128[5:0];
  _RAND_130 = {1{`RANDOM}};
  tensorFile_43_MPORT_107_en_pipe_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  tensorFile_43_MPORT_107_addr_pipe_0 = _RAND_131[5:0];
  _RAND_133 = {1{`RANDOM}};
  tensorFile_44_MPORT_108_en_pipe_0 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  tensorFile_44_MPORT_108_addr_pipe_0 = _RAND_134[5:0];
  _RAND_136 = {1{`RANDOM}};
  tensorFile_45_MPORT_109_en_pipe_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  tensorFile_45_MPORT_109_addr_pipe_0 = _RAND_137[5:0];
  _RAND_139 = {1{`RANDOM}};
  tensorFile_46_MPORT_110_en_pipe_0 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  tensorFile_46_MPORT_110_addr_pipe_0 = _RAND_140[5:0];
  _RAND_142 = {1{`RANDOM}};
  tensorFile_47_MPORT_111_en_pipe_0 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  tensorFile_47_MPORT_111_addr_pipe_0 = _RAND_143[5:0];
  _RAND_145 = {1{`RANDOM}};
  tensorFile_48_MPORT_112_en_pipe_0 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  tensorFile_48_MPORT_112_addr_pipe_0 = _RAND_146[5:0];
  _RAND_148 = {1{`RANDOM}};
  tensorFile_49_MPORT_113_en_pipe_0 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  tensorFile_49_MPORT_113_addr_pipe_0 = _RAND_149[5:0];
  _RAND_151 = {1{`RANDOM}};
  tensorFile_50_MPORT_114_en_pipe_0 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  tensorFile_50_MPORT_114_addr_pipe_0 = _RAND_152[5:0];
  _RAND_154 = {1{`RANDOM}};
  tensorFile_51_MPORT_115_en_pipe_0 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  tensorFile_51_MPORT_115_addr_pipe_0 = _RAND_155[5:0];
  _RAND_157 = {1{`RANDOM}};
  tensorFile_52_MPORT_116_en_pipe_0 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  tensorFile_52_MPORT_116_addr_pipe_0 = _RAND_158[5:0];
  _RAND_160 = {1{`RANDOM}};
  tensorFile_53_MPORT_117_en_pipe_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  tensorFile_53_MPORT_117_addr_pipe_0 = _RAND_161[5:0];
  _RAND_163 = {1{`RANDOM}};
  tensorFile_54_MPORT_118_en_pipe_0 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  tensorFile_54_MPORT_118_addr_pipe_0 = _RAND_164[5:0];
  _RAND_166 = {1{`RANDOM}};
  tensorFile_55_MPORT_119_en_pipe_0 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  tensorFile_55_MPORT_119_addr_pipe_0 = _RAND_167[5:0];
  _RAND_169 = {1{`RANDOM}};
  tensorFile_56_MPORT_120_en_pipe_0 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  tensorFile_56_MPORT_120_addr_pipe_0 = _RAND_170[5:0];
  _RAND_172 = {1{`RANDOM}};
  tensorFile_57_MPORT_121_en_pipe_0 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  tensorFile_57_MPORT_121_addr_pipe_0 = _RAND_173[5:0];
  _RAND_175 = {1{`RANDOM}};
  tensorFile_58_MPORT_122_en_pipe_0 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  tensorFile_58_MPORT_122_addr_pipe_0 = _RAND_176[5:0];
  _RAND_178 = {1{`RANDOM}};
  tensorFile_59_MPORT_123_en_pipe_0 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  tensorFile_59_MPORT_123_addr_pipe_0 = _RAND_179[5:0];
  _RAND_181 = {1{`RANDOM}};
  tensorFile_60_MPORT_124_en_pipe_0 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  tensorFile_60_MPORT_124_addr_pipe_0 = _RAND_182[5:0];
  _RAND_184 = {1{`RANDOM}};
  tensorFile_61_MPORT_125_en_pipe_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  tensorFile_61_MPORT_125_addr_pipe_0 = _RAND_185[5:0];
  _RAND_187 = {1{`RANDOM}};
  tensorFile_62_MPORT_126_en_pipe_0 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  tensorFile_62_MPORT_126_addr_pipe_0 = _RAND_188[5:0];
  _RAND_190 = {1{`RANDOM}};
  tensorFile_63_MPORT_127_en_pipe_0 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  tensorFile_63_MPORT_127_addr_pipe_0 = _RAND_191[5:0];
  _RAND_192 = {1{`RANDOM}};
  state = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  blocksInFlight = _RAND_193[11:0];
  _RAND_194 = {2{`RANDOM}};
  vmeDataBitsPipe_data = _RAND_194[63:0];
  _RAND_195 = {1{`RANDOM}};
  vmeDataBitsPipe_tag = _RAND_195[20:0];
  _RAND_196 = {1{`RANDOM}};
  vmeDataValidPipe = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  vmeDataReadyPipe = _RAND_197[0:0];
  _RAND_198 = {4{`RANDOM}};
  fillPadding_io_inst_REG = _RAND_198[127:0];
  _RAND_199 = {1{`RANDOM}};
  fillPadding_io_start_REG = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  rvalid = _RAND_200[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~io_start & ~_T_3 & ~_T_6 & _T_10 & ~reset) begin
      assert(blocksInFlight > 12'h0); // @[TensorLoadNarrowVME.scala 95:11]
    end
    //
    if (_T_13) begin
      assert(1'h1); // @[TensorLoadNarrowVME.scala 109:9]
    end
  end
endmodule
module TensorLoadWgt(
  input          clock,
  input          reset,
  input          io_start,
  output         io_done,
  input  [127:0] io_inst,
  input  [31:0]  io_baddr,
  input          io_vme_rd_cmd_ready,
  output         io_vme_rd_cmd_valid,
  output [31:0]  io_vme_rd_cmd_bits_addr,
  output [3:0]   io_vme_rd_cmd_bits_len,
  output [20:0]  io_vme_rd_cmd_bits_tag,
  input          io_vme_rd_data_valid,
  input  [63:0]  io_vme_rd_data_bits_data,
  input  [20:0]  io_vme_rd_data_bits_tag,
  input          io_tensor_rd_0_idx_valid,
  input  [5:0]   io_tensor_rd_0_idx_bits,
  output         io_tensor_rd_0_data_valid,
  output [7:0]   io_tensor_rd_0_data_bits_0_0,
  output [7:0]   io_tensor_rd_0_data_bits_0_1,
  output [7:0]   io_tensor_rd_0_data_bits_0_2,
  output [7:0]   io_tensor_rd_0_data_bits_0_3,
  output [7:0]   io_tensor_rd_0_data_bits_0_4,
  output [7:0]   io_tensor_rd_0_data_bits_0_5,
  output [7:0]   io_tensor_rd_0_data_bits_0_6,
  output [7:0]   io_tensor_rd_0_data_bits_0_7,
  output [7:0]   io_tensor_rd_0_data_bits_0_8,
  output [7:0]   io_tensor_rd_0_data_bits_0_9,
  output [7:0]   io_tensor_rd_0_data_bits_0_10,
  output [7:0]   io_tensor_rd_0_data_bits_0_11,
  output [7:0]   io_tensor_rd_0_data_bits_0_12,
  output [7:0]   io_tensor_rd_0_data_bits_0_13,
  output [7:0]   io_tensor_rd_0_data_bits_0_14,
  output [7:0]   io_tensor_rd_0_data_bits_0_15,
  output [7:0]   io_tensor_rd_0_data_bits_1_0,
  output [7:0]   io_tensor_rd_0_data_bits_1_1,
  output [7:0]   io_tensor_rd_0_data_bits_1_2,
  output [7:0]   io_tensor_rd_0_data_bits_1_3,
  output [7:0]   io_tensor_rd_0_data_bits_1_4,
  output [7:0]   io_tensor_rd_0_data_bits_1_5,
  output [7:0]   io_tensor_rd_0_data_bits_1_6,
  output [7:0]   io_tensor_rd_0_data_bits_1_7,
  output [7:0]   io_tensor_rd_0_data_bits_1_8,
  output [7:0]   io_tensor_rd_0_data_bits_1_9,
  output [7:0]   io_tensor_rd_0_data_bits_1_10,
  output [7:0]   io_tensor_rd_0_data_bits_1_11,
  output [7:0]   io_tensor_rd_0_data_bits_1_12,
  output [7:0]   io_tensor_rd_0_data_bits_1_13,
  output [7:0]   io_tensor_rd_0_data_bits_1_14,
  output [7:0]   io_tensor_rd_0_data_bits_1_15,
  output [7:0]   io_tensor_rd_0_data_bits_2_0,
  output [7:0]   io_tensor_rd_0_data_bits_2_1,
  output [7:0]   io_tensor_rd_0_data_bits_2_2,
  output [7:0]   io_tensor_rd_0_data_bits_2_3,
  output [7:0]   io_tensor_rd_0_data_bits_2_4,
  output [7:0]   io_tensor_rd_0_data_bits_2_5,
  output [7:0]   io_tensor_rd_0_data_bits_2_6,
  output [7:0]   io_tensor_rd_0_data_bits_2_7,
  output [7:0]   io_tensor_rd_0_data_bits_2_8,
  output [7:0]   io_tensor_rd_0_data_bits_2_9,
  output [7:0]   io_tensor_rd_0_data_bits_2_10,
  output [7:0]   io_tensor_rd_0_data_bits_2_11,
  output [7:0]   io_tensor_rd_0_data_bits_2_12,
  output [7:0]   io_tensor_rd_0_data_bits_2_13,
  output [7:0]   io_tensor_rd_0_data_bits_2_14,
  output [7:0]   io_tensor_rd_0_data_bits_2_15,
  output [7:0]   io_tensor_rd_0_data_bits_3_0,
  output [7:0]   io_tensor_rd_0_data_bits_3_1,
  output [7:0]   io_tensor_rd_0_data_bits_3_2,
  output [7:0]   io_tensor_rd_0_data_bits_3_3,
  output [7:0]   io_tensor_rd_0_data_bits_3_4,
  output [7:0]   io_tensor_rd_0_data_bits_3_5,
  output [7:0]   io_tensor_rd_0_data_bits_3_6,
  output [7:0]   io_tensor_rd_0_data_bits_3_7,
  output [7:0]   io_tensor_rd_0_data_bits_3_8,
  output [7:0]   io_tensor_rd_0_data_bits_3_9,
  output [7:0]   io_tensor_rd_0_data_bits_3_10,
  output [7:0]   io_tensor_rd_0_data_bits_3_11,
  output [7:0]   io_tensor_rd_0_data_bits_3_12,
  output [7:0]   io_tensor_rd_0_data_bits_3_13,
  output [7:0]   io_tensor_rd_0_data_bits_3_14,
  output [7:0]   io_tensor_rd_0_data_bits_3_15,
  output [7:0]   io_tensor_rd_0_data_bits_4_0,
  output [7:0]   io_tensor_rd_0_data_bits_4_1,
  output [7:0]   io_tensor_rd_0_data_bits_4_2,
  output [7:0]   io_tensor_rd_0_data_bits_4_3,
  output [7:0]   io_tensor_rd_0_data_bits_4_4,
  output [7:0]   io_tensor_rd_0_data_bits_4_5,
  output [7:0]   io_tensor_rd_0_data_bits_4_6,
  output [7:0]   io_tensor_rd_0_data_bits_4_7,
  output [7:0]   io_tensor_rd_0_data_bits_4_8,
  output [7:0]   io_tensor_rd_0_data_bits_4_9,
  output [7:0]   io_tensor_rd_0_data_bits_4_10,
  output [7:0]   io_tensor_rd_0_data_bits_4_11,
  output [7:0]   io_tensor_rd_0_data_bits_4_12,
  output [7:0]   io_tensor_rd_0_data_bits_4_13,
  output [7:0]   io_tensor_rd_0_data_bits_4_14,
  output [7:0]   io_tensor_rd_0_data_bits_4_15,
  output [7:0]   io_tensor_rd_0_data_bits_5_0,
  output [7:0]   io_tensor_rd_0_data_bits_5_1,
  output [7:0]   io_tensor_rd_0_data_bits_5_2,
  output [7:0]   io_tensor_rd_0_data_bits_5_3,
  output [7:0]   io_tensor_rd_0_data_bits_5_4,
  output [7:0]   io_tensor_rd_0_data_bits_5_5,
  output [7:0]   io_tensor_rd_0_data_bits_5_6,
  output [7:0]   io_tensor_rd_0_data_bits_5_7,
  output [7:0]   io_tensor_rd_0_data_bits_5_8,
  output [7:0]   io_tensor_rd_0_data_bits_5_9,
  output [7:0]   io_tensor_rd_0_data_bits_5_10,
  output [7:0]   io_tensor_rd_0_data_bits_5_11,
  output [7:0]   io_tensor_rd_0_data_bits_5_12,
  output [7:0]   io_tensor_rd_0_data_bits_5_13,
  output [7:0]   io_tensor_rd_0_data_bits_5_14,
  output [7:0]   io_tensor_rd_0_data_bits_5_15,
  output [7:0]   io_tensor_rd_0_data_bits_6_0,
  output [7:0]   io_tensor_rd_0_data_bits_6_1,
  output [7:0]   io_tensor_rd_0_data_bits_6_2,
  output [7:0]   io_tensor_rd_0_data_bits_6_3,
  output [7:0]   io_tensor_rd_0_data_bits_6_4,
  output [7:0]   io_tensor_rd_0_data_bits_6_5,
  output [7:0]   io_tensor_rd_0_data_bits_6_6,
  output [7:0]   io_tensor_rd_0_data_bits_6_7,
  output [7:0]   io_tensor_rd_0_data_bits_6_8,
  output [7:0]   io_tensor_rd_0_data_bits_6_9,
  output [7:0]   io_tensor_rd_0_data_bits_6_10,
  output [7:0]   io_tensor_rd_0_data_bits_6_11,
  output [7:0]   io_tensor_rd_0_data_bits_6_12,
  output [7:0]   io_tensor_rd_0_data_bits_6_13,
  output [7:0]   io_tensor_rd_0_data_bits_6_14,
  output [7:0]   io_tensor_rd_0_data_bits_6_15,
  output [7:0]   io_tensor_rd_0_data_bits_7_0,
  output [7:0]   io_tensor_rd_0_data_bits_7_1,
  output [7:0]   io_tensor_rd_0_data_bits_7_2,
  output [7:0]   io_tensor_rd_0_data_bits_7_3,
  output [7:0]   io_tensor_rd_0_data_bits_7_4,
  output [7:0]   io_tensor_rd_0_data_bits_7_5,
  output [7:0]   io_tensor_rd_0_data_bits_7_6,
  output [7:0]   io_tensor_rd_0_data_bits_7_7,
  output [7:0]   io_tensor_rd_0_data_bits_7_8,
  output [7:0]   io_tensor_rd_0_data_bits_7_9,
  output [7:0]   io_tensor_rd_0_data_bits_7_10,
  output [7:0]   io_tensor_rd_0_data_bits_7_11,
  output [7:0]   io_tensor_rd_0_data_bits_7_12,
  output [7:0]   io_tensor_rd_0_data_bits_7_13,
  output [7:0]   io_tensor_rd_0_data_bits_7_14,
  output [7:0]   io_tensor_rd_0_data_bits_7_15,
  output [7:0]   io_tensor_rd_0_data_bits_8_0,
  output [7:0]   io_tensor_rd_0_data_bits_8_1,
  output [7:0]   io_tensor_rd_0_data_bits_8_2,
  output [7:0]   io_tensor_rd_0_data_bits_8_3,
  output [7:0]   io_tensor_rd_0_data_bits_8_4,
  output [7:0]   io_tensor_rd_0_data_bits_8_5,
  output [7:0]   io_tensor_rd_0_data_bits_8_6,
  output [7:0]   io_tensor_rd_0_data_bits_8_7,
  output [7:0]   io_tensor_rd_0_data_bits_8_8,
  output [7:0]   io_tensor_rd_0_data_bits_8_9,
  output [7:0]   io_tensor_rd_0_data_bits_8_10,
  output [7:0]   io_tensor_rd_0_data_bits_8_11,
  output [7:0]   io_tensor_rd_0_data_bits_8_12,
  output [7:0]   io_tensor_rd_0_data_bits_8_13,
  output [7:0]   io_tensor_rd_0_data_bits_8_14,
  output [7:0]   io_tensor_rd_0_data_bits_8_15,
  output [7:0]   io_tensor_rd_0_data_bits_9_0,
  output [7:0]   io_tensor_rd_0_data_bits_9_1,
  output [7:0]   io_tensor_rd_0_data_bits_9_2,
  output [7:0]   io_tensor_rd_0_data_bits_9_3,
  output [7:0]   io_tensor_rd_0_data_bits_9_4,
  output [7:0]   io_tensor_rd_0_data_bits_9_5,
  output [7:0]   io_tensor_rd_0_data_bits_9_6,
  output [7:0]   io_tensor_rd_0_data_bits_9_7,
  output [7:0]   io_tensor_rd_0_data_bits_9_8,
  output [7:0]   io_tensor_rd_0_data_bits_9_9,
  output [7:0]   io_tensor_rd_0_data_bits_9_10,
  output [7:0]   io_tensor_rd_0_data_bits_9_11,
  output [7:0]   io_tensor_rd_0_data_bits_9_12,
  output [7:0]   io_tensor_rd_0_data_bits_9_13,
  output [7:0]   io_tensor_rd_0_data_bits_9_14,
  output [7:0]   io_tensor_rd_0_data_bits_9_15,
  output [7:0]   io_tensor_rd_0_data_bits_10_0,
  output [7:0]   io_tensor_rd_0_data_bits_10_1,
  output [7:0]   io_tensor_rd_0_data_bits_10_2,
  output [7:0]   io_tensor_rd_0_data_bits_10_3,
  output [7:0]   io_tensor_rd_0_data_bits_10_4,
  output [7:0]   io_tensor_rd_0_data_bits_10_5,
  output [7:0]   io_tensor_rd_0_data_bits_10_6,
  output [7:0]   io_tensor_rd_0_data_bits_10_7,
  output [7:0]   io_tensor_rd_0_data_bits_10_8,
  output [7:0]   io_tensor_rd_0_data_bits_10_9,
  output [7:0]   io_tensor_rd_0_data_bits_10_10,
  output [7:0]   io_tensor_rd_0_data_bits_10_11,
  output [7:0]   io_tensor_rd_0_data_bits_10_12,
  output [7:0]   io_tensor_rd_0_data_bits_10_13,
  output [7:0]   io_tensor_rd_0_data_bits_10_14,
  output [7:0]   io_tensor_rd_0_data_bits_10_15,
  output [7:0]   io_tensor_rd_0_data_bits_11_0,
  output [7:0]   io_tensor_rd_0_data_bits_11_1,
  output [7:0]   io_tensor_rd_0_data_bits_11_2,
  output [7:0]   io_tensor_rd_0_data_bits_11_3,
  output [7:0]   io_tensor_rd_0_data_bits_11_4,
  output [7:0]   io_tensor_rd_0_data_bits_11_5,
  output [7:0]   io_tensor_rd_0_data_bits_11_6,
  output [7:0]   io_tensor_rd_0_data_bits_11_7,
  output [7:0]   io_tensor_rd_0_data_bits_11_8,
  output [7:0]   io_tensor_rd_0_data_bits_11_9,
  output [7:0]   io_tensor_rd_0_data_bits_11_10,
  output [7:0]   io_tensor_rd_0_data_bits_11_11,
  output [7:0]   io_tensor_rd_0_data_bits_11_12,
  output [7:0]   io_tensor_rd_0_data_bits_11_13,
  output [7:0]   io_tensor_rd_0_data_bits_11_14,
  output [7:0]   io_tensor_rd_0_data_bits_11_15,
  output [7:0]   io_tensor_rd_0_data_bits_12_0,
  output [7:0]   io_tensor_rd_0_data_bits_12_1,
  output [7:0]   io_tensor_rd_0_data_bits_12_2,
  output [7:0]   io_tensor_rd_0_data_bits_12_3,
  output [7:0]   io_tensor_rd_0_data_bits_12_4,
  output [7:0]   io_tensor_rd_0_data_bits_12_5,
  output [7:0]   io_tensor_rd_0_data_bits_12_6,
  output [7:0]   io_tensor_rd_0_data_bits_12_7,
  output [7:0]   io_tensor_rd_0_data_bits_12_8,
  output [7:0]   io_tensor_rd_0_data_bits_12_9,
  output [7:0]   io_tensor_rd_0_data_bits_12_10,
  output [7:0]   io_tensor_rd_0_data_bits_12_11,
  output [7:0]   io_tensor_rd_0_data_bits_12_12,
  output [7:0]   io_tensor_rd_0_data_bits_12_13,
  output [7:0]   io_tensor_rd_0_data_bits_12_14,
  output [7:0]   io_tensor_rd_0_data_bits_12_15,
  output [7:0]   io_tensor_rd_0_data_bits_13_0,
  output [7:0]   io_tensor_rd_0_data_bits_13_1,
  output [7:0]   io_tensor_rd_0_data_bits_13_2,
  output [7:0]   io_tensor_rd_0_data_bits_13_3,
  output [7:0]   io_tensor_rd_0_data_bits_13_4,
  output [7:0]   io_tensor_rd_0_data_bits_13_5,
  output [7:0]   io_tensor_rd_0_data_bits_13_6,
  output [7:0]   io_tensor_rd_0_data_bits_13_7,
  output [7:0]   io_tensor_rd_0_data_bits_13_8,
  output [7:0]   io_tensor_rd_0_data_bits_13_9,
  output [7:0]   io_tensor_rd_0_data_bits_13_10,
  output [7:0]   io_tensor_rd_0_data_bits_13_11,
  output [7:0]   io_tensor_rd_0_data_bits_13_12,
  output [7:0]   io_tensor_rd_0_data_bits_13_13,
  output [7:0]   io_tensor_rd_0_data_bits_13_14,
  output [7:0]   io_tensor_rd_0_data_bits_13_15,
  output [7:0]   io_tensor_rd_0_data_bits_14_0,
  output [7:0]   io_tensor_rd_0_data_bits_14_1,
  output [7:0]   io_tensor_rd_0_data_bits_14_2,
  output [7:0]   io_tensor_rd_0_data_bits_14_3,
  output [7:0]   io_tensor_rd_0_data_bits_14_4,
  output [7:0]   io_tensor_rd_0_data_bits_14_5,
  output [7:0]   io_tensor_rd_0_data_bits_14_6,
  output [7:0]   io_tensor_rd_0_data_bits_14_7,
  output [7:0]   io_tensor_rd_0_data_bits_14_8,
  output [7:0]   io_tensor_rd_0_data_bits_14_9,
  output [7:0]   io_tensor_rd_0_data_bits_14_10,
  output [7:0]   io_tensor_rd_0_data_bits_14_11,
  output [7:0]   io_tensor_rd_0_data_bits_14_12,
  output [7:0]   io_tensor_rd_0_data_bits_14_13,
  output [7:0]   io_tensor_rd_0_data_bits_14_14,
  output [7:0]   io_tensor_rd_0_data_bits_14_15,
  output [7:0]   io_tensor_rd_0_data_bits_15_0,
  output [7:0]   io_tensor_rd_0_data_bits_15_1,
  output [7:0]   io_tensor_rd_0_data_bits_15_2,
  output [7:0]   io_tensor_rd_0_data_bits_15_3,
  output [7:0]   io_tensor_rd_0_data_bits_15_4,
  output [7:0]   io_tensor_rd_0_data_bits_15_5,
  output [7:0]   io_tensor_rd_0_data_bits_15_6,
  output [7:0]   io_tensor_rd_0_data_bits_15_7,
  output [7:0]   io_tensor_rd_0_data_bits_15_8,
  output [7:0]   io_tensor_rd_0_data_bits_15_9,
  output [7:0]   io_tensor_rd_0_data_bits_15_10,
  output [7:0]   io_tensor_rd_0_data_bits_15_11,
  output [7:0]   io_tensor_rd_0_data_bits_15_12,
  output [7:0]   io_tensor_rd_0_data_bits_15_13,
  output [7:0]   io_tensor_rd_0_data_bits_15_14,
  output [7:0]   io_tensor_rd_0_data_bits_15_15,
  output [7:0]   io_tensor_rd_0_data_bits_16_0,
  output [7:0]   io_tensor_rd_0_data_bits_16_1,
  output [7:0]   io_tensor_rd_0_data_bits_16_2,
  output [7:0]   io_tensor_rd_0_data_bits_16_3,
  output [7:0]   io_tensor_rd_0_data_bits_16_4,
  output [7:0]   io_tensor_rd_0_data_bits_16_5,
  output [7:0]   io_tensor_rd_0_data_bits_16_6,
  output [7:0]   io_tensor_rd_0_data_bits_16_7,
  output [7:0]   io_tensor_rd_0_data_bits_16_8,
  output [7:0]   io_tensor_rd_0_data_bits_16_9,
  output [7:0]   io_tensor_rd_0_data_bits_16_10,
  output [7:0]   io_tensor_rd_0_data_bits_16_11,
  output [7:0]   io_tensor_rd_0_data_bits_16_12,
  output [7:0]   io_tensor_rd_0_data_bits_16_13,
  output [7:0]   io_tensor_rd_0_data_bits_16_14,
  output [7:0]   io_tensor_rd_0_data_bits_16_15,
  output [7:0]   io_tensor_rd_0_data_bits_17_0,
  output [7:0]   io_tensor_rd_0_data_bits_17_1,
  output [7:0]   io_tensor_rd_0_data_bits_17_2,
  output [7:0]   io_tensor_rd_0_data_bits_17_3,
  output [7:0]   io_tensor_rd_0_data_bits_17_4,
  output [7:0]   io_tensor_rd_0_data_bits_17_5,
  output [7:0]   io_tensor_rd_0_data_bits_17_6,
  output [7:0]   io_tensor_rd_0_data_bits_17_7,
  output [7:0]   io_tensor_rd_0_data_bits_17_8,
  output [7:0]   io_tensor_rd_0_data_bits_17_9,
  output [7:0]   io_tensor_rd_0_data_bits_17_10,
  output [7:0]   io_tensor_rd_0_data_bits_17_11,
  output [7:0]   io_tensor_rd_0_data_bits_17_12,
  output [7:0]   io_tensor_rd_0_data_bits_17_13,
  output [7:0]   io_tensor_rd_0_data_bits_17_14,
  output [7:0]   io_tensor_rd_0_data_bits_17_15,
  output [7:0]   io_tensor_rd_0_data_bits_18_0,
  output [7:0]   io_tensor_rd_0_data_bits_18_1,
  output [7:0]   io_tensor_rd_0_data_bits_18_2,
  output [7:0]   io_tensor_rd_0_data_bits_18_3,
  output [7:0]   io_tensor_rd_0_data_bits_18_4,
  output [7:0]   io_tensor_rd_0_data_bits_18_5,
  output [7:0]   io_tensor_rd_0_data_bits_18_6,
  output [7:0]   io_tensor_rd_0_data_bits_18_7,
  output [7:0]   io_tensor_rd_0_data_bits_18_8,
  output [7:0]   io_tensor_rd_0_data_bits_18_9,
  output [7:0]   io_tensor_rd_0_data_bits_18_10,
  output [7:0]   io_tensor_rd_0_data_bits_18_11,
  output [7:0]   io_tensor_rd_0_data_bits_18_12,
  output [7:0]   io_tensor_rd_0_data_bits_18_13,
  output [7:0]   io_tensor_rd_0_data_bits_18_14,
  output [7:0]   io_tensor_rd_0_data_bits_18_15,
  output [7:0]   io_tensor_rd_0_data_bits_19_0,
  output [7:0]   io_tensor_rd_0_data_bits_19_1,
  output [7:0]   io_tensor_rd_0_data_bits_19_2,
  output [7:0]   io_tensor_rd_0_data_bits_19_3,
  output [7:0]   io_tensor_rd_0_data_bits_19_4,
  output [7:0]   io_tensor_rd_0_data_bits_19_5,
  output [7:0]   io_tensor_rd_0_data_bits_19_6,
  output [7:0]   io_tensor_rd_0_data_bits_19_7,
  output [7:0]   io_tensor_rd_0_data_bits_19_8,
  output [7:0]   io_tensor_rd_0_data_bits_19_9,
  output [7:0]   io_tensor_rd_0_data_bits_19_10,
  output [7:0]   io_tensor_rd_0_data_bits_19_11,
  output [7:0]   io_tensor_rd_0_data_bits_19_12,
  output [7:0]   io_tensor_rd_0_data_bits_19_13,
  output [7:0]   io_tensor_rd_0_data_bits_19_14,
  output [7:0]   io_tensor_rd_0_data_bits_19_15,
  output [7:0]   io_tensor_rd_0_data_bits_20_0,
  output [7:0]   io_tensor_rd_0_data_bits_20_1,
  output [7:0]   io_tensor_rd_0_data_bits_20_2,
  output [7:0]   io_tensor_rd_0_data_bits_20_3,
  output [7:0]   io_tensor_rd_0_data_bits_20_4,
  output [7:0]   io_tensor_rd_0_data_bits_20_5,
  output [7:0]   io_tensor_rd_0_data_bits_20_6,
  output [7:0]   io_tensor_rd_0_data_bits_20_7,
  output [7:0]   io_tensor_rd_0_data_bits_20_8,
  output [7:0]   io_tensor_rd_0_data_bits_20_9,
  output [7:0]   io_tensor_rd_0_data_bits_20_10,
  output [7:0]   io_tensor_rd_0_data_bits_20_11,
  output [7:0]   io_tensor_rd_0_data_bits_20_12,
  output [7:0]   io_tensor_rd_0_data_bits_20_13,
  output [7:0]   io_tensor_rd_0_data_bits_20_14,
  output [7:0]   io_tensor_rd_0_data_bits_20_15,
  output [7:0]   io_tensor_rd_0_data_bits_21_0,
  output [7:0]   io_tensor_rd_0_data_bits_21_1,
  output [7:0]   io_tensor_rd_0_data_bits_21_2,
  output [7:0]   io_tensor_rd_0_data_bits_21_3,
  output [7:0]   io_tensor_rd_0_data_bits_21_4,
  output [7:0]   io_tensor_rd_0_data_bits_21_5,
  output [7:0]   io_tensor_rd_0_data_bits_21_6,
  output [7:0]   io_tensor_rd_0_data_bits_21_7,
  output [7:0]   io_tensor_rd_0_data_bits_21_8,
  output [7:0]   io_tensor_rd_0_data_bits_21_9,
  output [7:0]   io_tensor_rd_0_data_bits_21_10,
  output [7:0]   io_tensor_rd_0_data_bits_21_11,
  output [7:0]   io_tensor_rd_0_data_bits_21_12,
  output [7:0]   io_tensor_rd_0_data_bits_21_13,
  output [7:0]   io_tensor_rd_0_data_bits_21_14,
  output [7:0]   io_tensor_rd_0_data_bits_21_15,
  output [7:0]   io_tensor_rd_0_data_bits_22_0,
  output [7:0]   io_tensor_rd_0_data_bits_22_1,
  output [7:0]   io_tensor_rd_0_data_bits_22_2,
  output [7:0]   io_tensor_rd_0_data_bits_22_3,
  output [7:0]   io_tensor_rd_0_data_bits_22_4,
  output [7:0]   io_tensor_rd_0_data_bits_22_5,
  output [7:0]   io_tensor_rd_0_data_bits_22_6,
  output [7:0]   io_tensor_rd_0_data_bits_22_7,
  output [7:0]   io_tensor_rd_0_data_bits_22_8,
  output [7:0]   io_tensor_rd_0_data_bits_22_9,
  output [7:0]   io_tensor_rd_0_data_bits_22_10,
  output [7:0]   io_tensor_rd_0_data_bits_22_11,
  output [7:0]   io_tensor_rd_0_data_bits_22_12,
  output [7:0]   io_tensor_rd_0_data_bits_22_13,
  output [7:0]   io_tensor_rd_0_data_bits_22_14,
  output [7:0]   io_tensor_rd_0_data_bits_22_15,
  output [7:0]   io_tensor_rd_0_data_bits_23_0,
  output [7:0]   io_tensor_rd_0_data_bits_23_1,
  output [7:0]   io_tensor_rd_0_data_bits_23_2,
  output [7:0]   io_tensor_rd_0_data_bits_23_3,
  output [7:0]   io_tensor_rd_0_data_bits_23_4,
  output [7:0]   io_tensor_rd_0_data_bits_23_5,
  output [7:0]   io_tensor_rd_0_data_bits_23_6,
  output [7:0]   io_tensor_rd_0_data_bits_23_7,
  output [7:0]   io_tensor_rd_0_data_bits_23_8,
  output [7:0]   io_tensor_rd_0_data_bits_23_9,
  output [7:0]   io_tensor_rd_0_data_bits_23_10,
  output [7:0]   io_tensor_rd_0_data_bits_23_11,
  output [7:0]   io_tensor_rd_0_data_bits_23_12,
  output [7:0]   io_tensor_rd_0_data_bits_23_13,
  output [7:0]   io_tensor_rd_0_data_bits_23_14,
  output [7:0]   io_tensor_rd_0_data_bits_23_15,
  output [7:0]   io_tensor_rd_0_data_bits_24_0,
  output [7:0]   io_tensor_rd_0_data_bits_24_1,
  output [7:0]   io_tensor_rd_0_data_bits_24_2,
  output [7:0]   io_tensor_rd_0_data_bits_24_3,
  output [7:0]   io_tensor_rd_0_data_bits_24_4,
  output [7:0]   io_tensor_rd_0_data_bits_24_5,
  output [7:0]   io_tensor_rd_0_data_bits_24_6,
  output [7:0]   io_tensor_rd_0_data_bits_24_7,
  output [7:0]   io_tensor_rd_0_data_bits_24_8,
  output [7:0]   io_tensor_rd_0_data_bits_24_9,
  output [7:0]   io_tensor_rd_0_data_bits_24_10,
  output [7:0]   io_tensor_rd_0_data_bits_24_11,
  output [7:0]   io_tensor_rd_0_data_bits_24_12,
  output [7:0]   io_tensor_rd_0_data_bits_24_13,
  output [7:0]   io_tensor_rd_0_data_bits_24_14,
  output [7:0]   io_tensor_rd_0_data_bits_24_15,
  output [7:0]   io_tensor_rd_0_data_bits_25_0,
  output [7:0]   io_tensor_rd_0_data_bits_25_1,
  output [7:0]   io_tensor_rd_0_data_bits_25_2,
  output [7:0]   io_tensor_rd_0_data_bits_25_3,
  output [7:0]   io_tensor_rd_0_data_bits_25_4,
  output [7:0]   io_tensor_rd_0_data_bits_25_5,
  output [7:0]   io_tensor_rd_0_data_bits_25_6,
  output [7:0]   io_tensor_rd_0_data_bits_25_7,
  output [7:0]   io_tensor_rd_0_data_bits_25_8,
  output [7:0]   io_tensor_rd_0_data_bits_25_9,
  output [7:0]   io_tensor_rd_0_data_bits_25_10,
  output [7:0]   io_tensor_rd_0_data_bits_25_11,
  output [7:0]   io_tensor_rd_0_data_bits_25_12,
  output [7:0]   io_tensor_rd_0_data_bits_25_13,
  output [7:0]   io_tensor_rd_0_data_bits_25_14,
  output [7:0]   io_tensor_rd_0_data_bits_25_15,
  output [7:0]   io_tensor_rd_0_data_bits_26_0,
  output [7:0]   io_tensor_rd_0_data_bits_26_1,
  output [7:0]   io_tensor_rd_0_data_bits_26_2,
  output [7:0]   io_tensor_rd_0_data_bits_26_3,
  output [7:0]   io_tensor_rd_0_data_bits_26_4,
  output [7:0]   io_tensor_rd_0_data_bits_26_5,
  output [7:0]   io_tensor_rd_0_data_bits_26_6,
  output [7:0]   io_tensor_rd_0_data_bits_26_7,
  output [7:0]   io_tensor_rd_0_data_bits_26_8,
  output [7:0]   io_tensor_rd_0_data_bits_26_9,
  output [7:0]   io_tensor_rd_0_data_bits_26_10,
  output [7:0]   io_tensor_rd_0_data_bits_26_11,
  output [7:0]   io_tensor_rd_0_data_bits_26_12,
  output [7:0]   io_tensor_rd_0_data_bits_26_13,
  output [7:0]   io_tensor_rd_0_data_bits_26_14,
  output [7:0]   io_tensor_rd_0_data_bits_26_15,
  output [7:0]   io_tensor_rd_0_data_bits_27_0,
  output [7:0]   io_tensor_rd_0_data_bits_27_1,
  output [7:0]   io_tensor_rd_0_data_bits_27_2,
  output [7:0]   io_tensor_rd_0_data_bits_27_3,
  output [7:0]   io_tensor_rd_0_data_bits_27_4,
  output [7:0]   io_tensor_rd_0_data_bits_27_5,
  output [7:0]   io_tensor_rd_0_data_bits_27_6,
  output [7:0]   io_tensor_rd_0_data_bits_27_7,
  output [7:0]   io_tensor_rd_0_data_bits_27_8,
  output [7:0]   io_tensor_rd_0_data_bits_27_9,
  output [7:0]   io_tensor_rd_0_data_bits_27_10,
  output [7:0]   io_tensor_rd_0_data_bits_27_11,
  output [7:0]   io_tensor_rd_0_data_bits_27_12,
  output [7:0]   io_tensor_rd_0_data_bits_27_13,
  output [7:0]   io_tensor_rd_0_data_bits_27_14,
  output [7:0]   io_tensor_rd_0_data_bits_27_15,
  output [7:0]   io_tensor_rd_0_data_bits_28_0,
  output [7:0]   io_tensor_rd_0_data_bits_28_1,
  output [7:0]   io_tensor_rd_0_data_bits_28_2,
  output [7:0]   io_tensor_rd_0_data_bits_28_3,
  output [7:0]   io_tensor_rd_0_data_bits_28_4,
  output [7:0]   io_tensor_rd_0_data_bits_28_5,
  output [7:0]   io_tensor_rd_0_data_bits_28_6,
  output [7:0]   io_tensor_rd_0_data_bits_28_7,
  output [7:0]   io_tensor_rd_0_data_bits_28_8,
  output [7:0]   io_tensor_rd_0_data_bits_28_9,
  output [7:0]   io_tensor_rd_0_data_bits_28_10,
  output [7:0]   io_tensor_rd_0_data_bits_28_11,
  output [7:0]   io_tensor_rd_0_data_bits_28_12,
  output [7:0]   io_tensor_rd_0_data_bits_28_13,
  output [7:0]   io_tensor_rd_0_data_bits_28_14,
  output [7:0]   io_tensor_rd_0_data_bits_28_15,
  output [7:0]   io_tensor_rd_0_data_bits_29_0,
  output [7:0]   io_tensor_rd_0_data_bits_29_1,
  output [7:0]   io_tensor_rd_0_data_bits_29_2,
  output [7:0]   io_tensor_rd_0_data_bits_29_3,
  output [7:0]   io_tensor_rd_0_data_bits_29_4,
  output [7:0]   io_tensor_rd_0_data_bits_29_5,
  output [7:0]   io_tensor_rd_0_data_bits_29_6,
  output [7:0]   io_tensor_rd_0_data_bits_29_7,
  output [7:0]   io_tensor_rd_0_data_bits_29_8,
  output [7:0]   io_tensor_rd_0_data_bits_29_9,
  output [7:0]   io_tensor_rd_0_data_bits_29_10,
  output [7:0]   io_tensor_rd_0_data_bits_29_11,
  output [7:0]   io_tensor_rd_0_data_bits_29_12,
  output [7:0]   io_tensor_rd_0_data_bits_29_13,
  output [7:0]   io_tensor_rd_0_data_bits_29_14,
  output [7:0]   io_tensor_rd_0_data_bits_29_15,
  output [7:0]   io_tensor_rd_0_data_bits_30_0,
  output [7:0]   io_tensor_rd_0_data_bits_30_1,
  output [7:0]   io_tensor_rd_0_data_bits_30_2,
  output [7:0]   io_tensor_rd_0_data_bits_30_3,
  output [7:0]   io_tensor_rd_0_data_bits_30_4,
  output [7:0]   io_tensor_rd_0_data_bits_30_5,
  output [7:0]   io_tensor_rd_0_data_bits_30_6,
  output [7:0]   io_tensor_rd_0_data_bits_30_7,
  output [7:0]   io_tensor_rd_0_data_bits_30_8,
  output [7:0]   io_tensor_rd_0_data_bits_30_9,
  output [7:0]   io_tensor_rd_0_data_bits_30_10,
  output [7:0]   io_tensor_rd_0_data_bits_30_11,
  output [7:0]   io_tensor_rd_0_data_bits_30_12,
  output [7:0]   io_tensor_rd_0_data_bits_30_13,
  output [7:0]   io_tensor_rd_0_data_bits_30_14,
  output [7:0]   io_tensor_rd_0_data_bits_30_15,
  output [7:0]   io_tensor_rd_0_data_bits_31_0,
  output [7:0]   io_tensor_rd_0_data_bits_31_1,
  output [7:0]   io_tensor_rd_0_data_bits_31_2,
  output [7:0]   io_tensor_rd_0_data_bits_31_3,
  output [7:0]   io_tensor_rd_0_data_bits_31_4,
  output [7:0]   io_tensor_rd_0_data_bits_31_5,
  output [7:0]   io_tensor_rd_0_data_bits_31_6,
  output [7:0]   io_tensor_rd_0_data_bits_31_7,
  output [7:0]   io_tensor_rd_0_data_bits_31_8,
  output [7:0]   io_tensor_rd_0_data_bits_31_9,
  output [7:0]   io_tensor_rd_0_data_bits_31_10,
  output [7:0]   io_tensor_rd_0_data_bits_31_11,
  output [7:0]   io_tensor_rd_0_data_bits_31_12,
  output [7:0]   io_tensor_rd_0_data_bits_31_13,
  output [7:0]   io_tensor_rd_0_data_bits_31_14,
  output [7:0]   io_tensor_rd_0_data_bits_31_15
);
  wire  tensorLoad_clock; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_reset; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_start; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_done; // @[TensorLoad.scala 71:28]
  wire [127:0] tensorLoad_io_inst; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_baddr; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_vme_rd_cmd_ready; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_vme_rd_cmd_valid; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_vme_rd_cmd_bits_addr; // @[TensorLoad.scala 71:28]
  wire [3:0] tensorLoad_io_vme_rd_cmd_bits_len; // @[TensorLoad.scala 71:28]
  wire [20:0] tensorLoad_io_vme_rd_cmd_bits_tag; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_vme_rd_data_ready; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_vme_rd_data_valid; // @[TensorLoad.scala 71:28]
  wire [63:0] tensorLoad_io_vme_rd_data_bits_data; // @[TensorLoad.scala 71:28]
  wire [20:0] tensorLoad_io_vme_rd_data_bits_tag; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_tensor_rd_0_idx_valid; // @[TensorLoad.scala 71:28]
  wire [5:0] tensorLoad_io_tensor_rd_0_idx_bits; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_tensor_rd_0_data_valid; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_0_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_1_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_1_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_1_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_1_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_1_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_1_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_1_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_1_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_1_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_1_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_1_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_1_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_1_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_1_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_1_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_1_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_2_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_2_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_2_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_2_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_2_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_2_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_2_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_2_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_2_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_2_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_2_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_2_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_2_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_2_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_2_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_2_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_3_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_3_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_3_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_3_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_3_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_3_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_3_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_3_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_3_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_3_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_3_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_3_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_3_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_3_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_3_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_3_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_4_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_4_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_4_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_4_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_4_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_4_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_4_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_4_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_4_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_4_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_4_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_4_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_4_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_4_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_4_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_4_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_5_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_5_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_5_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_5_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_5_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_5_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_5_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_5_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_5_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_5_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_5_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_5_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_5_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_5_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_5_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_5_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_6_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_6_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_6_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_6_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_6_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_6_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_6_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_6_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_6_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_6_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_6_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_6_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_6_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_6_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_6_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_6_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_7_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_7_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_7_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_7_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_7_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_7_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_7_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_7_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_7_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_7_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_7_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_7_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_7_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_7_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_7_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_7_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_8_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_8_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_8_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_8_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_8_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_8_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_8_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_8_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_8_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_8_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_8_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_8_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_8_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_8_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_8_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_8_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_9_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_9_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_9_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_9_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_9_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_9_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_9_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_9_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_9_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_9_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_9_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_9_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_9_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_9_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_9_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_9_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_10_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_10_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_10_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_10_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_10_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_10_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_10_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_10_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_10_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_10_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_10_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_10_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_10_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_10_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_10_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_10_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_11_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_11_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_11_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_11_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_11_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_11_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_11_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_11_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_11_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_11_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_11_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_11_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_11_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_11_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_11_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_11_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_12_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_12_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_12_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_12_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_12_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_12_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_12_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_12_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_12_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_12_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_12_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_12_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_12_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_12_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_12_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_12_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_13_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_13_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_13_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_13_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_13_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_13_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_13_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_13_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_13_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_13_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_13_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_13_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_13_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_13_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_13_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_13_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_14_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_14_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_14_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_14_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_14_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_14_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_14_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_14_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_14_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_14_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_14_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_14_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_14_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_14_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_14_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_14_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_15_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_15_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_15_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_15_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_15_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_15_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_15_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_15_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_15_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_15_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_15_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_15_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_15_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_15_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_15_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_15_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_16_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_16_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_16_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_16_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_16_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_16_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_16_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_16_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_16_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_16_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_16_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_16_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_16_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_16_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_16_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_16_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_17_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_17_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_17_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_17_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_17_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_17_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_17_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_17_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_17_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_17_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_17_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_17_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_17_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_17_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_17_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_17_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_18_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_18_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_18_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_18_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_18_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_18_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_18_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_18_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_18_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_18_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_18_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_18_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_18_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_18_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_18_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_18_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_19_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_19_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_19_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_19_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_19_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_19_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_19_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_19_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_19_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_19_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_19_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_19_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_19_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_19_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_19_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_19_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_20_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_20_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_20_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_20_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_20_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_20_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_20_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_20_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_20_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_20_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_20_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_20_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_20_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_20_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_20_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_20_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_21_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_21_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_21_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_21_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_21_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_21_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_21_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_21_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_21_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_21_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_21_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_21_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_21_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_21_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_21_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_21_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_22_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_22_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_22_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_22_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_22_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_22_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_22_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_22_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_22_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_22_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_22_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_22_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_22_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_22_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_22_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_22_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_23_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_23_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_23_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_23_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_23_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_23_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_23_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_23_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_23_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_23_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_23_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_23_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_23_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_23_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_23_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_23_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_24_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_24_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_24_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_24_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_24_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_24_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_24_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_24_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_24_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_24_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_24_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_24_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_24_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_24_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_24_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_24_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_25_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_25_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_25_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_25_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_25_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_25_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_25_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_25_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_25_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_25_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_25_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_25_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_25_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_25_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_25_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_25_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_26_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_26_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_26_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_26_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_26_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_26_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_26_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_26_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_26_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_26_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_26_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_26_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_26_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_26_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_26_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_26_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_27_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_27_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_27_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_27_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_27_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_27_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_27_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_27_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_27_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_27_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_27_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_27_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_27_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_27_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_27_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_27_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_28_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_28_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_28_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_28_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_28_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_28_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_28_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_28_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_28_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_28_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_28_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_28_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_28_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_28_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_28_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_28_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_29_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_29_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_29_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_29_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_29_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_29_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_29_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_29_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_29_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_29_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_29_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_29_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_29_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_29_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_29_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_29_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_30_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_30_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_30_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_30_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_30_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_30_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_30_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_30_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_30_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_30_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_30_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_30_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_30_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_30_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_30_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_30_15; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_31_0; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_31_1; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_31_2; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_31_3; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_31_4; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_31_5; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_31_6; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_31_7; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_31_8; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_31_9; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_31_10; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_31_11; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_31_12; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_31_13; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_31_14; // @[TensorLoad.scala 71:28]
  wire [7:0] tensorLoad_io_tensor_rd_0_data_bits_31_15; // @[TensorLoad.scala 71:28]
  TensorLoadNarrowVME_1 tensorLoad ( // @[TensorLoad.scala 71:28]
    .clock(tensorLoad_clock),
    .reset(tensorLoad_reset),
    .io_start(tensorLoad_io_start),
    .io_done(tensorLoad_io_done),
    .io_inst(tensorLoad_io_inst),
    .io_baddr(tensorLoad_io_baddr),
    .io_vme_rd_cmd_ready(tensorLoad_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(tensorLoad_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(tensorLoad_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(tensorLoad_io_vme_rd_cmd_bits_len),
    .io_vme_rd_cmd_bits_tag(tensorLoad_io_vme_rd_cmd_bits_tag),
    .io_vme_rd_data_ready(tensorLoad_io_vme_rd_data_ready),
    .io_vme_rd_data_valid(tensorLoad_io_vme_rd_data_valid),
    .io_vme_rd_data_bits_data(tensorLoad_io_vme_rd_data_bits_data),
    .io_vme_rd_data_bits_tag(tensorLoad_io_vme_rd_data_bits_tag),
    .io_tensor_rd_0_idx_valid(tensorLoad_io_tensor_rd_0_idx_valid),
    .io_tensor_rd_0_idx_bits(tensorLoad_io_tensor_rd_0_idx_bits),
    .io_tensor_rd_0_data_valid(tensorLoad_io_tensor_rd_0_data_valid),
    .io_tensor_rd_0_data_bits_0_0(tensorLoad_io_tensor_rd_0_data_bits_0_0),
    .io_tensor_rd_0_data_bits_0_1(tensorLoad_io_tensor_rd_0_data_bits_0_1),
    .io_tensor_rd_0_data_bits_0_2(tensorLoad_io_tensor_rd_0_data_bits_0_2),
    .io_tensor_rd_0_data_bits_0_3(tensorLoad_io_tensor_rd_0_data_bits_0_3),
    .io_tensor_rd_0_data_bits_0_4(tensorLoad_io_tensor_rd_0_data_bits_0_4),
    .io_tensor_rd_0_data_bits_0_5(tensorLoad_io_tensor_rd_0_data_bits_0_5),
    .io_tensor_rd_0_data_bits_0_6(tensorLoad_io_tensor_rd_0_data_bits_0_6),
    .io_tensor_rd_0_data_bits_0_7(tensorLoad_io_tensor_rd_0_data_bits_0_7),
    .io_tensor_rd_0_data_bits_0_8(tensorLoad_io_tensor_rd_0_data_bits_0_8),
    .io_tensor_rd_0_data_bits_0_9(tensorLoad_io_tensor_rd_0_data_bits_0_9),
    .io_tensor_rd_0_data_bits_0_10(tensorLoad_io_tensor_rd_0_data_bits_0_10),
    .io_tensor_rd_0_data_bits_0_11(tensorLoad_io_tensor_rd_0_data_bits_0_11),
    .io_tensor_rd_0_data_bits_0_12(tensorLoad_io_tensor_rd_0_data_bits_0_12),
    .io_tensor_rd_0_data_bits_0_13(tensorLoad_io_tensor_rd_0_data_bits_0_13),
    .io_tensor_rd_0_data_bits_0_14(tensorLoad_io_tensor_rd_0_data_bits_0_14),
    .io_tensor_rd_0_data_bits_0_15(tensorLoad_io_tensor_rd_0_data_bits_0_15),
    .io_tensor_rd_0_data_bits_1_0(tensorLoad_io_tensor_rd_0_data_bits_1_0),
    .io_tensor_rd_0_data_bits_1_1(tensorLoad_io_tensor_rd_0_data_bits_1_1),
    .io_tensor_rd_0_data_bits_1_2(tensorLoad_io_tensor_rd_0_data_bits_1_2),
    .io_tensor_rd_0_data_bits_1_3(tensorLoad_io_tensor_rd_0_data_bits_1_3),
    .io_tensor_rd_0_data_bits_1_4(tensorLoad_io_tensor_rd_0_data_bits_1_4),
    .io_tensor_rd_0_data_bits_1_5(tensorLoad_io_tensor_rd_0_data_bits_1_5),
    .io_tensor_rd_0_data_bits_1_6(tensorLoad_io_tensor_rd_0_data_bits_1_6),
    .io_tensor_rd_0_data_bits_1_7(tensorLoad_io_tensor_rd_0_data_bits_1_7),
    .io_tensor_rd_0_data_bits_1_8(tensorLoad_io_tensor_rd_0_data_bits_1_8),
    .io_tensor_rd_0_data_bits_1_9(tensorLoad_io_tensor_rd_0_data_bits_1_9),
    .io_tensor_rd_0_data_bits_1_10(tensorLoad_io_tensor_rd_0_data_bits_1_10),
    .io_tensor_rd_0_data_bits_1_11(tensorLoad_io_tensor_rd_0_data_bits_1_11),
    .io_tensor_rd_0_data_bits_1_12(tensorLoad_io_tensor_rd_0_data_bits_1_12),
    .io_tensor_rd_0_data_bits_1_13(tensorLoad_io_tensor_rd_0_data_bits_1_13),
    .io_tensor_rd_0_data_bits_1_14(tensorLoad_io_tensor_rd_0_data_bits_1_14),
    .io_tensor_rd_0_data_bits_1_15(tensorLoad_io_tensor_rd_0_data_bits_1_15),
    .io_tensor_rd_0_data_bits_2_0(tensorLoad_io_tensor_rd_0_data_bits_2_0),
    .io_tensor_rd_0_data_bits_2_1(tensorLoad_io_tensor_rd_0_data_bits_2_1),
    .io_tensor_rd_0_data_bits_2_2(tensorLoad_io_tensor_rd_0_data_bits_2_2),
    .io_tensor_rd_0_data_bits_2_3(tensorLoad_io_tensor_rd_0_data_bits_2_3),
    .io_tensor_rd_0_data_bits_2_4(tensorLoad_io_tensor_rd_0_data_bits_2_4),
    .io_tensor_rd_0_data_bits_2_5(tensorLoad_io_tensor_rd_0_data_bits_2_5),
    .io_tensor_rd_0_data_bits_2_6(tensorLoad_io_tensor_rd_0_data_bits_2_6),
    .io_tensor_rd_0_data_bits_2_7(tensorLoad_io_tensor_rd_0_data_bits_2_7),
    .io_tensor_rd_0_data_bits_2_8(tensorLoad_io_tensor_rd_0_data_bits_2_8),
    .io_tensor_rd_0_data_bits_2_9(tensorLoad_io_tensor_rd_0_data_bits_2_9),
    .io_tensor_rd_0_data_bits_2_10(tensorLoad_io_tensor_rd_0_data_bits_2_10),
    .io_tensor_rd_0_data_bits_2_11(tensorLoad_io_tensor_rd_0_data_bits_2_11),
    .io_tensor_rd_0_data_bits_2_12(tensorLoad_io_tensor_rd_0_data_bits_2_12),
    .io_tensor_rd_0_data_bits_2_13(tensorLoad_io_tensor_rd_0_data_bits_2_13),
    .io_tensor_rd_0_data_bits_2_14(tensorLoad_io_tensor_rd_0_data_bits_2_14),
    .io_tensor_rd_0_data_bits_2_15(tensorLoad_io_tensor_rd_0_data_bits_2_15),
    .io_tensor_rd_0_data_bits_3_0(tensorLoad_io_tensor_rd_0_data_bits_3_0),
    .io_tensor_rd_0_data_bits_3_1(tensorLoad_io_tensor_rd_0_data_bits_3_1),
    .io_tensor_rd_0_data_bits_3_2(tensorLoad_io_tensor_rd_0_data_bits_3_2),
    .io_tensor_rd_0_data_bits_3_3(tensorLoad_io_tensor_rd_0_data_bits_3_3),
    .io_tensor_rd_0_data_bits_3_4(tensorLoad_io_tensor_rd_0_data_bits_3_4),
    .io_tensor_rd_0_data_bits_3_5(tensorLoad_io_tensor_rd_0_data_bits_3_5),
    .io_tensor_rd_0_data_bits_3_6(tensorLoad_io_tensor_rd_0_data_bits_3_6),
    .io_tensor_rd_0_data_bits_3_7(tensorLoad_io_tensor_rd_0_data_bits_3_7),
    .io_tensor_rd_0_data_bits_3_8(tensorLoad_io_tensor_rd_0_data_bits_3_8),
    .io_tensor_rd_0_data_bits_3_9(tensorLoad_io_tensor_rd_0_data_bits_3_9),
    .io_tensor_rd_0_data_bits_3_10(tensorLoad_io_tensor_rd_0_data_bits_3_10),
    .io_tensor_rd_0_data_bits_3_11(tensorLoad_io_tensor_rd_0_data_bits_3_11),
    .io_tensor_rd_0_data_bits_3_12(tensorLoad_io_tensor_rd_0_data_bits_3_12),
    .io_tensor_rd_0_data_bits_3_13(tensorLoad_io_tensor_rd_0_data_bits_3_13),
    .io_tensor_rd_0_data_bits_3_14(tensorLoad_io_tensor_rd_0_data_bits_3_14),
    .io_tensor_rd_0_data_bits_3_15(tensorLoad_io_tensor_rd_0_data_bits_3_15),
    .io_tensor_rd_0_data_bits_4_0(tensorLoad_io_tensor_rd_0_data_bits_4_0),
    .io_tensor_rd_0_data_bits_4_1(tensorLoad_io_tensor_rd_0_data_bits_4_1),
    .io_tensor_rd_0_data_bits_4_2(tensorLoad_io_tensor_rd_0_data_bits_4_2),
    .io_tensor_rd_0_data_bits_4_3(tensorLoad_io_tensor_rd_0_data_bits_4_3),
    .io_tensor_rd_0_data_bits_4_4(tensorLoad_io_tensor_rd_0_data_bits_4_4),
    .io_tensor_rd_0_data_bits_4_5(tensorLoad_io_tensor_rd_0_data_bits_4_5),
    .io_tensor_rd_0_data_bits_4_6(tensorLoad_io_tensor_rd_0_data_bits_4_6),
    .io_tensor_rd_0_data_bits_4_7(tensorLoad_io_tensor_rd_0_data_bits_4_7),
    .io_tensor_rd_0_data_bits_4_8(tensorLoad_io_tensor_rd_0_data_bits_4_8),
    .io_tensor_rd_0_data_bits_4_9(tensorLoad_io_tensor_rd_0_data_bits_4_9),
    .io_tensor_rd_0_data_bits_4_10(tensorLoad_io_tensor_rd_0_data_bits_4_10),
    .io_tensor_rd_0_data_bits_4_11(tensorLoad_io_tensor_rd_0_data_bits_4_11),
    .io_tensor_rd_0_data_bits_4_12(tensorLoad_io_tensor_rd_0_data_bits_4_12),
    .io_tensor_rd_0_data_bits_4_13(tensorLoad_io_tensor_rd_0_data_bits_4_13),
    .io_tensor_rd_0_data_bits_4_14(tensorLoad_io_tensor_rd_0_data_bits_4_14),
    .io_tensor_rd_0_data_bits_4_15(tensorLoad_io_tensor_rd_0_data_bits_4_15),
    .io_tensor_rd_0_data_bits_5_0(tensorLoad_io_tensor_rd_0_data_bits_5_0),
    .io_tensor_rd_0_data_bits_5_1(tensorLoad_io_tensor_rd_0_data_bits_5_1),
    .io_tensor_rd_0_data_bits_5_2(tensorLoad_io_tensor_rd_0_data_bits_5_2),
    .io_tensor_rd_0_data_bits_5_3(tensorLoad_io_tensor_rd_0_data_bits_5_3),
    .io_tensor_rd_0_data_bits_5_4(tensorLoad_io_tensor_rd_0_data_bits_5_4),
    .io_tensor_rd_0_data_bits_5_5(tensorLoad_io_tensor_rd_0_data_bits_5_5),
    .io_tensor_rd_0_data_bits_5_6(tensorLoad_io_tensor_rd_0_data_bits_5_6),
    .io_tensor_rd_0_data_bits_5_7(tensorLoad_io_tensor_rd_0_data_bits_5_7),
    .io_tensor_rd_0_data_bits_5_8(tensorLoad_io_tensor_rd_0_data_bits_5_8),
    .io_tensor_rd_0_data_bits_5_9(tensorLoad_io_tensor_rd_0_data_bits_5_9),
    .io_tensor_rd_0_data_bits_5_10(tensorLoad_io_tensor_rd_0_data_bits_5_10),
    .io_tensor_rd_0_data_bits_5_11(tensorLoad_io_tensor_rd_0_data_bits_5_11),
    .io_tensor_rd_0_data_bits_5_12(tensorLoad_io_tensor_rd_0_data_bits_5_12),
    .io_tensor_rd_0_data_bits_5_13(tensorLoad_io_tensor_rd_0_data_bits_5_13),
    .io_tensor_rd_0_data_bits_5_14(tensorLoad_io_tensor_rd_0_data_bits_5_14),
    .io_tensor_rd_0_data_bits_5_15(tensorLoad_io_tensor_rd_0_data_bits_5_15),
    .io_tensor_rd_0_data_bits_6_0(tensorLoad_io_tensor_rd_0_data_bits_6_0),
    .io_tensor_rd_0_data_bits_6_1(tensorLoad_io_tensor_rd_0_data_bits_6_1),
    .io_tensor_rd_0_data_bits_6_2(tensorLoad_io_tensor_rd_0_data_bits_6_2),
    .io_tensor_rd_0_data_bits_6_3(tensorLoad_io_tensor_rd_0_data_bits_6_3),
    .io_tensor_rd_0_data_bits_6_4(tensorLoad_io_tensor_rd_0_data_bits_6_4),
    .io_tensor_rd_0_data_bits_6_5(tensorLoad_io_tensor_rd_0_data_bits_6_5),
    .io_tensor_rd_0_data_bits_6_6(tensorLoad_io_tensor_rd_0_data_bits_6_6),
    .io_tensor_rd_0_data_bits_6_7(tensorLoad_io_tensor_rd_0_data_bits_6_7),
    .io_tensor_rd_0_data_bits_6_8(tensorLoad_io_tensor_rd_0_data_bits_6_8),
    .io_tensor_rd_0_data_bits_6_9(tensorLoad_io_tensor_rd_0_data_bits_6_9),
    .io_tensor_rd_0_data_bits_6_10(tensorLoad_io_tensor_rd_0_data_bits_6_10),
    .io_tensor_rd_0_data_bits_6_11(tensorLoad_io_tensor_rd_0_data_bits_6_11),
    .io_tensor_rd_0_data_bits_6_12(tensorLoad_io_tensor_rd_0_data_bits_6_12),
    .io_tensor_rd_0_data_bits_6_13(tensorLoad_io_tensor_rd_0_data_bits_6_13),
    .io_tensor_rd_0_data_bits_6_14(tensorLoad_io_tensor_rd_0_data_bits_6_14),
    .io_tensor_rd_0_data_bits_6_15(tensorLoad_io_tensor_rd_0_data_bits_6_15),
    .io_tensor_rd_0_data_bits_7_0(tensorLoad_io_tensor_rd_0_data_bits_7_0),
    .io_tensor_rd_0_data_bits_7_1(tensorLoad_io_tensor_rd_0_data_bits_7_1),
    .io_tensor_rd_0_data_bits_7_2(tensorLoad_io_tensor_rd_0_data_bits_7_2),
    .io_tensor_rd_0_data_bits_7_3(tensorLoad_io_tensor_rd_0_data_bits_7_3),
    .io_tensor_rd_0_data_bits_7_4(tensorLoad_io_tensor_rd_0_data_bits_7_4),
    .io_tensor_rd_0_data_bits_7_5(tensorLoad_io_tensor_rd_0_data_bits_7_5),
    .io_tensor_rd_0_data_bits_7_6(tensorLoad_io_tensor_rd_0_data_bits_7_6),
    .io_tensor_rd_0_data_bits_7_7(tensorLoad_io_tensor_rd_0_data_bits_7_7),
    .io_tensor_rd_0_data_bits_7_8(tensorLoad_io_tensor_rd_0_data_bits_7_8),
    .io_tensor_rd_0_data_bits_7_9(tensorLoad_io_tensor_rd_0_data_bits_7_9),
    .io_tensor_rd_0_data_bits_7_10(tensorLoad_io_tensor_rd_0_data_bits_7_10),
    .io_tensor_rd_0_data_bits_7_11(tensorLoad_io_tensor_rd_0_data_bits_7_11),
    .io_tensor_rd_0_data_bits_7_12(tensorLoad_io_tensor_rd_0_data_bits_7_12),
    .io_tensor_rd_0_data_bits_7_13(tensorLoad_io_tensor_rd_0_data_bits_7_13),
    .io_tensor_rd_0_data_bits_7_14(tensorLoad_io_tensor_rd_0_data_bits_7_14),
    .io_tensor_rd_0_data_bits_7_15(tensorLoad_io_tensor_rd_0_data_bits_7_15),
    .io_tensor_rd_0_data_bits_8_0(tensorLoad_io_tensor_rd_0_data_bits_8_0),
    .io_tensor_rd_0_data_bits_8_1(tensorLoad_io_tensor_rd_0_data_bits_8_1),
    .io_tensor_rd_0_data_bits_8_2(tensorLoad_io_tensor_rd_0_data_bits_8_2),
    .io_tensor_rd_0_data_bits_8_3(tensorLoad_io_tensor_rd_0_data_bits_8_3),
    .io_tensor_rd_0_data_bits_8_4(tensorLoad_io_tensor_rd_0_data_bits_8_4),
    .io_tensor_rd_0_data_bits_8_5(tensorLoad_io_tensor_rd_0_data_bits_8_5),
    .io_tensor_rd_0_data_bits_8_6(tensorLoad_io_tensor_rd_0_data_bits_8_6),
    .io_tensor_rd_0_data_bits_8_7(tensorLoad_io_tensor_rd_0_data_bits_8_7),
    .io_tensor_rd_0_data_bits_8_8(tensorLoad_io_tensor_rd_0_data_bits_8_8),
    .io_tensor_rd_0_data_bits_8_9(tensorLoad_io_tensor_rd_0_data_bits_8_9),
    .io_tensor_rd_0_data_bits_8_10(tensorLoad_io_tensor_rd_0_data_bits_8_10),
    .io_tensor_rd_0_data_bits_8_11(tensorLoad_io_tensor_rd_0_data_bits_8_11),
    .io_tensor_rd_0_data_bits_8_12(tensorLoad_io_tensor_rd_0_data_bits_8_12),
    .io_tensor_rd_0_data_bits_8_13(tensorLoad_io_tensor_rd_0_data_bits_8_13),
    .io_tensor_rd_0_data_bits_8_14(tensorLoad_io_tensor_rd_0_data_bits_8_14),
    .io_tensor_rd_0_data_bits_8_15(tensorLoad_io_tensor_rd_0_data_bits_8_15),
    .io_tensor_rd_0_data_bits_9_0(tensorLoad_io_tensor_rd_0_data_bits_9_0),
    .io_tensor_rd_0_data_bits_9_1(tensorLoad_io_tensor_rd_0_data_bits_9_1),
    .io_tensor_rd_0_data_bits_9_2(tensorLoad_io_tensor_rd_0_data_bits_9_2),
    .io_tensor_rd_0_data_bits_9_3(tensorLoad_io_tensor_rd_0_data_bits_9_3),
    .io_tensor_rd_0_data_bits_9_4(tensorLoad_io_tensor_rd_0_data_bits_9_4),
    .io_tensor_rd_0_data_bits_9_5(tensorLoad_io_tensor_rd_0_data_bits_9_5),
    .io_tensor_rd_0_data_bits_9_6(tensorLoad_io_tensor_rd_0_data_bits_9_6),
    .io_tensor_rd_0_data_bits_9_7(tensorLoad_io_tensor_rd_0_data_bits_9_7),
    .io_tensor_rd_0_data_bits_9_8(tensorLoad_io_tensor_rd_0_data_bits_9_8),
    .io_tensor_rd_0_data_bits_9_9(tensorLoad_io_tensor_rd_0_data_bits_9_9),
    .io_tensor_rd_0_data_bits_9_10(tensorLoad_io_tensor_rd_0_data_bits_9_10),
    .io_tensor_rd_0_data_bits_9_11(tensorLoad_io_tensor_rd_0_data_bits_9_11),
    .io_tensor_rd_0_data_bits_9_12(tensorLoad_io_tensor_rd_0_data_bits_9_12),
    .io_tensor_rd_0_data_bits_9_13(tensorLoad_io_tensor_rd_0_data_bits_9_13),
    .io_tensor_rd_0_data_bits_9_14(tensorLoad_io_tensor_rd_0_data_bits_9_14),
    .io_tensor_rd_0_data_bits_9_15(tensorLoad_io_tensor_rd_0_data_bits_9_15),
    .io_tensor_rd_0_data_bits_10_0(tensorLoad_io_tensor_rd_0_data_bits_10_0),
    .io_tensor_rd_0_data_bits_10_1(tensorLoad_io_tensor_rd_0_data_bits_10_1),
    .io_tensor_rd_0_data_bits_10_2(tensorLoad_io_tensor_rd_0_data_bits_10_2),
    .io_tensor_rd_0_data_bits_10_3(tensorLoad_io_tensor_rd_0_data_bits_10_3),
    .io_tensor_rd_0_data_bits_10_4(tensorLoad_io_tensor_rd_0_data_bits_10_4),
    .io_tensor_rd_0_data_bits_10_5(tensorLoad_io_tensor_rd_0_data_bits_10_5),
    .io_tensor_rd_0_data_bits_10_6(tensorLoad_io_tensor_rd_0_data_bits_10_6),
    .io_tensor_rd_0_data_bits_10_7(tensorLoad_io_tensor_rd_0_data_bits_10_7),
    .io_tensor_rd_0_data_bits_10_8(tensorLoad_io_tensor_rd_0_data_bits_10_8),
    .io_tensor_rd_0_data_bits_10_9(tensorLoad_io_tensor_rd_0_data_bits_10_9),
    .io_tensor_rd_0_data_bits_10_10(tensorLoad_io_tensor_rd_0_data_bits_10_10),
    .io_tensor_rd_0_data_bits_10_11(tensorLoad_io_tensor_rd_0_data_bits_10_11),
    .io_tensor_rd_0_data_bits_10_12(tensorLoad_io_tensor_rd_0_data_bits_10_12),
    .io_tensor_rd_0_data_bits_10_13(tensorLoad_io_tensor_rd_0_data_bits_10_13),
    .io_tensor_rd_0_data_bits_10_14(tensorLoad_io_tensor_rd_0_data_bits_10_14),
    .io_tensor_rd_0_data_bits_10_15(tensorLoad_io_tensor_rd_0_data_bits_10_15),
    .io_tensor_rd_0_data_bits_11_0(tensorLoad_io_tensor_rd_0_data_bits_11_0),
    .io_tensor_rd_0_data_bits_11_1(tensorLoad_io_tensor_rd_0_data_bits_11_1),
    .io_tensor_rd_0_data_bits_11_2(tensorLoad_io_tensor_rd_0_data_bits_11_2),
    .io_tensor_rd_0_data_bits_11_3(tensorLoad_io_tensor_rd_0_data_bits_11_3),
    .io_tensor_rd_0_data_bits_11_4(tensorLoad_io_tensor_rd_0_data_bits_11_4),
    .io_tensor_rd_0_data_bits_11_5(tensorLoad_io_tensor_rd_0_data_bits_11_5),
    .io_tensor_rd_0_data_bits_11_6(tensorLoad_io_tensor_rd_0_data_bits_11_6),
    .io_tensor_rd_0_data_bits_11_7(tensorLoad_io_tensor_rd_0_data_bits_11_7),
    .io_tensor_rd_0_data_bits_11_8(tensorLoad_io_tensor_rd_0_data_bits_11_8),
    .io_tensor_rd_0_data_bits_11_9(tensorLoad_io_tensor_rd_0_data_bits_11_9),
    .io_tensor_rd_0_data_bits_11_10(tensorLoad_io_tensor_rd_0_data_bits_11_10),
    .io_tensor_rd_0_data_bits_11_11(tensorLoad_io_tensor_rd_0_data_bits_11_11),
    .io_tensor_rd_0_data_bits_11_12(tensorLoad_io_tensor_rd_0_data_bits_11_12),
    .io_tensor_rd_0_data_bits_11_13(tensorLoad_io_tensor_rd_0_data_bits_11_13),
    .io_tensor_rd_0_data_bits_11_14(tensorLoad_io_tensor_rd_0_data_bits_11_14),
    .io_tensor_rd_0_data_bits_11_15(tensorLoad_io_tensor_rd_0_data_bits_11_15),
    .io_tensor_rd_0_data_bits_12_0(tensorLoad_io_tensor_rd_0_data_bits_12_0),
    .io_tensor_rd_0_data_bits_12_1(tensorLoad_io_tensor_rd_0_data_bits_12_1),
    .io_tensor_rd_0_data_bits_12_2(tensorLoad_io_tensor_rd_0_data_bits_12_2),
    .io_tensor_rd_0_data_bits_12_3(tensorLoad_io_tensor_rd_0_data_bits_12_3),
    .io_tensor_rd_0_data_bits_12_4(tensorLoad_io_tensor_rd_0_data_bits_12_4),
    .io_tensor_rd_0_data_bits_12_5(tensorLoad_io_tensor_rd_0_data_bits_12_5),
    .io_tensor_rd_0_data_bits_12_6(tensorLoad_io_tensor_rd_0_data_bits_12_6),
    .io_tensor_rd_0_data_bits_12_7(tensorLoad_io_tensor_rd_0_data_bits_12_7),
    .io_tensor_rd_0_data_bits_12_8(tensorLoad_io_tensor_rd_0_data_bits_12_8),
    .io_tensor_rd_0_data_bits_12_9(tensorLoad_io_tensor_rd_0_data_bits_12_9),
    .io_tensor_rd_0_data_bits_12_10(tensorLoad_io_tensor_rd_0_data_bits_12_10),
    .io_tensor_rd_0_data_bits_12_11(tensorLoad_io_tensor_rd_0_data_bits_12_11),
    .io_tensor_rd_0_data_bits_12_12(tensorLoad_io_tensor_rd_0_data_bits_12_12),
    .io_tensor_rd_0_data_bits_12_13(tensorLoad_io_tensor_rd_0_data_bits_12_13),
    .io_tensor_rd_0_data_bits_12_14(tensorLoad_io_tensor_rd_0_data_bits_12_14),
    .io_tensor_rd_0_data_bits_12_15(tensorLoad_io_tensor_rd_0_data_bits_12_15),
    .io_tensor_rd_0_data_bits_13_0(tensorLoad_io_tensor_rd_0_data_bits_13_0),
    .io_tensor_rd_0_data_bits_13_1(tensorLoad_io_tensor_rd_0_data_bits_13_1),
    .io_tensor_rd_0_data_bits_13_2(tensorLoad_io_tensor_rd_0_data_bits_13_2),
    .io_tensor_rd_0_data_bits_13_3(tensorLoad_io_tensor_rd_0_data_bits_13_3),
    .io_tensor_rd_0_data_bits_13_4(tensorLoad_io_tensor_rd_0_data_bits_13_4),
    .io_tensor_rd_0_data_bits_13_5(tensorLoad_io_tensor_rd_0_data_bits_13_5),
    .io_tensor_rd_0_data_bits_13_6(tensorLoad_io_tensor_rd_0_data_bits_13_6),
    .io_tensor_rd_0_data_bits_13_7(tensorLoad_io_tensor_rd_0_data_bits_13_7),
    .io_tensor_rd_0_data_bits_13_8(tensorLoad_io_tensor_rd_0_data_bits_13_8),
    .io_tensor_rd_0_data_bits_13_9(tensorLoad_io_tensor_rd_0_data_bits_13_9),
    .io_tensor_rd_0_data_bits_13_10(tensorLoad_io_tensor_rd_0_data_bits_13_10),
    .io_tensor_rd_0_data_bits_13_11(tensorLoad_io_tensor_rd_0_data_bits_13_11),
    .io_tensor_rd_0_data_bits_13_12(tensorLoad_io_tensor_rd_0_data_bits_13_12),
    .io_tensor_rd_0_data_bits_13_13(tensorLoad_io_tensor_rd_0_data_bits_13_13),
    .io_tensor_rd_0_data_bits_13_14(tensorLoad_io_tensor_rd_0_data_bits_13_14),
    .io_tensor_rd_0_data_bits_13_15(tensorLoad_io_tensor_rd_0_data_bits_13_15),
    .io_tensor_rd_0_data_bits_14_0(tensorLoad_io_tensor_rd_0_data_bits_14_0),
    .io_tensor_rd_0_data_bits_14_1(tensorLoad_io_tensor_rd_0_data_bits_14_1),
    .io_tensor_rd_0_data_bits_14_2(tensorLoad_io_tensor_rd_0_data_bits_14_2),
    .io_tensor_rd_0_data_bits_14_3(tensorLoad_io_tensor_rd_0_data_bits_14_3),
    .io_tensor_rd_0_data_bits_14_4(tensorLoad_io_tensor_rd_0_data_bits_14_4),
    .io_tensor_rd_0_data_bits_14_5(tensorLoad_io_tensor_rd_0_data_bits_14_5),
    .io_tensor_rd_0_data_bits_14_6(tensorLoad_io_tensor_rd_0_data_bits_14_6),
    .io_tensor_rd_0_data_bits_14_7(tensorLoad_io_tensor_rd_0_data_bits_14_7),
    .io_tensor_rd_0_data_bits_14_8(tensorLoad_io_tensor_rd_0_data_bits_14_8),
    .io_tensor_rd_0_data_bits_14_9(tensorLoad_io_tensor_rd_0_data_bits_14_9),
    .io_tensor_rd_0_data_bits_14_10(tensorLoad_io_tensor_rd_0_data_bits_14_10),
    .io_tensor_rd_0_data_bits_14_11(tensorLoad_io_tensor_rd_0_data_bits_14_11),
    .io_tensor_rd_0_data_bits_14_12(tensorLoad_io_tensor_rd_0_data_bits_14_12),
    .io_tensor_rd_0_data_bits_14_13(tensorLoad_io_tensor_rd_0_data_bits_14_13),
    .io_tensor_rd_0_data_bits_14_14(tensorLoad_io_tensor_rd_0_data_bits_14_14),
    .io_tensor_rd_0_data_bits_14_15(tensorLoad_io_tensor_rd_0_data_bits_14_15),
    .io_tensor_rd_0_data_bits_15_0(tensorLoad_io_tensor_rd_0_data_bits_15_0),
    .io_tensor_rd_0_data_bits_15_1(tensorLoad_io_tensor_rd_0_data_bits_15_1),
    .io_tensor_rd_0_data_bits_15_2(tensorLoad_io_tensor_rd_0_data_bits_15_2),
    .io_tensor_rd_0_data_bits_15_3(tensorLoad_io_tensor_rd_0_data_bits_15_3),
    .io_tensor_rd_0_data_bits_15_4(tensorLoad_io_tensor_rd_0_data_bits_15_4),
    .io_tensor_rd_0_data_bits_15_5(tensorLoad_io_tensor_rd_0_data_bits_15_5),
    .io_tensor_rd_0_data_bits_15_6(tensorLoad_io_tensor_rd_0_data_bits_15_6),
    .io_tensor_rd_0_data_bits_15_7(tensorLoad_io_tensor_rd_0_data_bits_15_7),
    .io_tensor_rd_0_data_bits_15_8(tensorLoad_io_tensor_rd_0_data_bits_15_8),
    .io_tensor_rd_0_data_bits_15_9(tensorLoad_io_tensor_rd_0_data_bits_15_9),
    .io_tensor_rd_0_data_bits_15_10(tensorLoad_io_tensor_rd_0_data_bits_15_10),
    .io_tensor_rd_0_data_bits_15_11(tensorLoad_io_tensor_rd_0_data_bits_15_11),
    .io_tensor_rd_0_data_bits_15_12(tensorLoad_io_tensor_rd_0_data_bits_15_12),
    .io_tensor_rd_0_data_bits_15_13(tensorLoad_io_tensor_rd_0_data_bits_15_13),
    .io_tensor_rd_0_data_bits_15_14(tensorLoad_io_tensor_rd_0_data_bits_15_14),
    .io_tensor_rd_0_data_bits_15_15(tensorLoad_io_tensor_rd_0_data_bits_15_15),
    .io_tensor_rd_0_data_bits_16_0(tensorLoad_io_tensor_rd_0_data_bits_16_0),
    .io_tensor_rd_0_data_bits_16_1(tensorLoad_io_tensor_rd_0_data_bits_16_1),
    .io_tensor_rd_0_data_bits_16_2(tensorLoad_io_tensor_rd_0_data_bits_16_2),
    .io_tensor_rd_0_data_bits_16_3(tensorLoad_io_tensor_rd_0_data_bits_16_3),
    .io_tensor_rd_0_data_bits_16_4(tensorLoad_io_tensor_rd_0_data_bits_16_4),
    .io_tensor_rd_0_data_bits_16_5(tensorLoad_io_tensor_rd_0_data_bits_16_5),
    .io_tensor_rd_0_data_bits_16_6(tensorLoad_io_tensor_rd_0_data_bits_16_6),
    .io_tensor_rd_0_data_bits_16_7(tensorLoad_io_tensor_rd_0_data_bits_16_7),
    .io_tensor_rd_0_data_bits_16_8(tensorLoad_io_tensor_rd_0_data_bits_16_8),
    .io_tensor_rd_0_data_bits_16_9(tensorLoad_io_tensor_rd_0_data_bits_16_9),
    .io_tensor_rd_0_data_bits_16_10(tensorLoad_io_tensor_rd_0_data_bits_16_10),
    .io_tensor_rd_0_data_bits_16_11(tensorLoad_io_tensor_rd_0_data_bits_16_11),
    .io_tensor_rd_0_data_bits_16_12(tensorLoad_io_tensor_rd_0_data_bits_16_12),
    .io_tensor_rd_0_data_bits_16_13(tensorLoad_io_tensor_rd_0_data_bits_16_13),
    .io_tensor_rd_0_data_bits_16_14(tensorLoad_io_tensor_rd_0_data_bits_16_14),
    .io_tensor_rd_0_data_bits_16_15(tensorLoad_io_tensor_rd_0_data_bits_16_15),
    .io_tensor_rd_0_data_bits_17_0(tensorLoad_io_tensor_rd_0_data_bits_17_0),
    .io_tensor_rd_0_data_bits_17_1(tensorLoad_io_tensor_rd_0_data_bits_17_1),
    .io_tensor_rd_0_data_bits_17_2(tensorLoad_io_tensor_rd_0_data_bits_17_2),
    .io_tensor_rd_0_data_bits_17_3(tensorLoad_io_tensor_rd_0_data_bits_17_3),
    .io_tensor_rd_0_data_bits_17_4(tensorLoad_io_tensor_rd_0_data_bits_17_4),
    .io_tensor_rd_0_data_bits_17_5(tensorLoad_io_tensor_rd_0_data_bits_17_5),
    .io_tensor_rd_0_data_bits_17_6(tensorLoad_io_tensor_rd_0_data_bits_17_6),
    .io_tensor_rd_0_data_bits_17_7(tensorLoad_io_tensor_rd_0_data_bits_17_7),
    .io_tensor_rd_0_data_bits_17_8(tensorLoad_io_tensor_rd_0_data_bits_17_8),
    .io_tensor_rd_0_data_bits_17_9(tensorLoad_io_tensor_rd_0_data_bits_17_9),
    .io_tensor_rd_0_data_bits_17_10(tensorLoad_io_tensor_rd_0_data_bits_17_10),
    .io_tensor_rd_0_data_bits_17_11(tensorLoad_io_tensor_rd_0_data_bits_17_11),
    .io_tensor_rd_0_data_bits_17_12(tensorLoad_io_tensor_rd_0_data_bits_17_12),
    .io_tensor_rd_0_data_bits_17_13(tensorLoad_io_tensor_rd_0_data_bits_17_13),
    .io_tensor_rd_0_data_bits_17_14(tensorLoad_io_tensor_rd_0_data_bits_17_14),
    .io_tensor_rd_0_data_bits_17_15(tensorLoad_io_tensor_rd_0_data_bits_17_15),
    .io_tensor_rd_0_data_bits_18_0(tensorLoad_io_tensor_rd_0_data_bits_18_0),
    .io_tensor_rd_0_data_bits_18_1(tensorLoad_io_tensor_rd_0_data_bits_18_1),
    .io_tensor_rd_0_data_bits_18_2(tensorLoad_io_tensor_rd_0_data_bits_18_2),
    .io_tensor_rd_0_data_bits_18_3(tensorLoad_io_tensor_rd_0_data_bits_18_3),
    .io_tensor_rd_0_data_bits_18_4(tensorLoad_io_tensor_rd_0_data_bits_18_4),
    .io_tensor_rd_0_data_bits_18_5(tensorLoad_io_tensor_rd_0_data_bits_18_5),
    .io_tensor_rd_0_data_bits_18_6(tensorLoad_io_tensor_rd_0_data_bits_18_6),
    .io_tensor_rd_0_data_bits_18_7(tensorLoad_io_tensor_rd_0_data_bits_18_7),
    .io_tensor_rd_0_data_bits_18_8(tensorLoad_io_tensor_rd_0_data_bits_18_8),
    .io_tensor_rd_0_data_bits_18_9(tensorLoad_io_tensor_rd_0_data_bits_18_9),
    .io_tensor_rd_0_data_bits_18_10(tensorLoad_io_tensor_rd_0_data_bits_18_10),
    .io_tensor_rd_0_data_bits_18_11(tensorLoad_io_tensor_rd_0_data_bits_18_11),
    .io_tensor_rd_0_data_bits_18_12(tensorLoad_io_tensor_rd_0_data_bits_18_12),
    .io_tensor_rd_0_data_bits_18_13(tensorLoad_io_tensor_rd_0_data_bits_18_13),
    .io_tensor_rd_0_data_bits_18_14(tensorLoad_io_tensor_rd_0_data_bits_18_14),
    .io_tensor_rd_0_data_bits_18_15(tensorLoad_io_tensor_rd_0_data_bits_18_15),
    .io_tensor_rd_0_data_bits_19_0(tensorLoad_io_tensor_rd_0_data_bits_19_0),
    .io_tensor_rd_0_data_bits_19_1(tensorLoad_io_tensor_rd_0_data_bits_19_1),
    .io_tensor_rd_0_data_bits_19_2(tensorLoad_io_tensor_rd_0_data_bits_19_2),
    .io_tensor_rd_0_data_bits_19_3(tensorLoad_io_tensor_rd_0_data_bits_19_3),
    .io_tensor_rd_0_data_bits_19_4(tensorLoad_io_tensor_rd_0_data_bits_19_4),
    .io_tensor_rd_0_data_bits_19_5(tensorLoad_io_tensor_rd_0_data_bits_19_5),
    .io_tensor_rd_0_data_bits_19_6(tensorLoad_io_tensor_rd_0_data_bits_19_6),
    .io_tensor_rd_0_data_bits_19_7(tensorLoad_io_tensor_rd_0_data_bits_19_7),
    .io_tensor_rd_0_data_bits_19_8(tensorLoad_io_tensor_rd_0_data_bits_19_8),
    .io_tensor_rd_0_data_bits_19_9(tensorLoad_io_tensor_rd_0_data_bits_19_9),
    .io_tensor_rd_0_data_bits_19_10(tensorLoad_io_tensor_rd_0_data_bits_19_10),
    .io_tensor_rd_0_data_bits_19_11(tensorLoad_io_tensor_rd_0_data_bits_19_11),
    .io_tensor_rd_0_data_bits_19_12(tensorLoad_io_tensor_rd_0_data_bits_19_12),
    .io_tensor_rd_0_data_bits_19_13(tensorLoad_io_tensor_rd_0_data_bits_19_13),
    .io_tensor_rd_0_data_bits_19_14(tensorLoad_io_tensor_rd_0_data_bits_19_14),
    .io_tensor_rd_0_data_bits_19_15(tensorLoad_io_tensor_rd_0_data_bits_19_15),
    .io_tensor_rd_0_data_bits_20_0(tensorLoad_io_tensor_rd_0_data_bits_20_0),
    .io_tensor_rd_0_data_bits_20_1(tensorLoad_io_tensor_rd_0_data_bits_20_1),
    .io_tensor_rd_0_data_bits_20_2(tensorLoad_io_tensor_rd_0_data_bits_20_2),
    .io_tensor_rd_0_data_bits_20_3(tensorLoad_io_tensor_rd_0_data_bits_20_3),
    .io_tensor_rd_0_data_bits_20_4(tensorLoad_io_tensor_rd_0_data_bits_20_4),
    .io_tensor_rd_0_data_bits_20_5(tensorLoad_io_tensor_rd_0_data_bits_20_5),
    .io_tensor_rd_0_data_bits_20_6(tensorLoad_io_tensor_rd_0_data_bits_20_6),
    .io_tensor_rd_0_data_bits_20_7(tensorLoad_io_tensor_rd_0_data_bits_20_7),
    .io_tensor_rd_0_data_bits_20_8(tensorLoad_io_tensor_rd_0_data_bits_20_8),
    .io_tensor_rd_0_data_bits_20_9(tensorLoad_io_tensor_rd_0_data_bits_20_9),
    .io_tensor_rd_0_data_bits_20_10(tensorLoad_io_tensor_rd_0_data_bits_20_10),
    .io_tensor_rd_0_data_bits_20_11(tensorLoad_io_tensor_rd_0_data_bits_20_11),
    .io_tensor_rd_0_data_bits_20_12(tensorLoad_io_tensor_rd_0_data_bits_20_12),
    .io_tensor_rd_0_data_bits_20_13(tensorLoad_io_tensor_rd_0_data_bits_20_13),
    .io_tensor_rd_0_data_bits_20_14(tensorLoad_io_tensor_rd_0_data_bits_20_14),
    .io_tensor_rd_0_data_bits_20_15(tensorLoad_io_tensor_rd_0_data_bits_20_15),
    .io_tensor_rd_0_data_bits_21_0(tensorLoad_io_tensor_rd_0_data_bits_21_0),
    .io_tensor_rd_0_data_bits_21_1(tensorLoad_io_tensor_rd_0_data_bits_21_1),
    .io_tensor_rd_0_data_bits_21_2(tensorLoad_io_tensor_rd_0_data_bits_21_2),
    .io_tensor_rd_0_data_bits_21_3(tensorLoad_io_tensor_rd_0_data_bits_21_3),
    .io_tensor_rd_0_data_bits_21_4(tensorLoad_io_tensor_rd_0_data_bits_21_4),
    .io_tensor_rd_0_data_bits_21_5(tensorLoad_io_tensor_rd_0_data_bits_21_5),
    .io_tensor_rd_0_data_bits_21_6(tensorLoad_io_tensor_rd_0_data_bits_21_6),
    .io_tensor_rd_0_data_bits_21_7(tensorLoad_io_tensor_rd_0_data_bits_21_7),
    .io_tensor_rd_0_data_bits_21_8(tensorLoad_io_tensor_rd_0_data_bits_21_8),
    .io_tensor_rd_0_data_bits_21_9(tensorLoad_io_tensor_rd_0_data_bits_21_9),
    .io_tensor_rd_0_data_bits_21_10(tensorLoad_io_tensor_rd_0_data_bits_21_10),
    .io_tensor_rd_0_data_bits_21_11(tensorLoad_io_tensor_rd_0_data_bits_21_11),
    .io_tensor_rd_0_data_bits_21_12(tensorLoad_io_tensor_rd_0_data_bits_21_12),
    .io_tensor_rd_0_data_bits_21_13(tensorLoad_io_tensor_rd_0_data_bits_21_13),
    .io_tensor_rd_0_data_bits_21_14(tensorLoad_io_tensor_rd_0_data_bits_21_14),
    .io_tensor_rd_0_data_bits_21_15(tensorLoad_io_tensor_rd_0_data_bits_21_15),
    .io_tensor_rd_0_data_bits_22_0(tensorLoad_io_tensor_rd_0_data_bits_22_0),
    .io_tensor_rd_0_data_bits_22_1(tensorLoad_io_tensor_rd_0_data_bits_22_1),
    .io_tensor_rd_0_data_bits_22_2(tensorLoad_io_tensor_rd_0_data_bits_22_2),
    .io_tensor_rd_0_data_bits_22_3(tensorLoad_io_tensor_rd_0_data_bits_22_3),
    .io_tensor_rd_0_data_bits_22_4(tensorLoad_io_tensor_rd_0_data_bits_22_4),
    .io_tensor_rd_0_data_bits_22_5(tensorLoad_io_tensor_rd_0_data_bits_22_5),
    .io_tensor_rd_0_data_bits_22_6(tensorLoad_io_tensor_rd_0_data_bits_22_6),
    .io_tensor_rd_0_data_bits_22_7(tensorLoad_io_tensor_rd_0_data_bits_22_7),
    .io_tensor_rd_0_data_bits_22_8(tensorLoad_io_tensor_rd_0_data_bits_22_8),
    .io_tensor_rd_0_data_bits_22_9(tensorLoad_io_tensor_rd_0_data_bits_22_9),
    .io_tensor_rd_0_data_bits_22_10(tensorLoad_io_tensor_rd_0_data_bits_22_10),
    .io_tensor_rd_0_data_bits_22_11(tensorLoad_io_tensor_rd_0_data_bits_22_11),
    .io_tensor_rd_0_data_bits_22_12(tensorLoad_io_tensor_rd_0_data_bits_22_12),
    .io_tensor_rd_0_data_bits_22_13(tensorLoad_io_tensor_rd_0_data_bits_22_13),
    .io_tensor_rd_0_data_bits_22_14(tensorLoad_io_tensor_rd_0_data_bits_22_14),
    .io_tensor_rd_0_data_bits_22_15(tensorLoad_io_tensor_rd_0_data_bits_22_15),
    .io_tensor_rd_0_data_bits_23_0(tensorLoad_io_tensor_rd_0_data_bits_23_0),
    .io_tensor_rd_0_data_bits_23_1(tensorLoad_io_tensor_rd_0_data_bits_23_1),
    .io_tensor_rd_0_data_bits_23_2(tensorLoad_io_tensor_rd_0_data_bits_23_2),
    .io_tensor_rd_0_data_bits_23_3(tensorLoad_io_tensor_rd_0_data_bits_23_3),
    .io_tensor_rd_0_data_bits_23_4(tensorLoad_io_tensor_rd_0_data_bits_23_4),
    .io_tensor_rd_0_data_bits_23_5(tensorLoad_io_tensor_rd_0_data_bits_23_5),
    .io_tensor_rd_0_data_bits_23_6(tensorLoad_io_tensor_rd_0_data_bits_23_6),
    .io_tensor_rd_0_data_bits_23_7(tensorLoad_io_tensor_rd_0_data_bits_23_7),
    .io_tensor_rd_0_data_bits_23_8(tensorLoad_io_tensor_rd_0_data_bits_23_8),
    .io_tensor_rd_0_data_bits_23_9(tensorLoad_io_tensor_rd_0_data_bits_23_9),
    .io_tensor_rd_0_data_bits_23_10(tensorLoad_io_tensor_rd_0_data_bits_23_10),
    .io_tensor_rd_0_data_bits_23_11(tensorLoad_io_tensor_rd_0_data_bits_23_11),
    .io_tensor_rd_0_data_bits_23_12(tensorLoad_io_tensor_rd_0_data_bits_23_12),
    .io_tensor_rd_0_data_bits_23_13(tensorLoad_io_tensor_rd_0_data_bits_23_13),
    .io_tensor_rd_0_data_bits_23_14(tensorLoad_io_tensor_rd_0_data_bits_23_14),
    .io_tensor_rd_0_data_bits_23_15(tensorLoad_io_tensor_rd_0_data_bits_23_15),
    .io_tensor_rd_0_data_bits_24_0(tensorLoad_io_tensor_rd_0_data_bits_24_0),
    .io_tensor_rd_0_data_bits_24_1(tensorLoad_io_tensor_rd_0_data_bits_24_1),
    .io_tensor_rd_0_data_bits_24_2(tensorLoad_io_tensor_rd_0_data_bits_24_2),
    .io_tensor_rd_0_data_bits_24_3(tensorLoad_io_tensor_rd_0_data_bits_24_3),
    .io_tensor_rd_0_data_bits_24_4(tensorLoad_io_tensor_rd_0_data_bits_24_4),
    .io_tensor_rd_0_data_bits_24_5(tensorLoad_io_tensor_rd_0_data_bits_24_5),
    .io_tensor_rd_0_data_bits_24_6(tensorLoad_io_tensor_rd_0_data_bits_24_6),
    .io_tensor_rd_0_data_bits_24_7(tensorLoad_io_tensor_rd_0_data_bits_24_7),
    .io_tensor_rd_0_data_bits_24_8(tensorLoad_io_tensor_rd_0_data_bits_24_8),
    .io_tensor_rd_0_data_bits_24_9(tensorLoad_io_tensor_rd_0_data_bits_24_9),
    .io_tensor_rd_0_data_bits_24_10(tensorLoad_io_tensor_rd_0_data_bits_24_10),
    .io_tensor_rd_0_data_bits_24_11(tensorLoad_io_tensor_rd_0_data_bits_24_11),
    .io_tensor_rd_0_data_bits_24_12(tensorLoad_io_tensor_rd_0_data_bits_24_12),
    .io_tensor_rd_0_data_bits_24_13(tensorLoad_io_tensor_rd_0_data_bits_24_13),
    .io_tensor_rd_0_data_bits_24_14(tensorLoad_io_tensor_rd_0_data_bits_24_14),
    .io_tensor_rd_0_data_bits_24_15(tensorLoad_io_tensor_rd_0_data_bits_24_15),
    .io_tensor_rd_0_data_bits_25_0(tensorLoad_io_tensor_rd_0_data_bits_25_0),
    .io_tensor_rd_0_data_bits_25_1(tensorLoad_io_tensor_rd_0_data_bits_25_1),
    .io_tensor_rd_0_data_bits_25_2(tensorLoad_io_tensor_rd_0_data_bits_25_2),
    .io_tensor_rd_0_data_bits_25_3(tensorLoad_io_tensor_rd_0_data_bits_25_3),
    .io_tensor_rd_0_data_bits_25_4(tensorLoad_io_tensor_rd_0_data_bits_25_4),
    .io_tensor_rd_0_data_bits_25_5(tensorLoad_io_tensor_rd_0_data_bits_25_5),
    .io_tensor_rd_0_data_bits_25_6(tensorLoad_io_tensor_rd_0_data_bits_25_6),
    .io_tensor_rd_0_data_bits_25_7(tensorLoad_io_tensor_rd_0_data_bits_25_7),
    .io_tensor_rd_0_data_bits_25_8(tensorLoad_io_tensor_rd_0_data_bits_25_8),
    .io_tensor_rd_0_data_bits_25_9(tensorLoad_io_tensor_rd_0_data_bits_25_9),
    .io_tensor_rd_0_data_bits_25_10(tensorLoad_io_tensor_rd_0_data_bits_25_10),
    .io_tensor_rd_0_data_bits_25_11(tensorLoad_io_tensor_rd_0_data_bits_25_11),
    .io_tensor_rd_0_data_bits_25_12(tensorLoad_io_tensor_rd_0_data_bits_25_12),
    .io_tensor_rd_0_data_bits_25_13(tensorLoad_io_tensor_rd_0_data_bits_25_13),
    .io_tensor_rd_0_data_bits_25_14(tensorLoad_io_tensor_rd_0_data_bits_25_14),
    .io_tensor_rd_0_data_bits_25_15(tensorLoad_io_tensor_rd_0_data_bits_25_15),
    .io_tensor_rd_0_data_bits_26_0(tensorLoad_io_tensor_rd_0_data_bits_26_0),
    .io_tensor_rd_0_data_bits_26_1(tensorLoad_io_tensor_rd_0_data_bits_26_1),
    .io_tensor_rd_0_data_bits_26_2(tensorLoad_io_tensor_rd_0_data_bits_26_2),
    .io_tensor_rd_0_data_bits_26_3(tensorLoad_io_tensor_rd_0_data_bits_26_3),
    .io_tensor_rd_0_data_bits_26_4(tensorLoad_io_tensor_rd_0_data_bits_26_4),
    .io_tensor_rd_0_data_bits_26_5(tensorLoad_io_tensor_rd_0_data_bits_26_5),
    .io_tensor_rd_0_data_bits_26_6(tensorLoad_io_tensor_rd_0_data_bits_26_6),
    .io_tensor_rd_0_data_bits_26_7(tensorLoad_io_tensor_rd_0_data_bits_26_7),
    .io_tensor_rd_0_data_bits_26_8(tensorLoad_io_tensor_rd_0_data_bits_26_8),
    .io_tensor_rd_0_data_bits_26_9(tensorLoad_io_tensor_rd_0_data_bits_26_9),
    .io_tensor_rd_0_data_bits_26_10(tensorLoad_io_tensor_rd_0_data_bits_26_10),
    .io_tensor_rd_0_data_bits_26_11(tensorLoad_io_tensor_rd_0_data_bits_26_11),
    .io_tensor_rd_0_data_bits_26_12(tensorLoad_io_tensor_rd_0_data_bits_26_12),
    .io_tensor_rd_0_data_bits_26_13(tensorLoad_io_tensor_rd_0_data_bits_26_13),
    .io_tensor_rd_0_data_bits_26_14(tensorLoad_io_tensor_rd_0_data_bits_26_14),
    .io_tensor_rd_0_data_bits_26_15(tensorLoad_io_tensor_rd_0_data_bits_26_15),
    .io_tensor_rd_0_data_bits_27_0(tensorLoad_io_tensor_rd_0_data_bits_27_0),
    .io_tensor_rd_0_data_bits_27_1(tensorLoad_io_tensor_rd_0_data_bits_27_1),
    .io_tensor_rd_0_data_bits_27_2(tensorLoad_io_tensor_rd_0_data_bits_27_2),
    .io_tensor_rd_0_data_bits_27_3(tensorLoad_io_tensor_rd_0_data_bits_27_3),
    .io_tensor_rd_0_data_bits_27_4(tensorLoad_io_tensor_rd_0_data_bits_27_4),
    .io_tensor_rd_0_data_bits_27_5(tensorLoad_io_tensor_rd_0_data_bits_27_5),
    .io_tensor_rd_0_data_bits_27_6(tensorLoad_io_tensor_rd_0_data_bits_27_6),
    .io_tensor_rd_0_data_bits_27_7(tensorLoad_io_tensor_rd_0_data_bits_27_7),
    .io_tensor_rd_0_data_bits_27_8(tensorLoad_io_tensor_rd_0_data_bits_27_8),
    .io_tensor_rd_0_data_bits_27_9(tensorLoad_io_tensor_rd_0_data_bits_27_9),
    .io_tensor_rd_0_data_bits_27_10(tensorLoad_io_tensor_rd_0_data_bits_27_10),
    .io_tensor_rd_0_data_bits_27_11(tensorLoad_io_tensor_rd_0_data_bits_27_11),
    .io_tensor_rd_0_data_bits_27_12(tensorLoad_io_tensor_rd_0_data_bits_27_12),
    .io_tensor_rd_0_data_bits_27_13(tensorLoad_io_tensor_rd_0_data_bits_27_13),
    .io_tensor_rd_0_data_bits_27_14(tensorLoad_io_tensor_rd_0_data_bits_27_14),
    .io_tensor_rd_0_data_bits_27_15(tensorLoad_io_tensor_rd_0_data_bits_27_15),
    .io_tensor_rd_0_data_bits_28_0(tensorLoad_io_tensor_rd_0_data_bits_28_0),
    .io_tensor_rd_0_data_bits_28_1(tensorLoad_io_tensor_rd_0_data_bits_28_1),
    .io_tensor_rd_0_data_bits_28_2(tensorLoad_io_tensor_rd_0_data_bits_28_2),
    .io_tensor_rd_0_data_bits_28_3(tensorLoad_io_tensor_rd_0_data_bits_28_3),
    .io_tensor_rd_0_data_bits_28_4(tensorLoad_io_tensor_rd_0_data_bits_28_4),
    .io_tensor_rd_0_data_bits_28_5(tensorLoad_io_tensor_rd_0_data_bits_28_5),
    .io_tensor_rd_0_data_bits_28_6(tensorLoad_io_tensor_rd_0_data_bits_28_6),
    .io_tensor_rd_0_data_bits_28_7(tensorLoad_io_tensor_rd_0_data_bits_28_7),
    .io_tensor_rd_0_data_bits_28_8(tensorLoad_io_tensor_rd_0_data_bits_28_8),
    .io_tensor_rd_0_data_bits_28_9(tensorLoad_io_tensor_rd_0_data_bits_28_9),
    .io_tensor_rd_0_data_bits_28_10(tensorLoad_io_tensor_rd_0_data_bits_28_10),
    .io_tensor_rd_0_data_bits_28_11(tensorLoad_io_tensor_rd_0_data_bits_28_11),
    .io_tensor_rd_0_data_bits_28_12(tensorLoad_io_tensor_rd_0_data_bits_28_12),
    .io_tensor_rd_0_data_bits_28_13(tensorLoad_io_tensor_rd_0_data_bits_28_13),
    .io_tensor_rd_0_data_bits_28_14(tensorLoad_io_tensor_rd_0_data_bits_28_14),
    .io_tensor_rd_0_data_bits_28_15(tensorLoad_io_tensor_rd_0_data_bits_28_15),
    .io_tensor_rd_0_data_bits_29_0(tensorLoad_io_tensor_rd_0_data_bits_29_0),
    .io_tensor_rd_0_data_bits_29_1(tensorLoad_io_tensor_rd_0_data_bits_29_1),
    .io_tensor_rd_0_data_bits_29_2(tensorLoad_io_tensor_rd_0_data_bits_29_2),
    .io_tensor_rd_0_data_bits_29_3(tensorLoad_io_tensor_rd_0_data_bits_29_3),
    .io_tensor_rd_0_data_bits_29_4(tensorLoad_io_tensor_rd_0_data_bits_29_4),
    .io_tensor_rd_0_data_bits_29_5(tensorLoad_io_tensor_rd_0_data_bits_29_5),
    .io_tensor_rd_0_data_bits_29_6(tensorLoad_io_tensor_rd_0_data_bits_29_6),
    .io_tensor_rd_0_data_bits_29_7(tensorLoad_io_tensor_rd_0_data_bits_29_7),
    .io_tensor_rd_0_data_bits_29_8(tensorLoad_io_tensor_rd_0_data_bits_29_8),
    .io_tensor_rd_0_data_bits_29_9(tensorLoad_io_tensor_rd_0_data_bits_29_9),
    .io_tensor_rd_0_data_bits_29_10(tensorLoad_io_tensor_rd_0_data_bits_29_10),
    .io_tensor_rd_0_data_bits_29_11(tensorLoad_io_tensor_rd_0_data_bits_29_11),
    .io_tensor_rd_0_data_bits_29_12(tensorLoad_io_tensor_rd_0_data_bits_29_12),
    .io_tensor_rd_0_data_bits_29_13(tensorLoad_io_tensor_rd_0_data_bits_29_13),
    .io_tensor_rd_0_data_bits_29_14(tensorLoad_io_tensor_rd_0_data_bits_29_14),
    .io_tensor_rd_0_data_bits_29_15(tensorLoad_io_tensor_rd_0_data_bits_29_15),
    .io_tensor_rd_0_data_bits_30_0(tensorLoad_io_tensor_rd_0_data_bits_30_0),
    .io_tensor_rd_0_data_bits_30_1(tensorLoad_io_tensor_rd_0_data_bits_30_1),
    .io_tensor_rd_0_data_bits_30_2(tensorLoad_io_tensor_rd_0_data_bits_30_2),
    .io_tensor_rd_0_data_bits_30_3(tensorLoad_io_tensor_rd_0_data_bits_30_3),
    .io_tensor_rd_0_data_bits_30_4(tensorLoad_io_tensor_rd_0_data_bits_30_4),
    .io_tensor_rd_0_data_bits_30_5(tensorLoad_io_tensor_rd_0_data_bits_30_5),
    .io_tensor_rd_0_data_bits_30_6(tensorLoad_io_tensor_rd_0_data_bits_30_6),
    .io_tensor_rd_0_data_bits_30_7(tensorLoad_io_tensor_rd_0_data_bits_30_7),
    .io_tensor_rd_0_data_bits_30_8(tensorLoad_io_tensor_rd_0_data_bits_30_8),
    .io_tensor_rd_0_data_bits_30_9(tensorLoad_io_tensor_rd_0_data_bits_30_9),
    .io_tensor_rd_0_data_bits_30_10(tensorLoad_io_tensor_rd_0_data_bits_30_10),
    .io_tensor_rd_0_data_bits_30_11(tensorLoad_io_tensor_rd_0_data_bits_30_11),
    .io_tensor_rd_0_data_bits_30_12(tensorLoad_io_tensor_rd_0_data_bits_30_12),
    .io_tensor_rd_0_data_bits_30_13(tensorLoad_io_tensor_rd_0_data_bits_30_13),
    .io_tensor_rd_0_data_bits_30_14(tensorLoad_io_tensor_rd_0_data_bits_30_14),
    .io_tensor_rd_0_data_bits_30_15(tensorLoad_io_tensor_rd_0_data_bits_30_15),
    .io_tensor_rd_0_data_bits_31_0(tensorLoad_io_tensor_rd_0_data_bits_31_0),
    .io_tensor_rd_0_data_bits_31_1(tensorLoad_io_tensor_rd_0_data_bits_31_1),
    .io_tensor_rd_0_data_bits_31_2(tensorLoad_io_tensor_rd_0_data_bits_31_2),
    .io_tensor_rd_0_data_bits_31_3(tensorLoad_io_tensor_rd_0_data_bits_31_3),
    .io_tensor_rd_0_data_bits_31_4(tensorLoad_io_tensor_rd_0_data_bits_31_4),
    .io_tensor_rd_0_data_bits_31_5(tensorLoad_io_tensor_rd_0_data_bits_31_5),
    .io_tensor_rd_0_data_bits_31_6(tensorLoad_io_tensor_rd_0_data_bits_31_6),
    .io_tensor_rd_0_data_bits_31_7(tensorLoad_io_tensor_rd_0_data_bits_31_7),
    .io_tensor_rd_0_data_bits_31_8(tensorLoad_io_tensor_rd_0_data_bits_31_8),
    .io_tensor_rd_0_data_bits_31_9(tensorLoad_io_tensor_rd_0_data_bits_31_9),
    .io_tensor_rd_0_data_bits_31_10(tensorLoad_io_tensor_rd_0_data_bits_31_10),
    .io_tensor_rd_0_data_bits_31_11(tensorLoad_io_tensor_rd_0_data_bits_31_11),
    .io_tensor_rd_0_data_bits_31_12(tensorLoad_io_tensor_rd_0_data_bits_31_12),
    .io_tensor_rd_0_data_bits_31_13(tensorLoad_io_tensor_rd_0_data_bits_31_13),
    .io_tensor_rd_0_data_bits_31_14(tensorLoad_io_tensor_rd_0_data_bits_31_14),
    .io_tensor_rd_0_data_bits_31_15(tensorLoad_io_tensor_rd_0_data_bits_31_15)
  );
  assign io_done = tensorLoad_io_done; // @[TensorLoad.scala 72:8]
  assign io_vme_rd_cmd_valid = tensorLoad_io_vme_rd_cmd_valid; // @[TensorLoad.scala 72:8]
  assign io_vme_rd_cmd_bits_addr = tensorLoad_io_vme_rd_cmd_bits_addr; // @[TensorLoad.scala 72:8]
  assign io_vme_rd_cmd_bits_len = tensorLoad_io_vme_rd_cmd_bits_len; // @[TensorLoad.scala 72:8]
  assign io_vme_rd_cmd_bits_tag = tensorLoad_io_vme_rd_cmd_bits_tag; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_valid = tensorLoad_io_tensor_rd_0_data_valid; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_0 = tensorLoad_io_tensor_rd_0_data_bits_0_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_1 = tensorLoad_io_tensor_rd_0_data_bits_0_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_2 = tensorLoad_io_tensor_rd_0_data_bits_0_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_3 = tensorLoad_io_tensor_rd_0_data_bits_0_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_4 = tensorLoad_io_tensor_rd_0_data_bits_0_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_5 = tensorLoad_io_tensor_rd_0_data_bits_0_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_6 = tensorLoad_io_tensor_rd_0_data_bits_0_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_7 = tensorLoad_io_tensor_rd_0_data_bits_0_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_8 = tensorLoad_io_tensor_rd_0_data_bits_0_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_9 = tensorLoad_io_tensor_rd_0_data_bits_0_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_10 = tensorLoad_io_tensor_rd_0_data_bits_0_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_11 = tensorLoad_io_tensor_rd_0_data_bits_0_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_12 = tensorLoad_io_tensor_rd_0_data_bits_0_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_13 = tensorLoad_io_tensor_rd_0_data_bits_0_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_14 = tensorLoad_io_tensor_rd_0_data_bits_0_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_15 = tensorLoad_io_tensor_rd_0_data_bits_0_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_1_0 = tensorLoad_io_tensor_rd_0_data_bits_1_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_1_1 = tensorLoad_io_tensor_rd_0_data_bits_1_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_1_2 = tensorLoad_io_tensor_rd_0_data_bits_1_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_1_3 = tensorLoad_io_tensor_rd_0_data_bits_1_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_1_4 = tensorLoad_io_tensor_rd_0_data_bits_1_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_1_5 = tensorLoad_io_tensor_rd_0_data_bits_1_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_1_6 = tensorLoad_io_tensor_rd_0_data_bits_1_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_1_7 = tensorLoad_io_tensor_rd_0_data_bits_1_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_1_8 = tensorLoad_io_tensor_rd_0_data_bits_1_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_1_9 = tensorLoad_io_tensor_rd_0_data_bits_1_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_1_10 = tensorLoad_io_tensor_rd_0_data_bits_1_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_1_11 = tensorLoad_io_tensor_rd_0_data_bits_1_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_1_12 = tensorLoad_io_tensor_rd_0_data_bits_1_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_1_13 = tensorLoad_io_tensor_rd_0_data_bits_1_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_1_14 = tensorLoad_io_tensor_rd_0_data_bits_1_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_1_15 = tensorLoad_io_tensor_rd_0_data_bits_1_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_2_0 = tensorLoad_io_tensor_rd_0_data_bits_2_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_2_1 = tensorLoad_io_tensor_rd_0_data_bits_2_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_2_2 = tensorLoad_io_tensor_rd_0_data_bits_2_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_2_3 = tensorLoad_io_tensor_rd_0_data_bits_2_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_2_4 = tensorLoad_io_tensor_rd_0_data_bits_2_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_2_5 = tensorLoad_io_tensor_rd_0_data_bits_2_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_2_6 = tensorLoad_io_tensor_rd_0_data_bits_2_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_2_7 = tensorLoad_io_tensor_rd_0_data_bits_2_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_2_8 = tensorLoad_io_tensor_rd_0_data_bits_2_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_2_9 = tensorLoad_io_tensor_rd_0_data_bits_2_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_2_10 = tensorLoad_io_tensor_rd_0_data_bits_2_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_2_11 = tensorLoad_io_tensor_rd_0_data_bits_2_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_2_12 = tensorLoad_io_tensor_rd_0_data_bits_2_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_2_13 = tensorLoad_io_tensor_rd_0_data_bits_2_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_2_14 = tensorLoad_io_tensor_rd_0_data_bits_2_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_2_15 = tensorLoad_io_tensor_rd_0_data_bits_2_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_3_0 = tensorLoad_io_tensor_rd_0_data_bits_3_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_3_1 = tensorLoad_io_tensor_rd_0_data_bits_3_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_3_2 = tensorLoad_io_tensor_rd_0_data_bits_3_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_3_3 = tensorLoad_io_tensor_rd_0_data_bits_3_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_3_4 = tensorLoad_io_tensor_rd_0_data_bits_3_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_3_5 = tensorLoad_io_tensor_rd_0_data_bits_3_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_3_6 = tensorLoad_io_tensor_rd_0_data_bits_3_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_3_7 = tensorLoad_io_tensor_rd_0_data_bits_3_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_3_8 = tensorLoad_io_tensor_rd_0_data_bits_3_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_3_9 = tensorLoad_io_tensor_rd_0_data_bits_3_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_3_10 = tensorLoad_io_tensor_rd_0_data_bits_3_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_3_11 = tensorLoad_io_tensor_rd_0_data_bits_3_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_3_12 = tensorLoad_io_tensor_rd_0_data_bits_3_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_3_13 = tensorLoad_io_tensor_rd_0_data_bits_3_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_3_14 = tensorLoad_io_tensor_rd_0_data_bits_3_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_3_15 = tensorLoad_io_tensor_rd_0_data_bits_3_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_4_0 = tensorLoad_io_tensor_rd_0_data_bits_4_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_4_1 = tensorLoad_io_tensor_rd_0_data_bits_4_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_4_2 = tensorLoad_io_tensor_rd_0_data_bits_4_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_4_3 = tensorLoad_io_tensor_rd_0_data_bits_4_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_4_4 = tensorLoad_io_tensor_rd_0_data_bits_4_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_4_5 = tensorLoad_io_tensor_rd_0_data_bits_4_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_4_6 = tensorLoad_io_tensor_rd_0_data_bits_4_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_4_7 = tensorLoad_io_tensor_rd_0_data_bits_4_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_4_8 = tensorLoad_io_tensor_rd_0_data_bits_4_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_4_9 = tensorLoad_io_tensor_rd_0_data_bits_4_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_4_10 = tensorLoad_io_tensor_rd_0_data_bits_4_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_4_11 = tensorLoad_io_tensor_rd_0_data_bits_4_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_4_12 = tensorLoad_io_tensor_rd_0_data_bits_4_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_4_13 = tensorLoad_io_tensor_rd_0_data_bits_4_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_4_14 = tensorLoad_io_tensor_rd_0_data_bits_4_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_4_15 = tensorLoad_io_tensor_rd_0_data_bits_4_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_5_0 = tensorLoad_io_tensor_rd_0_data_bits_5_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_5_1 = tensorLoad_io_tensor_rd_0_data_bits_5_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_5_2 = tensorLoad_io_tensor_rd_0_data_bits_5_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_5_3 = tensorLoad_io_tensor_rd_0_data_bits_5_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_5_4 = tensorLoad_io_tensor_rd_0_data_bits_5_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_5_5 = tensorLoad_io_tensor_rd_0_data_bits_5_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_5_6 = tensorLoad_io_tensor_rd_0_data_bits_5_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_5_7 = tensorLoad_io_tensor_rd_0_data_bits_5_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_5_8 = tensorLoad_io_tensor_rd_0_data_bits_5_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_5_9 = tensorLoad_io_tensor_rd_0_data_bits_5_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_5_10 = tensorLoad_io_tensor_rd_0_data_bits_5_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_5_11 = tensorLoad_io_tensor_rd_0_data_bits_5_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_5_12 = tensorLoad_io_tensor_rd_0_data_bits_5_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_5_13 = tensorLoad_io_tensor_rd_0_data_bits_5_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_5_14 = tensorLoad_io_tensor_rd_0_data_bits_5_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_5_15 = tensorLoad_io_tensor_rd_0_data_bits_5_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_6_0 = tensorLoad_io_tensor_rd_0_data_bits_6_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_6_1 = tensorLoad_io_tensor_rd_0_data_bits_6_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_6_2 = tensorLoad_io_tensor_rd_0_data_bits_6_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_6_3 = tensorLoad_io_tensor_rd_0_data_bits_6_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_6_4 = tensorLoad_io_tensor_rd_0_data_bits_6_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_6_5 = tensorLoad_io_tensor_rd_0_data_bits_6_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_6_6 = tensorLoad_io_tensor_rd_0_data_bits_6_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_6_7 = tensorLoad_io_tensor_rd_0_data_bits_6_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_6_8 = tensorLoad_io_tensor_rd_0_data_bits_6_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_6_9 = tensorLoad_io_tensor_rd_0_data_bits_6_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_6_10 = tensorLoad_io_tensor_rd_0_data_bits_6_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_6_11 = tensorLoad_io_tensor_rd_0_data_bits_6_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_6_12 = tensorLoad_io_tensor_rd_0_data_bits_6_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_6_13 = tensorLoad_io_tensor_rd_0_data_bits_6_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_6_14 = tensorLoad_io_tensor_rd_0_data_bits_6_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_6_15 = tensorLoad_io_tensor_rd_0_data_bits_6_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_7_0 = tensorLoad_io_tensor_rd_0_data_bits_7_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_7_1 = tensorLoad_io_tensor_rd_0_data_bits_7_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_7_2 = tensorLoad_io_tensor_rd_0_data_bits_7_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_7_3 = tensorLoad_io_tensor_rd_0_data_bits_7_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_7_4 = tensorLoad_io_tensor_rd_0_data_bits_7_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_7_5 = tensorLoad_io_tensor_rd_0_data_bits_7_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_7_6 = tensorLoad_io_tensor_rd_0_data_bits_7_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_7_7 = tensorLoad_io_tensor_rd_0_data_bits_7_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_7_8 = tensorLoad_io_tensor_rd_0_data_bits_7_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_7_9 = tensorLoad_io_tensor_rd_0_data_bits_7_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_7_10 = tensorLoad_io_tensor_rd_0_data_bits_7_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_7_11 = tensorLoad_io_tensor_rd_0_data_bits_7_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_7_12 = tensorLoad_io_tensor_rd_0_data_bits_7_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_7_13 = tensorLoad_io_tensor_rd_0_data_bits_7_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_7_14 = tensorLoad_io_tensor_rd_0_data_bits_7_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_7_15 = tensorLoad_io_tensor_rd_0_data_bits_7_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_8_0 = tensorLoad_io_tensor_rd_0_data_bits_8_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_8_1 = tensorLoad_io_tensor_rd_0_data_bits_8_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_8_2 = tensorLoad_io_tensor_rd_0_data_bits_8_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_8_3 = tensorLoad_io_tensor_rd_0_data_bits_8_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_8_4 = tensorLoad_io_tensor_rd_0_data_bits_8_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_8_5 = tensorLoad_io_tensor_rd_0_data_bits_8_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_8_6 = tensorLoad_io_tensor_rd_0_data_bits_8_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_8_7 = tensorLoad_io_tensor_rd_0_data_bits_8_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_8_8 = tensorLoad_io_tensor_rd_0_data_bits_8_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_8_9 = tensorLoad_io_tensor_rd_0_data_bits_8_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_8_10 = tensorLoad_io_tensor_rd_0_data_bits_8_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_8_11 = tensorLoad_io_tensor_rd_0_data_bits_8_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_8_12 = tensorLoad_io_tensor_rd_0_data_bits_8_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_8_13 = tensorLoad_io_tensor_rd_0_data_bits_8_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_8_14 = tensorLoad_io_tensor_rd_0_data_bits_8_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_8_15 = tensorLoad_io_tensor_rd_0_data_bits_8_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_9_0 = tensorLoad_io_tensor_rd_0_data_bits_9_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_9_1 = tensorLoad_io_tensor_rd_0_data_bits_9_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_9_2 = tensorLoad_io_tensor_rd_0_data_bits_9_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_9_3 = tensorLoad_io_tensor_rd_0_data_bits_9_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_9_4 = tensorLoad_io_tensor_rd_0_data_bits_9_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_9_5 = tensorLoad_io_tensor_rd_0_data_bits_9_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_9_6 = tensorLoad_io_tensor_rd_0_data_bits_9_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_9_7 = tensorLoad_io_tensor_rd_0_data_bits_9_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_9_8 = tensorLoad_io_tensor_rd_0_data_bits_9_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_9_9 = tensorLoad_io_tensor_rd_0_data_bits_9_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_9_10 = tensorLoad_io_tensor_rd_0_data_bits_9_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_9_11 = tensorLoad_io_tensor_rd_0_data_bits_9_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_9_12 = tensorLoad_io_tensor_rd_0_data_bits_9_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_9_13 = tensorLoad_io_tensor_rd_0_data_bits_9_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_9_14 = tensorLoad_io_tensor_rd_0_data_bits_9_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_9_15 = tensorLoad_io_tensor_rd_0_data_bits_9_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_10_0 = tensorLoad_io_tensor_rd_0_data_bits_10_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_10_1 = tensorLoad_io_tensor_rd_0_data_bits_10_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_10_2 = tensorLoad_io_tensor_rd_0_data_bits_10_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_10_3 = tensorLoad_io_tensor_rd_0_data_bits_10_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_10_4 = tensorLoad_io_tensor_rd_0_data_bits_10_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_10_5 = tensorLoad_io_tensor_rd_0_data_bits_10_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_10_6 = tensorLoad_io_tensor_rd_0_data_bits_10_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_10_7 = tensorLoad_io_tensor_rd_0_data_bits_10_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_10_8 = tensorLoad_io_tensor_rd_0_data_bits_10_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_10_9 = tensorLoad_io_tensor_rd_0_data_bits_10_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_10_10 = tensorLoad_io_tensor_rd_0_data_bits_10_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_10_11 = tensorLoad_io_tensor_rd_0_data_bits_10_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_10_12 = tensorLoad_io_tensor_rd_0_data_bits_10_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_10_13 = tensorLoad_io_tensor_rd_0_data_bits_10_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_10_14 = tensorLoad_io_tensor_rd_0_data_bits_10_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_10_15 = tensorLoad_io_tensor_rd_0_data_bits_10_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_11_0 = tensorLoad_io_tensor_rd_0_data_bits_11_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_11_1 = tensorLoad_io_tensor_rd_0_data_bits_11_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_11_2 = tensorLoad_io_tensor_rd_0_data_bits_11_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_11_3 = tensorLoad_io_tensor_rd_0_data_bits_11_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_11_4 = tensorLoad_io_tensor_rd_0_data_bits_11_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_11_5 = tensorLoad_io_tensor_rd_0_data_bits_11_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_11_6 = tensorLoad_io_tensor_rd_0_data_bits_11_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_11_7 = tensorLoad_io_tensor_rd_0_data_bits_11_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_11_8 = tensorLoad_io_tensor_rd_0_data_bits_11_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_11_9 = tensorLoad_io_tensor_rd_0_data_bits_11_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_11_10 = tensorLoad_io_tensor_rd_0_data_bits_11_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_11_11 = tensorLoad_io_tensor_rd_0_data_bits_11_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_11_12 = tensorLoad_io_tensor_rd_0_data_bits_11_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_11_13 = tensorLoad_io_tensor_rd_0_data_bits_11_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_11_14 = tensorLoad_io_tensor_rd_0_data_bits_11_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_11_15 = tensorLoad_io_tensor_rd_0_data_bits_11_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_12_0 = tensorLoad_io_tensor_rd_0_data_bits_12_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_12_1 = tensorLoad_io_tensor_rd_0_data_bits_12_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_12_2 = tensorLoad_io_tensor_rd_0_data_bits_12_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_12_3 = tensorLoad_io_tensor_rd_0_data_bits_12_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_12_4 = tensorLoad_io_tensor_rd_0_data_bits_12_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_12_5 = tensorLoad_io_tensor_rd_0_data_bits_12_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_12_6 = tensorLoad_io_tensor_rd_0_data_bits_12_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_12_7 = tensorLoad_io_tensor_rd_0_data_bits_12_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_12_8 = tensorLoad_io_tensor_rd_0_data_bits_12_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_12_9 = tensorLoad_io_tensor_rd_0_data_bits_12_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_12_10 = tensorLoad_io_tensor_rd_0_data_bits_12_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_12_11 = tensorLoad_io_tensor_rd_0_data_bits_12_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_12_12 = tensorLoad_io_tensor_rd_0_data_bits_12_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_12_13 = tensorLoad_io_tensor_rd_0_data_bits_12_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_12_14 = tensorLoad_io_tensor_rd_0_data_bits_12_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_12_15 = tensorLoad_io_tensor_rd_0_data_bits_12_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_13_0 = tensorLoad_io_tensor_rd_0_data_bits_13_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_13_1 = tensorLoad_io_tensor_rd_0_data_bits_13_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_13_2 = tensorLoad_io_tensor_rd_0_data_bits_13_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_13_3 = tensorLoad_io_tensor_rd_0_data_bits_13_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_13_4 = tensorLoad_io_tensor_rd_0_data_bits_13_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_13_5 = tensorLoad_io_tensor_rd_0_data_bits_13_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_13_6 = tensorLoad_io_tensor_rd_0_data_bits_13_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_13_7 = tensorLoad_io_tensor_rd_0_data_bits_13_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_13_8 = tensorLoad_io_tensor_rd_0_data_bits_13_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_13_9 = tensorLoad_io_tensor_rd_0_data_bits_13_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_13_10 = tensorLoad_io_tensor_rd_0_data_bits_13_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_13_11 = tensorLoad_io_tensor_rd_0_data_bits_13_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_13_12 = tensorLoad_io_tensor_rd_0_data_bits_13_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_13_13 = tensorLoad_io_tensor_rd_0_data_bits_13_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_13_14 = tensorLoad_io_tensor_rd_0_data_bits_13_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_13_15 = tensorLoad_io_tensor_rd_0_data_bits_13_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_14_0 = tensorLoad_io_tensor_rd_0_data_bits_14_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_14_1 = tensorLoad_io_tensor_rd_0_data_bits_14_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_14_2 = tensorLoad_io_tensor_rd_0_data_bits_14_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_14_3 = tensorLoad_io_tensor_rd_0_data_bits_14_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_14_4 = tensorLoad_io_tensor_rd_0_data_bits_14_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_14_5 = tensorLoad_io_tensor_rd_0_data_bits_14_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_14_6 = tensorLoad_io_tensor_rd_0_data_bits_14_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_14_7 = tensorLoad_io_tensor_rd_0_data_bits_14_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_14_8 = tensorLoad_io_tensor_rd_0_data_bits_14_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_14_9 = tensorLoad_io_tensor_rd_0_data_bits_14_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_14_10 = tensorLoad_io_tensor_rd_0_data_bits_14_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_14_11 = tensorLoad_io_tensor_rd_0_data_bits_14_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_14_12 = tensorLoad_io_tensor_rd_0_data_bits_14_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_14_13 = tensorLoad_io_tensor_rd_0_data_bits_14_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_14_14 = tensorLoad_io_tensor_rd_0_data_bits_14_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_14_15 = tensorLoad_io_tensor_rd_0_data_bits_14_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_15_0 = tensorLoad_io_tensor_rd_0_data_bits_15_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_15_1 = tensorLoad_io_tensor_rd_0_data_bits_15_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_15_2 = tensorLoad_io_tensor_rd_0_data_bits_15_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_15_3 = tensorLoad_io_tensor_rd_0_data_bits_15_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_15_4 = tensorLoad_io_tensor_rd_0_data_bits_15_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_15_5 = tensorLoad_io_tensor_rd_0_data_bits_15_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_15_6 = tensorLoad_io_tensor_rd_0_data_bits_15_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_15_7 = tensorLoad_io_tensor_rd_0_data_bits_15_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_15_8 = tensorLoad_io_tensor_rd_0_data_bits_15_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_15_9 = tensorLoad_io_tensor_rd_0_data_bits_15_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_15_10 = tensorLoad_io_tensor_rd_0_data_bits_15_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_15_11 = tensorLoad_io_tensor_rd_0_data_bits_15_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_15_12 = tensorLoad_io_tensor_rd_0_data_bits_15_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_15_13 = tensorLoad_io_tensor_rd_0_data_bits_15_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_15_14 = tensorLoad_io_tensor_rd_0_data_bits_15_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_15_15 = tensorLoad_io_tensor_rd_0_data_bits_15_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_16_0 = tensorLoad_io_tensor_rd_0_data_bits_16_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_16_1 = tensorLoad_io_tensor_rd_0_data_bits_16_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_16_2 = tensorLoad_io_tensor_rd_0_data_bits_16_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_16_3 = tensorLoad_io_tensor_rd_0_data_bits_16_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_16_4 = tensorLoad_io_tensor_rd_0_data_bits_16_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_16_5 = tensorLoad_io_tensor_rd_0_data_bits_16_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_16_6 = tensorLoad_io_tensor_rd_0_data_bits_16_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_16_7 = tensorLoad_io_tensor_rd_0_data_bits_16_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_16_8 = tensorLoad_io_tensor_rd_0_data_bits_16_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_16_9 = tensorLoad_io_tensor_rd_0_data_bits_16_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_16_10 = tensorLoad_io_tensor_rd_0_data_bits_16_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_16_11 = tensorLoad_io_tensor_rd_0_data_bits_16_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_16_12 = tensorLoad_io_tensor_rd_0_data_bits_16_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_16_13 = tensorLoad_io_tensor_rd_0_data_bits_16_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_16_14 = tensorLoad_io_tensor_rd_0_data_bits_16_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_16_15 = tensorLoad_io_tensor_rd_0_data_bits_16_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_17_0 = tensorLoad_io_tensor_rd_0_data_bits_17_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_17_1 = tensorLoad_io_tensor_rd_0_data_bits_17_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_17_2 = tensorLoad_io_tensor_rd_0_data_bits_17_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_17_3 = tensorLoad_io_tensor_rd_0_data_bits_17_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_17_4 = tensorLoad_io_tensor_rd_0_data_bits_17_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_17_5 = tensorLoad_io_tensor_rd_0_data_bits_17_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_17_6 = tensorLoad_io_tensor_rd_0_data_bits_17_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_17_7 = tensorLoad_io_tensor_rd_0_data_bits_17_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_17_8 = tensorLoad_io_tensor_rd_0_data_bits_17_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_17_9 = tensorLoad_io_tensor_rd_0_data_bits_17_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_17_10 = tensorLoad_io_tensor_rd_0_data_bits_17_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_17_11 = tensorLoad_io_tensor_rd_0_data_bits_17_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_17_12 = tensorLoad_io_tensor_rd_0_data_bits_17_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_17_13 = tensorLoad_io_tensor_rd_0_data_bits_17_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_17_14 = tensorLoad_io_tensor_rd_0_data_bits_17_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_17_15 = tensorLoad_io_tensor_rd_0_data_bits_17_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_18_0 = tensorLoad_io_tensor_rd_0_data_bits_18_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_18_1 = tensorLoad_io_tensor_rd_0_data_bits_18_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_18_2 = tensorLoad_io_tensor_rd_0_data_bits_18_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_18_3 = tensorLoad_io_tensor_rd_0_data_bits_18_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_18_4 = tensorLoad_io_tensor_rd_0_data_bits_18_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_18_5 = tensorLoad_io_tensor_rd_0_data_bits_18_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_18_6 = tensorLoad_io_tensor_rd_0_data_bits_18_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_18_7 = tensorLoad_io_tensor_rd_0_data_bits_18_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_18_8 = tensorLoad_io_tensor_rd_0_data_bits_18_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_18_9 = tensorLoad_io_tensor_rd_0_data_bits_18_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_18_10 = tensorLoad_io_tensor_rd_0_data_bits_18_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_18_11 = tensorLoad_io_tensor_rd_0_data_bits_18_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_18_12 = tensorLoad_io_tensor_rd_0_data_bits_18_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_18_13 = tensorLoad_io_tensor_rd_0_data_bits_18_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_18_14 = tensorLoad_io_tensor_rd_0_data_bits_18_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_18_15 = tensorLoad_io_tensor_rd_0_data_bits_18_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_19_0 = tensorLoad_io_tensor_rd_0_data_bits_19_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_19_1 = tensorLoad_io_tensor_rd_0_data_bits_19_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_19_2 = tensorLoad_io_tensor_rd_0_data_bits_19_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_19_3 = tensorLoad_io_tensor_rd_0_data_bits_19_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_19_4 = tensorLoad_io_tensor_rd_0_data_bits_19_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_19_5 = tensorLoad_io_tensor_rd_0_data_bits_19_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_19_6 = tensorLoad_io_tensor_rd_0_data_bits_19_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_19_7 = tensorLoad_io_tensor_rd_0_data_bits_19_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_19_8 = tensorLoad_io_tensor_rd_0_data_bits_19_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_19_9 = tensorLoad_io_tensor_rd_0_data_bits_19_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_19_10 = tensorLoad_io_tensor_rd_0_data_bits_19_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_19_11 = tensorLoad_io_tensor_rd_0_data_bits_19_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_19_12 = tensorLoad_io_tensor_rd_0_data_bits_19_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_19_13 = tensorLoad_io_tensor_rd_0_data_bits_19_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_19_14 = tensorLoad_io_tensor_rd_0_data_bits_19_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_19_15 = tensorLoad_io_tensor_rd_0_data_bits_19_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_20_0 = tensorLoad_io_tensor_rd_0_data_bits_20_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_20_1 = tensorLoad_io_tensor_rd_0_data_bits_20_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_20_2 = tensorLoad_io_tensor_rd_0_data_bits_20_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_20_3 = tensorLoad_io_tensor_rd_0_data_bits_20_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_20_4 = tensorLoad_io_tensor_rd_0_data_bits_20_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_20_5 = tensorLoad_io_tensor_rd_0_data_bits_20_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_20_6 = tensorLoad_io_tensor_rd_0_data_bits_20_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_20_7 = tensorLoad_io_tensor_rd_0_data_bits_20_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_20_8 = tensorLoad_io_tensor_rd_0_data_bits_20_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_20_9 = tensorLoad_io_tensor_rd_0_data_bits_20_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_20_10 = tensorLoad_io_tensor_rd_0_data_bits_20_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_20_11 = tensorLoad_io_tensor_rd_0_data_bits_20_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_20_12 = tensorLoad_io_tensor_rd_0_data_bits_20_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_20_13 = tensorLoad_io_tensor_rd_0_data_bits_20_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_20_14 = tensorLoad_io_tensor_rd_0_data_bits_20_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_20_15 = tensorLoad_io_tensor_rd_0_data_bits_20_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_21_0 = tensorLoad_io_tensor_rd_0_data_bits_21_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_21_1 = tensorLoad_io_tensor_rd_0_data_bits_21_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_21_2 = tensorLoad_io_tensor_rd_0_data_bits_21_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_21_3 = tensorLoad_io_tensor_rd_0_data_bits_21_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_21_4 = tensorLoad_io_tensor_rd_0_data_bits_21_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_21_5 = tensorLoad_io_tensor_rd_0_data_bits_21_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_21_6 = tensorLoad_io_tensor_rd_0_data_bits_21_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_21_7 = tensorLoad_io_tensor_rd_0_data_bits_21_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_21_8 = tensorLoad_io_tensor_rd_0_data_bits_21_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_21_9 = tensorLoad_io_tensor_rd_0_data_bits_21_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_21_10 = tensorLoad_io_tensor_rd_0_data_bits_21_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_21_11 = tensorLoad_io_tensor_rd_0_data_bits_21_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_21_12 = tensorLoad_io_tensor_rd_0_data_bits_21_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_21_13 = tensorLoad_io_tensor_rd_0_data_bits_21_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_21_14 = tensorLoad_io_tensor_rd_0_data_bits_21_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_21_15 = tensorLoad_io_tensor_rd_0_data_bits_21_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_22_0 = tensorLoad_io_tensor_rd_0_data_bits_22_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_22_1 = tensorLoad_io_tensor_rd_0_data_bits_22_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_22_2 = tensorLoad_io_tensor_rd_0_data_bits_22_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_22_3 = tensorLoad_io_tensor_rd_0_data_bits_22_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_22_4 = tensorLoad_io_tensor_rd_0_data_bits_22_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_22_5 = tensorLoad_io_tensor_rd_0_data_bits_22_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_22_6 = tensorLoad_io_tensor_rd_0_data_bits_22_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_22_7 = tensorLoad_io_tensor_rd_0_data_bits_22_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_22_8 = tensorLoad_io_tensor_rd_0_data_bits_22_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_22_9 = tensorLoad_io_tensor_rd_0_data_bits_22_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_22_10 = tensorLoad_io_tensor_rd_0_data_bits_22_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_22_11 = tensorLoad_io_tensor_rd_0_data_bits_22_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_22_12 = tensorLoad_io_tensor_rd_0_data_bits_22_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_22_13 = tensorLoad_io_tensor_rd_0_data_bits_22_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_22_14 = tensorLoad_io_tensor_rd_0_data_bits_22_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_22_15 = tensorLoad_io_tensor_rd_0_data_bits_22_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_23_0 = tensorLoad_io_tensor_rd_0_data_bits_23_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_23_1 = tensorLoad_io_tensor_rd_0_data_bits_23_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_23_2 = tensorLoad_io_tensor_rd_0_data_bits_23_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_23_3 = tensorLoad_io_tensor_rd_0_data_bits_23_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_23_4 = tensorLoad_io_tensor_rd_0_data_bits_23_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_23_5 = tensorLoad_io_tensor_rd_0_data_bits_23_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_23_6 = tensorLoad_io_tensor_rd_0_data_bits_23_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_23_7 = tensorLoad_io_tensor_rd_0_data_bits_23_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_23_8 = tensorLoad_io_tensor_rd_0_data_bits_23_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_23_9 = tensorLoad_io_tensor_rd_0_data_bits_23_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_23_10 = tensorLoad_io_tensor_rd_0_data_bits_23_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_23_11 = tensorLoad_io_tensor_rd_0_data_bits_23_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_23_12 = tensorLoad_io_tensor_rd_0_data_bits_23_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_23_13 = tensorLoad_io_tensor_rd_0_data_bits_23_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_23_14 = tensorLoad_io_tensor_rd_0_data_bits_23_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_23_15 = tensorLoad_io_tensor_rd_0_data_bits_23_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_24_0 = tensorLoad_io_tensor_rd_0_data_bits_24_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_24_1 = tensorLoad_io_tensor_rd_0_data_bits_24_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_24_2 = tensorLoad_io_tensor_rd_0_data_bits_24_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_24_3 = tensorLoad_io_tensor_rd_0_data_bits_24_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_24_4 = tensorLoad_io_tensor_rd_0_data_bits_24_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_24_5 = tensorLoad_io_tensor_rd_0_data_bits_24_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_24_6 = tensorLoad_io_tensor_rd_0_data_bits_24_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_24_7 = tensorLoad_io_tensor_rd_0_data_bits_24_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_24_8 = tensorLoad_io_tensor_rd_0_data_bits_24_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_24_9 = tensorLoad_io_tensor_rd_0_data_bits_24_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_24_10 = tensorLoad_io_tensor_rd_0_data_bits_24_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_24_11 = tensorLoad_io_tensor_rd_0_data_bits_24_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_24_12 = tensorLoad_io_tensor_rd_0_data_bits_24_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_24_13 = tensorLoad_io_tensor_rd_0_data_bits_24_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_24_14 = tensorLoad_io_tensor_rd_0_data_bits_24_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_24_15 = tensorLoad_io_tensor_rd_0_data_bits_24_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_25_0 = tensorLoad_io_tensor_rd_0_data_bits_25_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_25_1 = tensorLoad_io_tensor_rd_0_data_bits_25_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_25_2 = tensorLoad_io_tensor_rd_0_data_bits_25_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_25_3 = tensorLoad_io_tensor_rd_0_data_bits_25_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_25_4 = tensorLoad_io_tensor_rd_0_data_bits_25_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_25_5 = tensorLoad_io_tensor_rd_0_data_bits_25_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_25_6 = tensorLoad_io_tensor_rd_0_data_bits_25_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_25_7 = tensorLoad_io_tensor_rd_0_data_bits_25_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_25_8 = tensorLoad_io_tensor_rd_0_data_bits_25_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_25_9 = tensorLoad_io_tensor_rd_0_data_bits_25_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_25_10 = tensorLoad_io_tensor_rd_0_data_bits_25_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_25_11 = tensorLoad_io_tensor_rd_0_data_bits_25_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_25_12 = tensorLoad_io_tensor_rd_0_data_bits_25_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_25_13 = tensorLoad_io_tensor_rd_0_data_bits_25_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_25_14 = tensorLoad_io_tensor_rd_0_data_bits_25_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_25_15 = tensorLoad_io_tensor_rd_0_data_bits_25_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_26_0 = tensorLoad_io_tensor_rd_0_data_bits_26_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_26_1 = tensorLoad_io_tensor_rd_0_data_bits_26_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_26_2 = tensorLoad_io_tensor_rd_0_data_bits_26_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_26_3 = tensorLoad_io_tensor_rd_0_data_bits_26_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_26_4 = tensorLoad_io_tensor_rd_0_data_bits_26_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_26_5 = tensorLoad_io_tensor_rd_0_data_bits_26_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_26_6 = tensorLoad_io_tensor_rd_0_data_bits_26_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_26_7 = tensorLoad_io_tensor_rd_0_data_bits_26_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_26_8 = tensorLoad_io_tensor_rd_0_data_bits_26_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_26_9 = tensorLoad_io_tensor_rd_0_data_bits_26_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_26_10 = tensorLoad_io_tensor_rd_0_data_bits_26_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_26_11 = tensorLoad_io_tensor_rd_0_data_bits_26_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_26_12 = tensorLoad_io_tensor_rd_0_data_bits_26_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_26_13 = tensorLoad_io_tensor_rd_0_data_bits_26_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_26_14 = tensorLoad_io_tensor_rd_0_data_bits_26_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_26_15 = tensorLoad_io_tensor_rd_0_data_bits_26_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_27_0 = tensorLoad_io_tensor_rd_0_data_bits_27_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_27_1 = tensorLoad_io_tensor_rd_0_data_bits_27_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_27_2 = tensorLoad_io_tensor_rd_0_data_bits_27_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_27_3 = tensorLoad_io_tensor_rd_0_data_bits_27_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_27_4 = tensorLoad_io_tensor_rd_0_data_bits_27_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_27_5 = tensorLoad_io_tensor_rd_0_data_bits_27_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_27_6 = tensorLoad_io_tensor_rd_0_data_bits_27_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_27_7 = tensorLoad_io_tensor_rd_0_data_bits_27_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_27_8 = tensorLoad_io_tensor_rd_0_data_bits_27_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_27_9 = tensorLoad_io_tensor_rd_0_data_bits_27_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_27_10 = tensorLoad_io_tensor_rd_0_data_bits_27_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_27_11 = tensorLoad_io_tensor_rd_0_data_bits_27_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_27_12 = tensorLoad_io_tensor_rd_0_data_bits_27_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_27_13 = tensorLoad_io_tensor_rd_0_data_bits_27_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_27_14 = tensorLoad_io_tensor_rd_0_data_bits_27_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_27_15 = tensorLoad_io_tensor_rd_0_data_bits_27_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_28_0 = tensorLoad_io_tensor_rd_0_data_bits_28_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_28_1 = tensorLoad_io_tensor_rd_0_data_bits_28_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_28_2 = tensorLoad_io_tensor_rd_0_data_bits_28_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_28_3 = tensorLoad_io_tensor_rd_0_data_bits_28_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_28_4 = tensorLoad_io_tensor_rd_0_data_bits_28_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_28_5 = tensorLoad_io_tensor_rd_0_data_bits_28_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_28_6 = tensorLoad_io_tensor_rd_0_data_bits_28_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_28_7 = tensorLoad_io_tensor_rd_0_data_bits_28_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_28_8 = tensorLoad_io_tensor_rd_0_data_bits_28_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_28_9 = tensorLoad_io_tensor_rd_0_data_bits_28_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_28_10 = tensorLoad_io_tensor_rd_0_data_bits_28_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_28_11 = tensorLoad_io_tensor_rd_0_data_bits_28_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_28_12 = tensorLoad_io_tensor_rd_0_data_bits_28_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_28_13 = tensorLoad_io_tensor_rd_0_data_bits_28_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_28_14 = tensorLoad_io_tensor_rd_0_data_bits_28_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_28_15 = tensorLoad_io_tensor_rd_0_data_bits_28_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_29_0 = tensorLoad_io_tensor_rd_0_data_bits_29_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_29_1 = tensorLoad_io_tensor_rd_0_data_bits_29_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_29_2 = tensorLoad_io_tensor_rd_0_data_bits_29_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_29_3 = tensorLoad_io_tensor_rd_0_data_bits_29_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_29_4 = tensorLoad_io_tensor_rd_0_data_bits_29_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_29_5 = tensorLoad_io_tensor_rd_0_data_bits_29_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_29_6 = tensorLoad_io_tensor_rd_0_data_bits_29_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_29_7 = tensorLoad_io_tensor_rd_0_data_bits_29_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_29_8 = tensorLoad_io_tensor_rd_0_data_bits_29_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_29_9 = tensorLoad_io_tensor_rd_0_data_bits_29_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_29_10 = tensorLoad_io_tensor_rd_0_data_bits_29_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_29_11 = tensorLoad_io_tensor_rd_0_data_bits_29_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_29_12 = tensorLoad_io_tensor_rd_0_data_bits_29_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_29_13 = tensorLoad_io_tensor_rd_0_data_bits_29_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_29_14 = tensorLoad_io_tensor_rd_0_data_bits_29_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_29_15 = tensorLoad_io_tensor_rd_0_data_bits_29_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_30_0 = tensorLoad_io_tensor_rd_0_data_bits_30_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_30_1 = tensorLoad_io_tensor_rd_0_data_bits_30_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_30_2 = tensorLoad_io_tensor_rd_0_data_bits_30_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_30_3 = tensorLoad_io_tensor_rd_0_data_bits_30_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_30_4 = tensorLoad_io_tensor_rd_0_data_bits_30_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_30_5 = tensorLoad_io_tensor_rd_0_data_bits_30_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_30_6 = tensorLoad_io_tensor_rd_0_data_bits_30_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_30_7 = tensorLoad_io_tensor_rd_0_data_bits_30_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_30_8 = tensorLoad_io_tensor_rd_0_data_bits_30_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_30_9 = tensorLoad_io_tensor_rd_0_data_bits_30_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_30_10 = tensorLoad_io_tensor_rd_0_data_bits_30_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_30_11 = tensorLoad_io_tensor_rd_0_data_bits_30_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_30_12 = tensorLoad_io_tensor_rd_0_data_bits_30_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_30_13 = tensorLoad_io_tensor_rd_0_data_bits_30_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_30_14 = tensorLoad_io_tensor_rd_0_data_bits_30_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_30_15 = tensorLoad_io_tensor_rd_0_data_bits_30_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_31_0 = tensorLoad_io_tensor_rd_0_data_bits_31_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_31_1 = tensorLoad_io_tensor_rd_0_data_bits_31_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_31_2 = tensorLoad_io_tensor_rd_0_data_bits_31_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_31_3 = tensorLoad_io_tensor_rd_0_data_bits_31_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_31_4 = tensorLoad_io_tensor_rd_0_data_bits_31_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_31_5 = tensorLoad_io_tensor_rd_0_data_bits_31_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_31_6 = tensorLoad_io_tensor_rd_0_data_bits_31_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_31_7 = tensorLoad_io_tensor_rd_0_data_bits_31_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_31_8 = tensorLoad_io_tensor_rd_0_data_bits_31_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_31_9 = tensorLoad_io_tensor_rd_0_data_bits_31_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_31_10 = tensorLoad_io_tensor_rd_0_data_bits_31_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_31_11 = tensorLoad_io_tensor_rd_0_data_bits_31_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_31_12 = tensorLoad_io_tensor_rd_0_data_bits_31_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_31_13 = tensorLoad_io_tensor_rd_0_data_bits_31_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_31_14 = tensorLoad_io_tensor_rd_0_data_bits_31_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_31_15 = tensorLoad_io_tensor_rd_0_data_bits_31_15; // @[TensorLoad.scala 72:8]
  assign tensorLoad_clock = clock;
  assign tensorLoad_reset = reset;
  assign tensorLoad_io_start = io_start; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_inst = io_inst; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_baddr = io_baddr; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_vme_rd_cmd_ready = io_vme_rd_cmd_ready; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_vme_rd_data_valid = io_vme_rd_data_valid; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_vme_rd_data_bits_data = io_vme_rd_data_bits_data; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_vme_rd_data_bits_tag = io_vme_rd_data_bits_tag; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_rd_0_idx_valid = io_tensor_rd_0_idx_valid; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_rd_0_idx_bits = io_tensor_rd_0_idx_bits; // @[TensorLoad.scala 72:8]
endmodule
module Load(
  input          clock,
  input          reset,
  input          io_i_post,
  output         io_o_post,
  output         io_inst_ready,
  input          io_inst_valid,
  input  [127:0] io_inst_bits,
  input  [31:0]  io_inp_baddr,
  input  [31:0]  io_wgt_baddr,
  input          io_vme_rd_0_cmd_ready,
  output         io_vme_rd_0_cmd_valid,
  output [31:0]  io_vme_rd_0_cmd_bits_addr,
  output [3:0]   io_vme_rd_0_cmd_bits_len,
  output [20:0]  io_vme_rd_0_cmd_bits_tag,
  input          io_vme_rd_0_data_valid,
  input  [63:0]  io_vme_rd_0_data_bits_data,
  input  [20:0]  io_vme_rd_0_data_bits_tag,
  input          io_vme_rd_1_cmd_ready,
  output         io_vme_rd_1_cmd_valid,
  output [31:0]  io_vme_rd_1_cmd_bits_addr,
  output [3:0]   io_vme_rd_1_cmd_bits_len,
  output [20:0]  io_vme_rd_1_cmd_bits_tag,
  input          io_vme_rd_1_data_valid,
  input  [63:0]  io_vme_rd_1_data_bits_data,
  input  [20:0]  io_vme_rd_1_data_bits_tag,
  input          io_inp_rd_0_idx_valid,
  input  [6:0]   io_inp_rd_0_idx_bits,
  output         io_inp_rd_0_data_valid,
  output [7:0]   io_inp_rd_0_data_bits_0_0,
  output [7:0]   io_inp_rd_0_data_bits_0_1,
  output [7:0]   io_inp_rd_0_data_bits_0_2,
  output [7:0]   io_inp_rd_0_data_bits_0_3,
  output [7:0]   io_inp_rd_0_data_bits_0_4,
  output [7:0]   io_inp_rd_0_data_bits_0_5,
  output [7:0]   io_inp_rd_0_data_bits_0_6,
  output [7:0]   io_inp_rd_0_data_bits_0_7,
  output [7:0]   io_inp_rd_0_data_bits_0_8,
  output [7:0]   io_inp_rd_0_data_bits_0_9,
  output [7:0]   io_inp_rd_0_data_bits_0_10,
  output [7:0]   io_inp_rd_0_data_bits_0_11,
  output [7:0]   io_inp_rd_0_data_bits_0_12,
  output [7:0]   io_inp_rd_0_data_bits_0_13,
  output [7:0]   io_inp_rd_0_data_bits_0_14,
  output [7:0]   io_inp_rd_0_data_bits_0_15,
  input          io_wgt_rd_0_idx_valid,
  input  [5:0]   io_wgt_rd_0_idx_bits,
  output         io_wgt_rd_0_data_valid,
  output [7:0]   io_wgt_rd_0_data_bits_0_0,
  output [7:0]   io_wgt_rd_0_data_bits_0_1,
  output [7:0]   io_wgt_rd_0_data_bits_0_2,
  output [7:0]   io_wgt_rd_0_data_bits_0_3,
  output [7:0]   io_wgt_rd_0_data_bits_0_4,
  output [7:0]   io_wgt_rd_0_data_bits_0_5,
  output [7:0]   io_wgt_rd_0_data_bits_0_6,
  output [7:0]   io_wgt_rd_0_data_bits_0_7,
  output [7:0]   io_wgt_rd_0_data_bits_0_8,
  output [7:0]   io_wgt_rd_0_data_bits_0_9,
  output [7:0]   io_wgt_rd_0_data_bits_0_10,
  output [7:0]   io_wgt_rd_0_data_bits_0_11,
  output [7:0]   io_wgt_rd_0_data_bits_0_12,
  output [7:0]   io_wgt_rd_0_data_bits_0_13,
  output [7:0]   io_wgt_rd_0_data_bits_0_14,
  output [7:0]   io_wgt_rd_0_data_bits_0_15,
  output [7:0]   io_wgt_rd_0_data_bits_1_0,
  output [7:0]   io_wgt_rd_0_data_bits_1_1,
  output [7:0]   io_wgt_rd_0_data_bits_1_2,
  output [7:0]   io_wgt_rd_0_data_bits_1_3,
  output [7:0]   io_wgt_rd_0_data_bits_1_4,
  output [7:0]   io_wgt_rd_0_data_bits_1_5,
  output [7:0]   io_wgt_rd_0_data_bits_1_6,
  output [7:0]   io_wgt_rd_0_data_bits_1_7,
  output [7:0]   io_wgt_rd_0_data_bits_1_8,
  output [7:0]   io_wgt_rd_0_data_bits_1_9,
  output [7:0]   io_wgt_rd_0_data_bits_1_10,
  output [7:0]   io_wgt_rd_0_data_bits_1_11,
  output [7:0]   io_wgt_rd_0_data_bits_1_12,
  output [7:0]   io_wgt_rd_0_data_bits_1_13,
  output [7:0]   io_wgt_rd_0_data_bits_1_14,
  output [7:0]   io_wgt_rd_0_data_bits_1_15,
  output [7:0]   io_wgt_rd_0_data_bits_2_0,
  output [7:0]   io_wgt_rd_0_data_bits_2_1,
  output [7:0]   io_wgt_rd_0_data_bits_2_2,
  output [7:0]   io_wgt_rd_0_data_bits_2_3,
  output [7:0]   io_wgt_rd_0_data_bits_2_4,
  output [7:0]   io_wgt_rd_0_data_bits_2_5,
  output [7:0]   io_wgt_rd_0_data_bits_2_6,
  output [7:0]   io_wgt_rd_0_data_bits_2_7,
  output [7:0]   io_wgt_rd_0_data_bits_2_8,
  output [7:0]   io_wgt_rd_0_data_bits_2_9,
  output [7:0]   io_wgt_rd_0_data_bits_2_10,
  output [7:0]   io_wgt_rd_0_data_bits_2_11,
  output [7:0]   io_wgt_rd_0_data_bits_2_12,
  output [7:0]   io_wgt_rd_0_data_bits_2_13,
  output [7:0]   io_wgt_rd_0_data_bits_2_14,
  output [7:0]   io_wgt_rd_0_data_bits_2_15,
  output [7:0]   io_wgt_rd_0_data_bits_3_0,
  output [7:0]   io_wgt_rd_0_data_bits_3_1,
  output [7:0]   io_wgt_rd_0_data_bits_3_2,
  output [7:0]   io_wgt_rd_0_data_bits_3_3,
  output [7:0]   io_wgt_rd_0_data_bits_3_4,
  output [7:0]   io_wgt_rd_0_data_bits_3_5,
  output [7:0]   io_wgt_rd_0_data_bits_3_6,
  output [7:0]   io_wgt_rd_0_data_bits_3_7,
  output [7:0]   io_wgt_rd_0_data_bits_3_8,
  output [7:0]   io_wgt_rd_0_data_bits_3_9,
  output [7:0]   io_wgt_rd_0_data_bits_3_10,
  output [7:0]   io_wgt_rd_0_data_bits_3_11,
  output [7:0]   io_wgt_rd_0_data_bits_3_12,
  output [7:0]   io_wgt_rd_0_data_bits_3_13,
  output [7:0]   io_wgt_rd_0_data_bits_3_14,
  output [7:0]   io_wgt_rd_0_data_bits_3_15,
  output [7:0]   io_wgt_rd_0_data_bits_4_0,
  output [7:0]   io_wgt_rd_0_data_bits_4_1,
  output [7:0]   io_wgt_rd_0_data_bits_4_2,
  output [7:0]   io_wgt_rd_0_data_bits_4_3,
  output [7:0]   io_wgt_rd_0_data_bits_4_4,
  output [7:0]   io_wgt_rd_0_data_bits_4_5,
  output [7:0]   io_wgt_rd_0_data_bits_4_6,
  output [7:0]   io_wgt_rd_0_data_bits_4_7,
  output [7:0]   io_wgt_rd_0_data_bits_4_8,
  output [7:0]   io_wgt_rd_0_data_bits_4_9,
  output [7:0]   io_wgt_rd_0_data_bits_4_10,
  output [7:0]   io_wgt_rd_0_data_bits_4_11,
  output [7:0]   io_wgt_rd_0_data_bits_4_12,
  output [7:0]   io_wgt_rd_0_data_bits_4_13,
  output [7:0]   io_wgt_rd_0_data_bits_4_14,
  output [7:0]   io_wgt_rd_0_data_bits_4_15,
  output [7:0]   io_wgt_rd_0_data_bits_5_0,
  output [7:0]   io_wgt_rd_0_data_bits_5_1,
  output [7:0]   io_wgt_rd_0_data_bits_5_2,
  output [7:0]   io_wgt_rd_0_data_bits_5_3,
  output [7:0]   io_wgt_rd_0_data_bits_5_4,
  output [7:0]   io_wgt_rd_0_data_bits_5_5,
  output [7:0]   io_wgt_rd_0_data_bits_5_6,
  output [7:0]   io_wgt_rd_0_data_bits_5_7,
  output [7:0]   io_wgt_rd_0_data_bits_5_8,
  output [7:0]   io_wgt_rd_0_data_bits_5_9,
  output [7:0]   io_wgt_rd_0_data_bits_5_10,
  output [7:0]   io_wgt_rd_0_data_bits_5_11,
  output [7:0]   io_wgt_rd_0_data_bits_5_12,
  output [7:0]   io_wgt_rd_0_data_bits_5_13,
  output [7:0]   io_wgt_rd_0_data_bits_5_14,
  output [7:0]   io_wgt_rd_0_data_bits_5_15,
  output [7:0]   io_wgt_rd_0_data_bits_6_0,
  output [7:0]   io_wgt_rd_0_data_bits_6_1,
  output [7:0]   io_wgt_rd_0_data_bits_6_2,
  output [7:0]   io_wgt_rd_0_data_bits_6_3,
  output [7:0]   io_wgt_rd_0_data_bits_6_4,
  output [7:0]   io_wgt_rd_0_data_bits_6_5,
  output [7:0]   io_wgt_rd_0_data_bits_6_6,
  output [7:0]   io_wgt_rd_0_data_bits_6_7,
  output [7:0]   io_wgt_rd_0_data_bits_6_8,
  output [7:0]   io_wgt_rd_0_data_bits_6_9,
  output [7:0]   io_wgt_rd_0_data_bits_6_10,
  output [7:0]   io_wgt_rd_0_data_bits_6_11,
  output [7:0]   io_wgt_rd_0_data_bits_6_12,
  output [7:0]   io_wgt_rd_0_data_bits_6_13,
  output [7:0]   io_wgt_rd_0_data_bits_6_14,
  output [7:0]   io_wgt_rd_0_data_bits_6_15,
  output [7:0]   io_wgt_rd_0_data_bits_7_0,
  output [7:0]   io_wgt_rd_0_data_bits_7_1,
  output [7:0]   io_wgt_rd_0_data_bits_7_2,
  output [7:0]   io_wgt_rd_0_data_bits_7_3,
  output [7:0]   io_wgt_rd_0_data_bits_7_4,
  output [7:0]   io_wgt_rd_0_data_bits_7_5,
  output [7:0]   io_wgt_rd_0_data_bits_7_6,
  output [7:0]   io_wgt_rd_0_data_bits_7_7,
  output [7:0]   io_wgt_rd_0_data_bits_7_8,
  output [7:0]   io_wgt_rd_0_data_bits_7_9,
  output [7:0]   io_wgt_rd_0_data_bits_7_10,
  output [7:0]   io_wgt_rd_0_data_bits_7_11,
  output [7:0]   io_wgt_rd_0_data_bits_7_12,
  output [7:0]   io_wgt_rd_0_data_bits_7_13,
  output [7:0]   io_wgt_rd_0_data_bits_7_14,
  output [7:0]   io_wgt_rd_0_data_bits_7_15,
  output [7:0]   io_wgt_rd_0_data_bits_8_0,
  output [7:0]   io_wgt_rd_0_data_bits_8_1,
  output [7:0]   io_wgt_rd_0_data_bits_8_2,
  output [7:0]   io_wgt_rd_0_data_bits_8_3,
  output [7:0]   io_wgt_rd_0_data_bits_8_4,
  output [7:0]   io_wgt_rd_0_data_bits_8_5,
  output [7:0]   io_wgt_rd_0_data_bits_8_6,
  output [7:0]   io_wgt_rd_0_data_bits_8_7,
  output [7:0]   io_wgt_rd_0_data_bits_8_8,
  output [7:0]   io_wgt_rd_0_data_bits_8_9,
  output [7:0]   io_wgt_rd_0_data_bits_8_10,
  output [7:0]   io_wgt_rd_0_data_bits_8_11,
  output [7:0]   io_wgt_rd_0_data_bits_8_12,
  output [7:0]   io_wgt_rd_0_data_bits_8_13,
  output [7:0]   io_wgt_rd_0_data_bits_8_14,
  output [7:0]   io_wgt_rd_0_data_bits_8_15,
  output [7:0]   io_wgt_rd_0_data_bits_9_0,
  output [7:0]   io_wgt_rd_0_data_bits_9_1,
  output [7:0]   io_wgt_rd_0_data_bits_9_2,
  output [7:0]   io_wgt_rd_0_data_bits_9_3,
  output [7:0]   io_wgt_rd_0_data_bits_9_4,
  output [7:0]   io_wgt_rd_0_data_bits_9_5,
  output [7:0]   io_wgt_rd_0_data_bits_9_6,
  output [7:0]   io_wgt_rd_0_data_bits_9_7,
  output [7:0]   io_wgt_rd_0_data_bits_9_8,
  output [7:0]   io_wgt_rd_0_data_bits_9_9,
  output [7:0]   io_wgt_rd_0_data_bits_9_10,
  output [7:0]   io_wgt_rd_0_data_bits_9_11,
  output [7:0]   io_wgt_rd_0_data_bits_9_12,
  output [7:0]   io_wgt_rd_0_data_bits_9_13,
  output [7:0]   io_wgt_rd_0_data_bits_9_14,
  output [7:0]   io_wgt_rd_0_data_bits_9_15,
  output [7:0]   io_wgt_rd_0_data_bits_10_0,
  output [7:0]   io_wgt_rd_0_data_bits_10_1,
  output [7:0]   io_wgt_rd_0_data_bits_10_2,
  output [7:0]   io_wgt_rd_0_data_bits_10_3,
  output [7:0]   io_wgt_rd_0_data_bits_10_4,
  output [7:0]   io_wgt_rd_0_data_bits_10_5,
  output [7:0]   io_wgt_rd_0_data_bits_10_6,
  output [7:0]   io_wgt_rd_0_data_bits_10_7,
  output [7:0]   io_wgt_rd_0_data_bits_10_8,
  output [7:0]   io_wgt_rd_0_data_bits_10_9,
  output [7:0]   io_wgt_rd_0_data_bits_10_10,
  output [7:0]   io_wgt_rd_0_data_bits_10_11,
  output [7:0]   io_wgt_rd_0_data_bits_10_12,
  output [7:0]   io_wgt_rd_0_data_bits_10_13,
  output [7:0]   io_wgt_rd_0_data_bits_10_14,
  output [7:0]   io_wgt_rd_0_data_bits_10_15,
  output [7:0]   io_wgt_rd_0_data_bits_11_0,
  output [7:0]   io_wgt_rd_0_data_bits_11_1,
  output [7:0]   io_wgt_rd_0_data_bits_11_2,
  output [7:0]   io_wgt_rd_0_data_bits_11_3,
  output [7:0]   io_wgt_rd_0_data_bits_11_4,
  output [7:0]   io_wgt_rd_0_data_bits_11_5,
  output [7:0]   io_wgt_rd_0_data_bits_11_6,
  output [7:0]   io_wgt_rd_0_data_bits_11_7,
  output [7:0]   io_wgt_rd_0_data_bits_11_8,
  output [7:0]   io_wgt_rd_0_data_bits_11_9,
  output [7:0]   io_wgt_rd_0_data_bits_11_10,
  output [7:0]   io_wgt_rd_0_data_bits_11_11,
  output [7:0]   io_wgt_rd_0_data_bits_11_12,
  output [7:0]   io_wgt_rd_0_data_bits_11_13,
  output [7:0]   io_wgt_rd_0_data_bits_11_14,
  output [7:0]   io_wgt_rd_0_data_bits_11_15,
  output [7:0]   io_wgt_rd_0_data_bits_12_0,
  output [7:0]   io_wgt_rd_0_data_bits_12_1,
  output [7:0]   io_wgt_rd_0_data_bits_12_2,
  output [7:0]   io_wgt_rd_0_data_bits_12_3,
  output [7:0]   io_wgt_rd_0_data_bits_12_4,
  output [7:0]   io_wgt_rd_0_data_bits_12_5,
  output [7:0]   io_wgt_rd_0_data_bits_12_6,
  output [7:0]   io_wgt_rd_0_data_bits_12_7,
  output [7:0]   io_wgt_rd_0_data_bits_12_8,
  output [7:0]   io_wgt_rd_0_data_bits_12_9,
  output [7:0]   io_wgt_rd_0_data_bits_12_10,
  output [7:0]   io_wgt_rd_0_data_bits_12_11,
  output [7:0]   io_wgt_rd_0_data_bits_12_12,
  output [7:0]   io_wgt_rd_0_data_bits_12_13,
  output [7:0]   io_wgt_rd_0_data_bits_12_14,
  output [7:0]   io_wgt_rd_0_data_bits_12_15,
  output [7:0]   io_wgt_rd_0_data_bits_13_0,
  output [7:0]   io_wgt_rd_0_data_bits_13_1,
  output [7:0]   io_wgt_rd_0_data_bits_13_2,
  output [7:0]   io_wgt_rd_0_data_bits_13_3,
  output [7:0]   io_wgt_rd_0_data_bits_13_4,
  output [7:0]   io_wgt_rd_0_data_bits_13_5,
  output [7:0]   io_wgt_rd_0_data_bits_13_6,
  output [7:0]   io_wgt_rd_0_data_bits_13_7,
  output [7:0]   io_wgt_rd_0_data_bits_13_8,
  output [7:0]   io_wgt_rd_0_data_bits_13_9,
  output [7:0]   io_wgt_rd_0_data_bits_13_10,
  output [7:0]   io_wgt_rd_0_data_bits_13_11,
  output [7:0]   io_wgt_rd_0_data_bits_13_12,
  output [7:0]   io_wgt_rd_0_data_bits_13_13,
  output [7:0]   io_wgt_rd_0_data_bits_13_14,
  output [7:0]   io_wgt_rd_0_data_bits_13_15,
  output [7:0]   io_wgt_rd_0_data_bits_14_0,
  output [7:0]   io_wgt_rd_0_data_bits_14_1,
  output [7:0]   io_wgt_rd_0_data_bits_14_2,
  output [7:0]   io_wgt_rd_0_data_bits_14_3,
  output [7:0]   io_wgt_rd_0_data_bits_14_4,
  output [7:0]   io_wgt_rd_0_data_bits_14_5,
  output [7:0]   io_wgt_rd_0_data_bits_14_6,
  output [7:0]   io_wgt_rd_0_data_bits_14_7,
  output [7:0]   io_wgt_rd_0_data_bits_14_8,
  output [7:0]   io_wgt_rd_0_data_bits_14_9,
  output [7:0]   io_wgt_rd_0_data_bits_14_10,
  output [7:0]   io_wgt_rd_0_data_bits_14_11,
  output [7:0]   io_wgt_rd_0_data_bits_14_12,
  output [7:0]   io_wgt_rd_0_data_bits_14_13,
  output [7:0]   io_wgt_rd_0_data_bits_14_14,
  output [7:0]   io_wgt_rd_0_data_bits_14_15,
  output [7:0]   io_wgt_rd_0_data_bits_15_0,
  output [7:0]   io_wgt_rd_0_data_bits_15_1,
  output [7:0]   io_wgt_rd_0_data_bits_15_2,
  output [7:0]   io_wgt_rd_0_data_bits_15_3,
  output [7:0]   io_wgt_rd_0_data_bits_15_4,
  output [7:0]   io_wgt_rd_0_data_bits_15_5,
  output [7:0]   io_wgt_rd_0_data_bits_15_6,
  output [7:0]   io_wgt_rd_0_data_bits_15_7,
  output [7:0]   io_wgt_rd_0_data_bits_15_8,
  output [7:0]   io_wgt_rd_0_data_bits_15_9,
  output [7:0]   io_wgt_rd_0_data_bits_15_10,
  output [7:0]   io_wgt_rd_0_data_bits_15_11,
  output [7:0]   io_wgt_rd_0_data_bits_15_12,
  output [7:0]   io_wgt_rd_0_data_bits_15_13,
  output [7:0]   io_wgt_rd_0_data_bits_15_14,
  output [7:0]   io_wgt_rd_0_data_bits_15_15,
  output [7:0]   io_wgt_rd_0_data_bits_16_0,
  output [7:0]   io_wgt_rd_0_data_bits_16_1,
  output [7:0]   io_wgt_rd_0_data_bits_16_2,
  output [7:0]   io_wgt_rd_0_data_bits_16_3,
  output [7:0]   io_wgt_rd_0_data_bits_16_4,
  output [7:0]   io_wgt_rd_0_data_bits_16_5,
  output [7:0]   io_wgt_rd_0_data_bits_16_6,
  output [7:0]   io_wgt_rd_0_data_bits_16_7,
  output [7:0]   io_wgt_rd_0_data_bits_16_8,
  output [7:0]   io_wgt_rd_0_data_bits_16_9,
  output [7:0]   io_wgt_rd_0_data_bits_16_10,
  output [7:0]   io_wgt_rd_0_data_bits_16_11,
  output [7:0]   io_wgt_rd_0_data_bits_16_12,
  output [7:0]   io_wgt_rd_0_data_bits_16_13,
  output [7:0]   io_wgt_rd_0_data_bits_16_14,
  output [7:0]   io_wgt_rd_0_data_bits_16_15,
  output [7:0]   io_wgt_rd_0_data_bits_17_0,
  output [7:0]   io_wgt_rd_0_data_bits_17_1,
  output [7:0]   io_wgt_rd_0_data_bits_17_2,
  output [7:0]   io_wgt_rd_0_data_bits_17_3,
  output [7:0]   io_wgt_rd_0_data_bits_17_4,
  output [7:0]   io_wgt_rd_0_data_bits_17_5,
  output [7:0]   io_wgt_rd_0_data_bits_17_6,
  output [7:0]   io_wgt_rd_0_data_bits_17_7,
  output [7:0]   io_wgt_rd_0_data_bits_17_8,
  output [7:0]   io_wgt_rd_0_data_bits_17_9,
  output [7:0]   io_wgt_rd_0_data_bits_17_10,
  output [7:0]   io_wgt_rd_0_data_bits_17_11,
  output [7:0]   io_wgt_rd_0_data_bits_17_12,
  output [7:0]   io_wgt_rd_0_data_bits_17_13,
  output [7:0]   io_wgt_rd_0_data_bits_17_14,
  output [7:0]   io_wgt_rd_0_data_bits_17_15,
  output [7:0]   io_wgt_rd_0_data_bits_18_0,
  output [7:0]   io_wgt_rd_0_data_bits_18_1,
  output [7:0]   io_wgt_rd_0_data_bits_18_2,
  output [7:0]   io_wgt_rd_0_data_bits_18_3,
  output [7:0]   io_wgt_rd_0_data_bits_18_4,
  output [7:0]   io_wgt_rd_0_data_bits_18_5,
  output [7:0]   io_wgt_rd_0_data_bits_18_6,
  output [7:0]   io_wgt_rd_0_data_bits_18_7,
  output [7:0]   io_wgt_rd_0_data_bits_18_8,
  output [7:0]   io_wgt_rd_0_data_bits_18_9,
  output [7:0]   io_wgt_rd_0_data_bits_18_10,
  output [7:0]   io_wgt_rd_0_data_bits_18_11,
  output [7:0]   io_wgt_rd_0_data_bits_18_12,
  output [7:0]   io_wgt_rd_0_data_bits_18_13,
  output [7:0]   io_wgt_rd_0_data_bits_18_14,
  output [7:0]   io_wgt_rd_0_data_bits_18_15,
  output [7:0]   io_wgt_rd_0_data_bits_19_0,
  output [7:0]   io_wgt_rd_0_data_bits_19_1,
  output [7:0]   io_wgt_rd_0_data_bits_19_2,
  output [7:0]   io_wgt_rd_0_data_bits_19_3,
  output [7:0]   io_wgt_rd_0_data_bits_19_4,
  output [7:0]   io_wgt_rd_0_data_bits_19_5,
  output [7:0]   io_wgt_rd_0_data_bits_19_6,
  output [7:0]   io_wgt_rd_0_data_bits_19_7,
  output [7:0]   io_wgt_rd_0_data_bits_19_8,
  output [7:0]   io_wgt_rd_0_data_bits_19_9,
  output [7:0]   io_wgt_rd_0_data_bits_19_10,
  output [7:0]   io_wgt_rd_0_data_bits_19_11,
  output [7:0]   io_wgt_rd_0_data_bits_19_12,
  output [7:0]   io_wgt_rd_0_data_bits_19_13,
  output [7:0]   io_wgt_rd_0_data_bits_19_14,
  output [7:0]   io_wgt_rd_0_data_bits_19_15,
  output [7:0]   io_wgt_rd_0_data_bits_20_0,
  output [7:0]   io_wgt_rd_0_data_bits_20_1,
  output [7:0]   io_wgt_rd_0_data_bits_20_2,
  output [7:0]   io_wgt_rd_0_data_bits_20_3,
  output [7:0]   io_wgt_rd_0_data_bits_20_4,
  output [7:0]   io_wgt_rd_0_data_bits_20_5,
  output [7:0]   io_wgt_rd_0_data_bits_20_6,
  output [7:0]   io_wgt_rd_0_data_bits_20_7,
  output [7:0]   io_wgt_rd_0_data_bits_20_8,
  output [7:0]   io_wgt_rd_0_data_bits_20_9,
  output [7:0]   io_wgt_rd_0_data_bits_20_10,
  output [7:0]   io_wgt_rd_0_data_bits_20_11,
  output [7:0]   io_wgt_rd_0_data_bits_20_12,
  output [7:0]   io_wgt_rd_0_data_bits_20_13,
  output [7:0]   io_wgt_rd_0_data_bits_20_14,
  output [7:0]   io_wgt_rd_0_data_bits_20_15,
  output [7:0]   io_wgt_rd_0_data_bits_21_0,
  output [7:0]   io_wgt_rd_0_data_bits_21_1,
  output [7:0]   io_wgt_rd_0_data_bits_21_2,
  output [7:0]   io_wgt_rd_0_data_bits_21_3,
  output [7:0]   io_wgt_rd_0_data_bits_21_4,
  output [7:0]   io_wgt_rd_0_data_bits_21_5,
  output [7:0]   io_wgt_rd_0_data_bits_21_6,
  output [7:0]   io_wgt_rd_0_data_bits_21_7,
  output [7:0]   io_wgt_rd_0_data_bits_21_8,
  output [7:0]   io_wgt_rd_0_data_bits_21_9,
  output [7:0]   io_wgt_rd_0_data_bits_21_10,
  output [7:0]   io_wgt_rd_0_data_bits_21_11,
  output [7:0]   io_wgt_rd_0_data_bits_21_12,
  output [7:0]   io_wgt_rd_0_data_bits_21_13,
  output [7:0]   io_wgt_rd_0_data_bits_21_14,
  output [7:0]   io_wgt_rd_0_data_bits_21_15,
  output [7:0]   io_wgt_rd_0_data_bits_22_0,
  output [7:0]   io_wgt_rd_0_data_bits_22_1,
  output [7:0]   io_wgt_rd_0_data_bits_22_2,
  output [7:0]   io_wgt_rd_0_data_bits_22_3,
  output [7:0]   io_wgt_rd_0_data_bits_22_4,
  output [7:0]   io_wgt_rd_0_data_bits_22_5,
  output [7:0]   io_wgt_rd_0_data_bits_22_6,
  output [7:0]   io_wgt_rd_0_data_bits_22_7,
  output [7:0]   io_wgt_rd_0_data_bits_22_8,
  output [7:0]   io_wgt_rd_0_data_bits_22_9,
  output [7:0]   io_wgt_rd_0_data_bits_22_10,
  output [7:0]   io_wgt_rd_0_data_bits_22_11,
  output [7:0]   io_wgt_rd_0_data_bits_22_12,
  output [7:0]   io_wgt_rd_0_data_bits_22_13,
  output [7:0]   io_wgt_rd_0_data_bits_22_14,
  output [7:0]   io_wgt_rd_0_data_bits_22_15,
  output [7:0]   io_wgt_rd_0_data_bits_23_0,
  output [7:0]   io_wgt_rd_0_data_bits_23_1,
  output [7:0]   io_wgt_rd_0_data_bits_23_2,
  output [7:0]   io_wgt_rd_0_data_bits_23_3,
  output [7:0]   io_wgt_rd_0_data_bits_23_4,
  output [7:0]   io_wgt_rd_0_data_bits_23_5,
  output [7:0]   io_wgt_rd_0_data_bits_23_6,
  output [7:0]   io_wgt_rd_0_data_bits_23_7,
  output [7:0]   io_wgt_rd_0_data_bits_23_8,
  output [7:0]   io_wgt_rd_0_data_bits_23_9,
  output [7:0]   io_wgt_rd_0_data_bits_23_10,
  output [7:0]   io_wgt_rd_0_data_bits_23_11,
  output [7:0]   io_wgt_rd_0_data_bits_23_12,
  output [7:0]   io_wgt_rd_0_data_bits_23_13,
  output [7:0]   io_wgt_rd_0_data_bits_23_14,
  output [7:0]   io_wgt_rd_0_data_bits_23_15,
  output [7:0]   io_wgt_rd_0_data_bits_24_0,
  output [7:0]   io_wgt_rd_0_data_bits_24_1,
  output [7:0]   io_wgt_rd_0_data_bits_24_2,
  output [7:0]   io_wgt_rd_0_data_bits_24_3,
  output [7:0]   io_wgt_rd_0_data_bits_24_4,
  output [7:0]   io_wgt_rd_0_data_bits_24_5,
  output [7:0]   io_wgt_rd_0_data_bits_24_6,
  output [7:0]   io_wgt_rd_0_data_bits_24_7,
  output [7:0]   io_wgt_rd_0_data_bits_24_8,
  output [7:0]   io_wgt_rd_0_data_bits_24_9,
  output [7:0]   io_wgt_rd_0_data_bits_24_10,
  output [7:0]   io_wgt_rd_0_data_bits_24_11,
  output [7:0]   io_wgt_rd_0_data_bits_24_12,
  output [7:0]   io_wgt_rd_0_data_bits_24_13,
  output [7:0]   io_wgt_rd_0_data_bits_24_14,
  output [7:0]   io_wgt_rd_0_data_bits_24_15,
  output [7:0]   io_wgt_rd_0_data_bits_25_0,
  output [7:0]   io_wgt_rd_0_data_bits_25_1,
  output [7:0]   io_wgt_rd_0_data_bits_25_2,
  output [7:0]   io_wgt_rd_0_data_bits_25_3,
  output [7:0]   io_wgt_rd_0_data_bits_25_4,
  output [7:0]   io_wgt_rd_0_data_bits_25_5,
  output [7:0]   io_wgt_rd_0_data_bits_25_6,
  output [7:0]   io_wgt_rd_0_data_bits_25_7,
  output [7:0]   io_wgt_rd_0_data_bits_25_8,
  output [7:0]   io_wgt_rd_0_data_bits_25_9,
  output [7:0]   io_wgt_rd_0_data_bits_25_10,
  output [7:0]   io_wgt_rd_0_data_bits_25_11,
  output [7:0]   io_wgt_rd_0_data_bits_25_12,
  output [7:0]   io_wgt_rd_0_data_bits_25_13,
  output [7:0]   io_wgt_rd_0_data_bits_25_14,
  output [7:0]   io_wgt_rd_0_data_bits_25_15,
  output [7:0]   io_wgt_rd_0_data_bits_26_0,
  output [7:0]   io_wgt_rd_0_data_bits_26_1,
  output [7:0]   io_wgt_rd_0_data_bits_26_2,
  output [7:0]   io_wgt_rd_0_data_bits_26_3,
  output [7:0]   io_wgt_rd_0_data_bits_26_4,
  output [7:0]   io_wgt_rd_0_data_bits_26_5,
  output [7:0]   io_wgt_rd_0_data_bits_26_6,
  output [7:0]   io_wgt_rd_0_data_bits_26_7,
  output [7:0]   io_wgt_rd_0_data_bits_26_8,
  output [7:0]   io_wgt_rd_0_data_bits_26_9,
  output [7:0]   io_wgt_rd_0_data_bits_26_10,
  output [7:0]   io_wgt_rd_0_data_bits_26_11,
  output [7:0]   io_wgt_rd_0_data_bits_26_12,
  output [7:0]   io_wgt_rd_0_data_bits_26_13,
  output [7:0]   io_wgt_rd_0_data_bits_26_14,
  output [7:0]   io_wgt_rd_0_data_bits_26_15,
  output [7:0]   io_wgt_rd_0_data_bits_27_0,
  output [7:0]   io_wgt_rd_0_data_bits_27_1,
  output [7:0]   io_wgt_rd_0_data_bits_27_2,
  output [7:0]   io_wgt_rd_0_data_bits_27_3,
  output [7:0]   io_wgt_rd_0_data_bits_27_4,
  output [7:0]   io_wgt_rd_0_data_bits_27_5,
  output [7:0]   io_wgt_rd_0_data_bits_27_6,
  output [7:0]   io_wgt_rd_0_data_bits_27_7,
  output [7:0]   io_wgt_rd_0_data_bits_27_8,
  output [7:0]   io_wgt_rd_0_data_bits_27_9,
  output [7:0]   io_wgt_rd_0_data_bits_27_10,
  output [7:0]   io_wgt_rd_0_data_bits_27_11,
  output [7:0]   io_wgt_rd_0_data_bits_27_12,
  output [7:0]   io_wgt_rd_0_data_bits_27_13,
  output [7:0]   io_wgt_rd_0_data_bits_27_14,
  output [7:0]   io_wgt_rd_0_data_bits_27_15,
  output [7:0]   io_wgt_rd_0_data_bits_28_0,
  output [7:0]   io_wgt_rd_0_data_bits_28_1,
  output [7:0]   io_wgt_rd_0_data_bits_28_2,
  output [7:0]   io_wgt_rd_0_data_bits_28_3,
  output [7:0]   io_wgt_rd_0_data_bits_28_4,
  output [7:0]   io_wgt_rd_0_data_bits_28_5,
  output [7:0]   io_wgt_rd_0_data_bits_28_6,
  output [7:0]   io_wgt_rd_0_data_bits_28_7,
  output [7:0]   io_wgt_rd_0_data_bits_28_8,
  output [7:0]   io_wgt_rd_0_data_bits_28_9,
  output [7:0]   io_wgt_rd_0_data_bits_28_10,
  output [7:0]   io_wgt_rd_0_data_bits_28_11,
  output [7:0]   io_wgt_rd_0_data_bits_28_12,
  output [7:0]   io_wgt_rd_0_data_bits_28_13,
  output [7:0]   io_wgt_rd_0_data_bits_28_14,
  output [7:0]   io_wgt_rd_0_data_bits_28_15,
  output [7:0]   io_wgt_rd_0_data_bits_29_0,
  output [7:0]   io_wgt_rd_0_data_bits_29_1,
  output [7:0]   io_wgt_rd_0_data_bits_29_2,
  output [7:0]   io_wgt_rd_0_data_bits_29_3,
  output [7:0]   io_wgt_rd_0_data_bits_29_4,
  output [7:0]   io_wgt_rd_0_data_bits_29_5,
  output [7:0]   io_wgt_rd_0_data_bits_29_6,
  output [7:0]   io_wgt_rd_0_data_bits_29_7,
  output [7:0]   io_wgt_rd_0_data_bits_29_8,
  output [7:0]   io_wgt_rd_0_data_bits_29_9,
  output [7:0]   io_wgt_rd_0_data_bits_29_10,
  output [7:0]   io_wgt_rd_0_data_bits_29_11,
  output [7:0]   io_wgt_rd_0_data_bits_29_12,
  output [7:0]   io_wgt_rd_0_data_bits_29_13,
  output [7:0]   io_wgt_rd_0_data_bits_29_14,
  output [7:0]   io_wgt_rd_0_data_bits_29_15,
  output [7:0]   io_wgt_rd_0_data_bits_30_0,
  output [7:0]   io_wgt_rd_0_data_bits_30_1,
  output [7:0]   io_wgt_rd_0_data_bits_30_2,
  output [7:0]   io_wgt_rd_0_data_bits_30_3,
  output [7:0]   io_wgt_rd_0_data_bits_30_4,
  output [7:0]   io_wgt_rd_0_data_bits_30_5,
  output [7:0]   io_wgt_rd_0_data_bits_30_6,
  output [7:0]   io_wgt_rd_0_data_bits_30_7,
  output [7:0]   io_wgt_rd_0_data_bits_30_8,
  output [7:0]   io_wgt_rd_0_data_bits_30_9,
  output [7:0]   io_wgt_rd_0_data_bits_30_10,
  output [7:0]   io_wgt_rd_0_data_bits_30_11,
  output [7:0]   io_wgt_rd_0_data_bits_30_12,
  output [7:0]   io_wgt_rd_0_data_bits_30_13,
  output [7:0]   io_wgt_rd_0_data_bits_30_14,
  output [7:0]   io_wgt_rd_0_data_bits_30_15,
  output [7:0]   io_wgt_rd_0_data_bits_31_0,
  output [7:0]   io_wgt_rd_0_data_bits_31_1,
  output [7:0]   io_wgt_rd_0_data_bits_31_2,
  output [7:0]   io_wgt_rd_0_data_bits_31_3,
  output [7:0]   io_wgt_rd_0_data_bits_31_4,
  output [7:0]   io_wgt_rd_0_data_bits_31_5,
  output [7:0]   io_wgt_rd_0_data_bits_31_6,
  output [7:0]   io_wgt_rd_0_data_bits_31_7,
  output [7:0]   io_wgt_rd_0_data_bits_31_8,
  output [7:0]   io_wgt_rd_0_data_bits_31_9,
  output [7:0]   io_wgt_rd_0_data_bits_31_10,
  output [7:0]   io_wgt_rd_0_data_bits_31_11,
  output [7:0]   io_wgt_rd_0_data_bits_31_12,
  output [7:0]   io_wgt_rd_0_data_bits_31_13,
  output [7:0]   io_wgt_rd_0_data_bits_31_14,
  output [7:0]   io_wgt_rd_0_data_bits_31_15
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  s_clock; // @[Load.scala 49:17]
  wire  s_reset; // @[Load.scala 49:17]
  wire  s_io_spost; // @[Load.scala 49:17]
  wire  s_io_swait; // @[Load.scala 49:17]
  wire  s_io_sready; // @[Load.scala 49:17]
  wire  inst_q_clock; // @[Load.scala 50:22]
  wire  inst_q_reset; // @[Load.scala 50:22]
  wire  inst_q_io_enq_ready; // @[Load.scala 50:22]
  wire  inst_q_io_enq_valid; // @[Load.scala 50:22]
  wire [127:0] inst_q_io_enq_bits; // @[Load.scala 50:22]
  wire  inst_q_io_deq_ready; // @[Load.scala 50:22]
  wire  inst_q_io_deq_valid; // @[Load.scala 50:22]
  wire [127:0] inst_q_io_deq_bits; // @[Load.scala 50:22]
  wire [127:0] dec_io_inst; // @[Load.scala 52:19]
  wire  dec_io_push_next; // @[Load.scala 52:19]
  wire  dec_io_pop_next; // @[Load.scala 52:19]
  wire  dec_io_isInput; // @[Load.scala 52:19]
  wire  dec_io_isWeight; // @[Load.scala 52:19]
  wire  dec_io_isSync; // @[Load.scala 52:19]
  wire  tensorLoad_0_clock; // @[Load.scala 58:32]
  wire  tensorLoad_0_reset; // @[Load.scala 58:32]
  wire  tensorLoad_0_io_start; // @[Load.scala 58:32]
  wire  tensorLoad_0_io_done; // @[Load.scala 58:32]
  wire [127:0] tensorLoad_0_io_inst; // @[Load.scala 58:32]
  wire [31:0] tensorLoad_0_io_baddr; // @[Load.scala 58:32]
  wire  tensorLoad_0_io_vme_rd_cmd_ready; // @[Load.scala 58:32]
  wire  tensorLoad_0_io_vme_rd_cmd_valid; // @[Load.scala 58:32]
  wire [31:0] tensorLoad_0_io_vme_rd_cmd_bits_addr; // @[Load.scala 58:32]
  wire [3:0] tensorLoad_0_io_vme_rd_cmd_bits_len; // @[Load.scala 58:32]
  wire [20:0] tensorLoad_0_io_vme_rd_cmd_bits_tag; // @[Load.scala 58:32]
  wire  tensorLoad_0_io_vme_rd_data_valid; // @[Load.scala 58:32]
  wire [63:0] tensorLoad_0_io_vme_rd_data_bits_data; // @[Load.scala 58:32]
  wire [20:0] tensorLoad_0_io_vme_rd_data_bits_tag; // @[Load.scala 58:32]
  wire  tensorLoad_0_io_tensor_rd_0_idx_valid; // @[Load.scala 58:32]
  wire [6:0] tensorLoad_0_io_tensor_rd_0_idx_bits; // @[Load.scala 58:32]
  wire  tensorLoad_0_io_tensor_rd_0_data_valid; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_0_io_tensor_rd_0_data_bits_0_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_0_io_tensor_rd_0_data_bits_0_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_0_io_tensor_rd_0_data_bits_0_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_0_io_tensor_rd_0_data_bits_0_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_0_io_tensor_rd_0_data_bits_0_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_0_io_tensor_rd_0_data_bits_0_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_0_io_tensor_rd_0_data_bits_0_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_0_io_tensor_rd_0_data_bits_0_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_0_io_tensor_rd_0_data_bits_0_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_0_io_tensor_rd_0_data_bits_0_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_0_io_tensor_rd_0_data_bits_0_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_0_io_tensor_rd_0_data_bits_0_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_0_io_tensor_rd_0_data_bits_0_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_0_io_tensor_rd_0_data_bits_0_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_0_io_tensor_rd_0_data_bits_0_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_0_io_tensor_rd_0_data_bits_0_15; // @[Load.scala 58:32]
  wire  tensorLoad_1_clock; // @[Load.scala 58:32]
  wire  tensorLoad_1_reset; // @[Load.scala 58:32]
  wire  tensorLoad_1_io_start; // @[Load.scala 58:32]
  wire  tensorLoad_1_io_done; // @[Load.scala 58:32]
  wire [127:0] tensorLoad_1_io_inst; // @[Load.scala 58:32]
  wire [31:0] tensorLoad_1_io_baddr; // @[Load.scala 58:32]
  wire  tensorLoad_1_io_vme_rd_cmd_ready; // @[Load.scala 58:32]
  wire  tensorLoad_1_io_vme_rd_cmd_valid; // @[Load.scala 58:32]
  wire [31:0] tensorLoad_1_io_vme_rd_cmd_bits_addr; // @[Load.scala 58:32]
  wire [3:0] tensorLoad_1_io_vme_rd_cmd_bits_len; // @[Load.scala 58:32]
  wire [20:0] tensorLoad_1_io_vme_rd_cmd_bits_tag; // @[Load.scala 58:32]
  wire  tensorLoad_1_io_vme_rd_data_valid; // @[Load.scala 58:32]
  wire [63:0] tensorLoad_1_io_vme_rd_data_bits_data; // @[Load.scala 58:32]
  wire [20:0] tensorLoad_1_io_vme_rd_data_bits_tag; // @[Load.scala 58:32]
  wire  tensorLoad_1_io_tensor_rd_0_idx_valid; // @[Load.scala 58:32]
  wire [5:0] tensorLoad_1_io_tensor_rd_0_idx_bits; // @[Load.scala 58:32]
  wire  tensorLoad_1_io_tensor_rd_0_data_valid; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_0_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_0_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_0_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_0_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_0_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_0_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_0_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_0_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_0_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_0_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_0_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_0_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_0_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_0_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_0_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_0_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_1_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_1_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_1_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_1_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_1_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_1_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_1_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_1_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_1_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_1_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_1_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_1_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_1_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_1_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_1_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_1_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_2_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_2_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_2_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_2_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_2_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_2_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_2_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_2_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_2_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_2_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_2_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_2_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_2_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_2_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_2_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_2_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_3_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_3_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_3_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_3_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_3_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_3_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_3_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_3_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_3_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_3_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_3_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_3_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_3_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_3_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_3_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_3_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_4_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_4_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_4_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_4_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_4_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_4_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_4_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_4_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_4_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_4_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_4_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_4_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_4_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_4_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_4_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_4_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_5_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_5_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_5_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_5_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_5_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_5_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_5_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_5_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_5_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_5_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_5_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_5_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_5_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_5_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_5_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_5_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_6_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_6_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_6_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_6_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_6_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_6_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_6_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_6_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_6_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_6_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_6_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_6_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_6_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_6_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_6_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_6_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_7_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_7_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_7_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_7_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_7_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_7_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_7_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_7_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_7_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_7_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_7_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_7_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_7_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_7_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_7_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_7_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_8_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_8_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_8_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_8_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_8_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_8_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_8_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_8_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_8_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_8_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_8_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_8_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_8_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_8_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_8_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_8_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_9_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_9_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_9_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_9_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_9_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_9_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_9_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_9_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_9_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_9_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_9_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_9_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_9_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_9_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_9_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_9_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_10_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_10_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_10_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_10_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_10_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_10_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_10_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_10_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_10_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_10_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_10_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_10_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_10_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_10_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_10_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_10_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_11_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_11_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_11_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_11_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_11_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_11_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_11_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_11_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_11_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_11_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_11_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_11_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_11_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_11_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_11_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_11_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_12_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_12_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_12_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_12_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_12_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_12_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_12_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_12_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_12_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_12_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_12_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_12_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_12_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_12_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_12_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_12_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_13_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_13_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_13_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_13_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_13_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_13_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_13_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_13_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_13_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_13_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_13_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_13_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_13_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_13_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_13_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_13_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_14_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_14_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_14_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_14_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_14_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_14_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_14_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_14_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_14_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_14_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_14_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_14_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_14_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_14_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_14_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_14_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_15_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_15_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_15_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_15_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_15_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_15_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_15_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_15_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_15_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_15_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_15_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_15_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_15_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_15_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_15_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_15_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_16_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_16_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_16_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_16_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_16_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_16_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_16_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_16_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_16_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_16_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_16_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_16_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_16_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_16_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_16_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_16_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_17_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_17_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_17_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_17_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_17_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_17_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_17_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_17_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_17_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_17_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_17_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_17_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_17_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_17_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_17_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_17_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_18_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_18_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_18_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_18_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_18_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_18_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_18_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_18_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_18_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_18_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_18_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_18_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_18_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_18_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_18_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_18_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_19_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_19_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_19_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_19_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_19_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_19_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_19_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_19_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_19_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_19_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_19_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_19_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_19_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_19_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_19_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_19_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_20_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_20_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_20_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_20_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_20_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_20_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_20_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_20_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_20_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_20_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_20_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_20_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_20_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_20_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_20_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_20_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_21_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_21_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_21_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_21_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_21_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_21_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_21_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_21_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_21_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_21_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_21_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_21_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_21_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_21_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_21_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_21_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_22_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_22_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_22_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_22_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_22_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_22_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_22_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_22_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_22_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_22_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_22_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_22_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_22_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_22_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_22_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_22_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_23_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_23_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_23_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_23_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_23_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_23_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_23_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_23_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_23_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_23_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_23_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_23_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_23_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_23_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_23_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_23_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_24_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_24_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_24_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_24_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_24_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_24_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_24_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_24_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_24_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_24_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_24_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_24_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_24_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_24_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_24_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_24_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_25_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_25_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_25_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_25_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_25_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_25_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_25_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_25_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_25_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_25_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_25_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_25_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_25_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_25_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_25_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_25_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_26_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_26_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_26_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_26_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_26_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_26_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_26_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_26_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_26_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_26_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_26_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_26_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_26_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_26_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_26_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_26_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_27_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_27_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_27_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_27_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_27_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_27_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_27_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_27_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_27_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_27_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_27_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_27_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_27_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_27_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_27_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_27_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_28_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_28_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_28_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_28_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_28_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_28_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_28_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_28_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_28_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_28_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_28_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_28_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_28_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_28_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_28_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_28_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_29_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_29_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_29_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_29_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_29_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_29_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_29_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_29_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_29_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_29_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_29_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_29_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_29_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_29_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_29_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_29_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_30_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_30_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_30_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_30_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_30_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_30_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_30_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_30_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_30_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_30_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_30_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_30_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_30_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_30_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_30_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_30_15; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_31_0; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_31_1; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_31_2; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_31_3; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_31_4; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_31_5; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_31_6; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_31_7; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_31_8; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_31_9; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_31_10; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_31_11; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_31_12; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_31_13; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_31_14; // @[Load.scala 58:32]
  wire [7:0] tensorLoad_1_io_tensor_rd_0_data_bits_31_15; // @[Load.scala 58:32]
  reg [1:0] state; // @[Load.scala 47:22]
  wire  _start_T = dec_io_pop_next ? s_io_sready : 1'h1; // @[Load.scala 60:40]
  wire  start = inst_q_io_deq_valid & _start_T; // @[Load.scala 60:35]
  wire  done = dec_io_isInput ? tensorLoad_0_io_done : tensorLoad_1_io_done; // @[Load.scala 61:17]
  wire [1:0] _GEN_0 = dec_io_isInput | dec_io_isWeight ? 2'h2 : state; // @[Load.scala 69:55 70:17 47:22]
  wire [1:0] _GEN_3 = done ? 2'h0 : state; // @[Load.scala 78:18 79:15 47:22]
  wire  _inst_q_io_deq_ready_T_3 = state == 2'h2 & done | state == 2'h1; // @[Load.scala 86:50]
  wire  _tensorLoad_0_io_start_T_1 = state == 2'h0 & start; // @[Load.scala 94:47]
  Semaphore s ( // @[Load.scala 49:17]
    .clock(s_clock),
    .reset(s_reset),
    .io_spost(s_io_spost),
    .io_swait(s_io_swait),
    .io_sready(s_io_sready)
  );
  Queue_6 inst_q ( // @[Load.scala 50:22]
    .clock(inst_q_clock),
    .reset(inst_q_reset),
    .io_enq_ready(inst_q_io_enq_ready),
    .io_enq_valid(inst_q_io_enq_valid),
    .io_enq_bits(inst_q_io_enq_bits),
    .io_deq_ready(inst_q_io_deq_ready),
    .io_deq_valid(inst_q_io_deq_valid),
    .io_deq_bits(inst_q_io_deq_bits)
  );
  LoadDecode dec ( // @[Load.scala 52:19]
    .io_inst(dec_io_inst),
    .io_push_next(dec_io_push_next),
    .io_pop_next(dec_io_pop_next),
    .io_isInput(dec_io_isInput),
    .io_isWeight(dec_io_isWeight),
    .io_isSync(dec_io_isSync)
  );
  TensorLoadInp tensorLoad_0 ( // @[Load.scala 58:32]
    .clock(tensorLoad_0_clock),
    .reset(tensorLoad_0_reset),
    .io_start(tensorLoad_0_io_start),
    .io_done(tensorLoad_0_io_done),
    .io_inst(tensorLoad_0_io_inst),
    .io_baddr(tensorLoad_0_io_baddr),
    .io_vme_rd_cmd_ready(tensorLoad_0_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(tensorLoad_0_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(tensorLoad_0_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(tensorLoad_0_io_vme_rd_cmd_bits_len),
    .io_vme_rd_cmd_bits_tag(tensorLoad_0_io_vme_rd_cmd_bits_tag),
    .io_vme_rd_data_valid(tensorLoad_0_io_vme_rd_data_valid),
    .io_vme_rd_data_bits_data(tensorLoad_0_io_vme_rd_data_bits_data),
    .io_vme_rd_data_bits_tag(tensorLoad_0_io_vme_rd_data_bits_tag),
    .io_tensor_rd_0_idx_valid(tensorLoad_0_io_tensor_rd_0_idx_valid),
    .io_tensor_rd_0_idx_bits(tensorLoad_0_io_tensor_rd_0_idx_bits),
    .io_tensor_rd_0_data_valid(tensorLoad_0_io_tensor_rd_0_data_valid),
    .io_tensor_rd_0_data_bits_0_0(tensorLoad_0_io_tensor_rd_0_data_bits_0_0),
    .io_tensor_rd_0_data_bits_0_1(tensorLoad_0_io_tensor_rd_0_data_bits_0_1),
    .io_tensor_rd_0_data_bits_0_2(tensorLoad_0_io_tensor_rd_0_data_bits_0_2),
    .io_tensor_rd_0_data_bits_0_3(tensorLoad_0_io_tensor_rd_0_data_bits_0_3),
    .io_tensor_rd_0_data_bits_0_4(tensorLoad_0_io_tensor_rd_0_data_bits_0_4),
    .io_tensor_rd_0_data_bits_0_5(tensorLoad_0_io_tensor_rd_0_data_bits_0_5),
    .io_tensor_rd_0_data_bits_0_6(tensorLoad_0_io_tensor_rd_0_data_bits_0_6),
    .io_tensor_rd_0_data_bits_0_7(tensorLoad_0_io_tensor_rd_0_data_bits_0_7),
    .io_tensor_rd_0_data_bits_0_8(tensorLoad_0_io_tensor_rd_0_data_bits_0_8),
    .io_tensor_rd_0_data_bits_0_9(tensorLoad_0_io_tensor_rd_0_data_bits_0_9),
    .io_tensor_rd_0_data_bits_0_10(tensorLoad_0_io_tensor_rd_0_data_bits_0_10),
    .io_tensor_rd_0_data_bits_0_11(tensorLoad_0_io_tensor_rd_0_data_bits_0_11),
    .io_tensor_rd_0_data_bits_0_12(tensorLoad_0_io_tensor_rd_0_data_bits_0_12),
    .io_tensor_rd_0_data_bits_0_13(tensorLoad_0_io_tensor_rd_0_data_bits_0_13),
    .io_tensor_rd_0_data_bits_0_14(tensorLoad_0_io_tensor_rd_0_data_bits_0_14),
    .io_tensor_rd_0_data_bits_0_15(tensorLoad_0_io_tensor_rd_0_data_bits_0_15)
  );
  TensorLoadWgt tensorLoad_1 ( // @[Load.scala 58:32]
    .clock(tensorLoad_1_clock),
    .reset(tensorLoad_1_reset),
    .io_start(tensorLoad_1_io_start),
    .io_done(tensorLoad_1_io_done),
    .io_inst(tensorLoad_1_io_inst),
    .io_baddr(tensorLoad_1_io_baddr),
    .io_vme_rd_cmd_ready(tensorLoad_1_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(tensorLoad_1_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(tensorLoad_1_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(tensorLoad_1_io_vme_rd_cmd_bits_len),
    .io_vme_rd_cmd_bits_tag(tensorLoad_1_io_vme_rd_cmd_bits_tag),
    .io_vme_rd_data_valid(tensorLoad_1_io_vme_rd_data_valid),
    .io_vme_rd_data_bits_data(tensorLoad_1_io_vme_rd_data_bits_data),
    .io_vme_rd_data_bits_tag(tensorLoad_1_io_vme_rd_data_bits_tag),
    .io_tensor_rd_0_idx_valid(tensorLoad_1_io_tensor_rd_0_idx_valid),
    .io_tensor_rd_0_idx_bits(tensorLoad_1_io_tensor_rd_0_idx_bits),
    .io_tensor_rd_0_data_valid(tensorLoad_1_io_tensor_rd_0_data_valid),
    .io_tensor_rd_0_data_bits_0_0(tensorLoad_1_io_tensor_rd_0_data_bits_0_0),
    .io_tensor_rd_0_data_bits_0_1(tensorLoad_1_io_tensor_rd_0_data_bits_0_1),
    .io_tensor_rd_0_data_bits_0_2(tensorLoad_1_io_tensor_rd_0_data_bits_0_2),
    .io_tensor_rd_0_data_bits_0_3(tensorLoad_1_io_tensor_rd_0_data_bits_0_3),
    .io_tensor_rd_0_data_bits_0_4(tensorLoad_1_io_tensor_rd_0_data_bits_0_4),
    .io_tensor_rd_0_data_bits_0_5(tensorLoad_1_io_tensor_rd_0_data_bits_0_5),
    .io_tensor_rd_0_data_bits_0_6(tensorLoad_1_io_tensor_rd_0_data_bits_0_6),
    .io_tensor_rd_0_data_bits_0_7(tensorLoad_1_io_tensor_rd_0_data_bits_0_7),
    .io_tensor_rd_0_data_bits_0_8(tensorLoad_1_io_tensor_rd_0_data_bits_0_8),
    .io_tensor_rd_0_data_bits_0_9(tensorLoad_1_io_tensor_rd_0_data_bits_0_9),
    .io_tensor_rd_0_data_bits_0_10(tensorLoad_1_io_tensor_rd_0_data_bits_0_10),
    .io_tensor_rd_0_data_bits_0_11(tensorLoad_1_io_tensor_rd_0_data_bits_0_11),
    .io_tensor_rd_0_data_bits_0_12(tensorLoad_1_io_tensor_rd_0_data_bits_0_12),
    .io_tensor_rd_0_data_bits_0_13(tensorLoad_1_io_tensor_rd_0_data_bits_0_13),
    .io_tensor_rd_0_data_bits_0_14(tensorLoad_1_io_tensor_rd_0_data_bits_0_14),
    .io_tensor_rd_0_data_bits_0_15(tensorLoad_1_io_tensor_rd_0_data_bits_0_15),
    .io_tensor_rd_0_data_bits_1_0(tensorLoad_1_io_tensor_rd_0_data_bits_1_0),
    .io_tensor_rd_0_data_bits_1_1(tensorLoad_1_io_tensor_rd_0_data_bits_1_1),
    .io_tensor_rd_0_data_bits_1_2(tensorLoad_1_io_tensor_rd_0_data_bits_1_2),
    .io_tensor_rd_0_data_bits_1_3(tensorLoad_1_io_tensor_rd_0_data_bits_1_3),
    .io_tensor_rd_0_data_bits_1_4(tensorLoad_1_io_tensor_rd_0_data_bits_1_4),
    .io_tensor_rd_0_data_bits_1_5(tensorLoad_1_io_tensor_rd_0_data_bits_1_5),
    .io_tensor_rd_0_data_bits_1_6(tensorLoad_1_io_tensor_rd_0_data_bits_1_6),
    .io_tensor_rd_0_data_bits_1_7(tensorLoad_1_io_tensor_rd_0_data_bits_1_7),
    .io_tensor_rd_0_data_bits_1_8(tensorLoad_1_io_tensor_rd_0_data_bits_1_8),
    .io_tensor_rd_0_data_bits_1_9(tensorLoad_1_io_tensor_rd_0_data_bits_1_9),
    .io_tensor_rd_0_data_bits_1_10(tensorLoad_1_io_tensor_rd_0_data_bits_1_10),
    .io_tensor_rd_0_data_bits_1_11(tensorLoad_1_io_tensor_rd_0_data_bits_1_11),
    .io_tensor_rd_0_data_bits_1_12(tensorLoad_1_io_tensor_rd_0_data_bits_1_12),
    .io_tensor_rd_0_data_bits_1_13(tensorLoad_1_io_tensor_rd_0_data_bits_1_13),
    .io_tensor_rd_0_data_bits_1_14(tensorLoad_1_io_tensor_rd_0_data_bits_1_14),
    .io_tensor_rd_0_data_bits_1_15(tensorLoad_1_io_tensor_rd_0_data_bits_1_15),
    .io_tensor_rd_0_data_bits_2_0(tensorLoad_1_io_tensor_rd_0_data_bits_2_0),
    .io_tensor_rd_0_data_bits_2_1(tensorLoad_1_io_tensor_rd_0_data_bits_2_1),
    .io_tensor_rd_0_data_bits_2_2(tensorLoad_1_io_tensor_rd_0_data_bits_2_2),
    .io_tensor_rd_0_data_bits_2_3(tensorLoad_1_io_tensor_rd_0_data_bits_2_3),
    .io_tensor_rd_0_data_bits_2_4(tensorLoad_1_io_tensor_rd_0_data_bits_2_4),
    .io_tensor_rd_0_data_bits_2_5(tensorLoad_1_io_tensor_rd_0_data_bits_2_5),
    .io_tensor_rd_0_data_bits_2_6(tensorLoad_1_io_tensor_rd_0_data_bits_2_6),
    .io_tensor_rd_0_data_bits_2_7(tensorLoad_1_io_tensor_rd_0_data_bits_2_7),
    .io_tensor_rd_0_data_bits_2_8(tensorLoad_1_io_tensor_rd_0_data_bits_2_8),
    .io_tensor_rd_0_data_bits_2_9(tensorLoad_1_io_tensor_rd_0_data_bits_2_9),
    .io_tensor_rd_0_data_bits_2_10(tensorLoad_1_io_tensor_rd_0_data_bits_2_10),
    .io_tensor_rd_0_data_bits_2_11(tensorLoad_1_io_tensor_rd_0_data_bits_2_11),
    .io_tensor_rd_0_data_bits_2_12(tensorLoad_1_io_tensor_rd_0_data_bits_2_12),
    .io_tensor_rd_0_data_bits_2_13(tensorLoad_1_io_tensor_rd_0_data_bits_2_13),
    .io_tensor_rd_0_data_bits_2_14(tensorLoad_1_io_tensor_rd_0_data_bits_2_14),
    .io_tensor_rd_0_data_bits_2_15(tensorLoad_1_io_tensor_rd_0_data_bits_2_15),
    .io_tensor_rd_0_data_bits_3_0(tensorLoad_1_io_tensor_rd_0_data_bits_3_0),
    .io_tensor_rd_0_data_bits_3_1(tensorLoad_1_io_tensor_rd_0_data_bits_3_1),
    .io_tensor_rd_0_data_bits_3_2(tensorLoad_1_io_tensor_rd_0_data_bits_3_2),
    .io_tensor_rd_0_data_bits_3_3(tensorLoad_1_io_tensor_rd_0_data_bits_3_3),
    .io_tensor_rd_0_data_bits_3_4(tensorLoad_1_io_tensor_rd_0_data_bits_3_4),
    .io_tensor_rd_0_data_bits_3_5(tensorLoad_1_io_tensor_rd_0_data_bits_3_5),
    .io_tensor_rd_0_data_bits_3_6(tensorLoad_1_io_tensor_rd_0_data_bits_3_6),
    .io_tensor_rd_0_data_bits_3_7(tensorLoad_1_io_tensor_rd_0_data_bits_3_7),
    .io_tensor_rd_0_data_bits_3_8(tensorLoad_1_io_tensor_rd_0_data_bits_3_8),
    .io_tensor_rd_0_data_bits_3_9(tensorLoad_1_io_tensor_rd_0_data_bits_3_9),
    .io_tensor_rd_0_data_bits_3_10(tensorLoad_1_io_tensor_rd_0_data_bits_3_10),
    .io_tensor_rd_0_data_bits_3_11(tensorLoad_1_io_tensor_rd_0_data_bits_3_11),
    .io_tensor_rd_0_data_bits_3_12(tensorLoad_1_io_tensor_rd_0_data_bits_3_12),
    .io_tensor_rd_0_data_bits_3_13(tensorLoad_1_io_tensor_rd_0_data_bits_3_13),
    .io_tensor_rd_0_data_bits_3_14(tensorLoad_1_io_tensor_rd_0_data_bits_3_14),
    .io_tensor_rd_0_data_bits_3_15(tensorLoad_1_io_tensor_rd_0_data_bits_3_15),
    .io_tensor_rd_0_data_bits_4_0(tensorLoad_1_io_tensor_rd_0_data_bits_4_0),
    .io_tensor_rd_0_data_bits_4_1(tensorLoad_1_io_tensor_rd_0_data_bits_4_1),
    .io_tensor_rd_0_data_bits_4_2(tensorLoad_1_io_tensor_rd_0_data_bits_4_2),
    .io_tensor_rd_0_data_bits_4_3(tensorLoad_1_io_tensor_rd_0_data_bits_4_3),
    .io_tensor_rd_0_data_bits_4_4(tensorLoad_1_io_tensor_rd_0_data_bits_4_4),
    .io_tensor_rd_0_data_bits_4_5(tensorLoad_1_io_tensor_rd_0_data_bits_4_5),
    .io_tensor_rd_0_data_bits_4_6(tensorLoad_1_io_tensor_rd_0_data_bits_4_6),
    .io_tensor_rd_0_data_bits_4_7(tensorLoad_1_io_tensor_rd_0_data_bits_4_7),
    .io_tensor_rd_0_data_bits_4_8(tensorLoad_1_io_tensor_rd_0_data_bits_4_8),
    .io_tensor_rd_0_data_bits_4_9(tensorLoad_1_io_tensor_rd_0_data_bits_4_9),
    .io_tensor_rd_0_data_bits_4_10(tensorLoad_1_io_tensor_rd_0_data_bits_4_10),
    .io_tensor_rd_0_data_bits_4_11(tensorLoad_1_io_tensor_rd_0_data_bits_4_11),
    .io_tensor_rd_0_data_bits_4_12(tensorLoad_1_io_tensor_rd_0_data_bits_4_12),
    .io_tensor_rd_0_data_bits_4_13(tensorLoad_1_io_tensor_rd_0_data_bits_4_13),
    .io_tensor_rd_0_data_bits_4_14(tensorLoad_1_io_tensor_rd_0_data_bits_4_14),
    .io_tensor_rd_0_data_bits_4_15(tensorLoad_1_io_tensor_rd_0_data_bits_4_15),
    .io_tensor_rd_0_data_bits_5_0(tensorLoad_1_io_tensor_rd_0_data_bits_5_0),
    .io_tensor_rd_0_data_bits_5_1(tensorLoad_1_io_tensor_rd_0_data_bits_5_1),
    .io_tensor_rd_0_data_bits_5_2(tensorLoad_1_io_tensor_rd_0_data_bits_5_2),
    .io_tensor_rd_0_data_bits_5_3(tensorLoad_1_io_tensor_rd_0_data_bits_5_3),
    .io_tensor_rd_0_data_bits_5_4(tensorLoad_1_io_tensor_rd_0_data_bits_5_4),
    .io_tensor_rd_0_data_bits_5_5(tensorLoad_1_io_tensor_rd_0_data_bits_5_5),
    .io_tensor_rd_0_data_bits_5_6(tensorLoad_1_io_tensor_rd_0_data_bits_5_6),
    .io_tensor_rd_0_data_bits_5_7(tensorLoad_1_io_tensor_rd_0_data_bits_5_7),
    .io_tensor_rd_0_data_bits_5_8(tensorLoad_1_io_tensor_rd_0_data_bits_5_8),
    .io_tensor_rd_0_data_bits_5_9(tensorLoad_1_io_tensor_rd_0_data_bits_5_9),
    .io_tensor_rd_0_data_bits_5_10(tensorLoad_1_io_tensor_rd_0_data_bits_5_10),
    .io_tensor_rd_0_data_bits_5_11(tensorLoad_1_io_tensor_rd_0_data_bits_5_11),
    .io_tensor_rd_0_data_bits_5_12(tensorLoad_1_io_tensor_rd_0_data_bits_5_12),
    .io_tensor_rd_0_data_bits_5_13(tensorLoad_1_io_tensor_rd_0_data_bits_5_13),
    .io_tensor_rd_0_data_bits_5_14(tensorLoad_1_io_tensor_rd_0_data_bits_5_14),
    .io_tensor_rd_0_data_bits_5_15(tensorLoad_1_io_tensor_rd_0_data_bits_5_15),
    .io_tensor_rd_0_data_bits_6_0(tensorLoad_1_io_tensor_rd_0_data_bits_6_0),
    .io_tensor_rd_0_data_bits_6_1(tensorLoad_1_io_tensor_rd_0_data_bits_6_1),
    .io_tensor_rd_0_data_bits_6_2(tensorLoad_1_io_tensor_rd_0_data_bits_6_2),
    .io_tensor_rd_0_data_bits_6_3(tensorLoad_1_io_tensor_rd_0_data_bits_6_3),
    .io_tensor_rd_0_data_bits_6_4(tensorLoad_1_io_tensor_rd_0_data_bits_6_4),
    .io_tensor_rd_0_data_bits_6_5(tensorLoad_1_io_tensor_rd_0_data_bits_6_5),
    .io_tensor_rd_0_data_bits_6_6(tensorLoad_1_io_tensor_rd_0_data_bits_6_6),
    .io_tensor_rd_0_data_bits_6_7(tensorLoad_1_io_tensor_rd_0_data_bits_6_7),
    .io_tensor_rd_0_data_bits_6_8(tensorLoad_1_io_tensor_rd_0_data_bits_6_8),
    .io_tensor_rd_0_data_bits_6_9(tensorLoad_1_io_tensor_rd_0_data_bits_6_9),
    .io_tensor_rd_0_data_bits_6_10(tensorLoad_1_io_tensor_rd_0_data_bits_6_10),
    .io_tensor_rd_0_data_bits_6_11(tensorLoad_1_io_tensor_rd_0_data_bits_6_11),
    .io_tensor_rd_0_data_bits_6_12(tensorLoad_1_io_tensor_rd_0_data_bits_6_12),
    .io_tensor_rd_0_data_bits_6_13(tensorLoad_1_io_tensor_rd_0_data_bits_6_13),
    .io_tensor_rd_0_data_bits_6_14(tensorLoad_1_io_tensor_rd_0_data_bits_6_14),
    .io_tensor_rd_0_data_bits_6_15(tensorLoad_1_io_tensor_rd_0_data_bits_6_15),
    .io_tensor_rd_0_data_bits_7_0(tensorLoad_1_io_tensor_rd_0_data_bits_7_0),
    .io_tensor_rd_0_data_bits_7_1(tensorLoad_1_io_tensor_rd_0_data_bits_7_1),
    .io_tensor_rd_0_data_bits_7_2(tensorLoad_1_io_tensor_rd_0_data_bits_7_2),
    .io_tensor_rd_0_data_bits_7_3(tensorLoad_1_io_tensor_rd_0_data_bits_7_3),
    .io_tensor_rd_0_data_bits_7_4(tensorLoad_1_io_tensor_rd_0_data_bits_7_4),
    .io_tensor_rd_0_data_bits_7_5(tensorLoad_1_io_tensor_rd_0_data_bits_7_5),
    .io_tensor_rd_0_data_bits_7_6(tensorLoad_1_io_tensor_rd_0_data_bits_7_6),
    .io_tensor_rd_0_data_bits_7_7(tensorLoad_1_io_tensor_rd_0_data_bits_7_7),
    .io_tensor_rd_0_data_bits_7_8(tensorLoad_1_io_tensor_rd_0_data_bits_7_8),
    .io_tensor_rd_0_data_bits_7_9(tensorLoad_1_io_tensor_rd_0_data_bits_7_9),
    .io_tensor_rd_0_data_bits_7_10(tensorLoad_1_io_tensor_rd_0_data_bits_7_10),
    .io_tensor_rd_0_data_bits_7_11(tensorLoad_1_io_tensor_rd_0_data_bits_7_11),
    .io_tensor_rd_0_data_bits_7_12(tensorLoad_1_io_tensor_rd_0_data_bits_7_12),
    .io_tensor_rd_0_data_bits_7_13(tensorLoad_1_io_tensor_rd_0_data_bits_7_13),
    .io_tensor_rd_0_data_bits_7_14(tensorLoad_1_io_tensor_rd_0_data_bits_7_14),
    .io_tensor_rd_0_data_bits_7_15(tensorLoad_1_io_tensor_rd_0_data_bits_7_15),
    .io_tensor_rd_0_data_bits_8_0(tensorLoad_1_io_tensor_rd_0_data_bits_8_0),
    .io_tensor_rd_0_data_bits_8_1(tensorLoad_1_io_tensor_rd_0_data_bits_8_1),
    .io_tensor_rd_0_data_bits_8_2(tensorLoad_1_io_tensor_rd_0_data_bits_8_2),
    .io_tensor_rd_0_data_bits_8_3(tensorLoad_1_io_tensor_rd_0_data_bits_8_3),
    .io_tensor_rd_0_data_bits_8_4(tensorLoad_1_io_tensor_rd_0_data_bits_8_4),
    .io_tensor_rd_0_data_bits_8_5(tensorLoad_1_io_tensor_rd_0_data_bits_8_5),
    .io_tensor_rd_0_data_bits_8_6(tensorLoad_1_io_tensor_rd_0_data_bits_8_6),
    .io_tensor_rd_0_data_bits_8_7(tensorLoad_1_io_tensor_rd_0_data_bits_8_7),
    .io_tensor_rd_0_data_bits_8_8(tensorLoad_1_io_tensor_rd_0_data_bits_8_8),
    .io_tensor_rd_0_data_bits_8_9(tensorLoad_1_io_tensor_rd_0_data_bits_8_9),
    .io_tensor_rd_0_data_bits_8_10(tensorLoad_1_io_tensor_rd_0_data_bits_8_10),
    .io_tensor_rd_0_data_bits_8_11(tensorLoad_1_io_tensor_rd_0_data_bits_8_11),
    .io_tensor_rd_0_data_bits_8_12(tensorLoad_1_io_tensor_rd_0_data_bits_8_12),
    .io_tensor_rd_0_data_bits_8_13(tensorLoad_1_io_tensor_rd_0_data_bits_8_13),
    .io_tensor_rd_0_data_bits_8_14(tensorLoad_1_io_tensor_rd_0_data_bits_8_14),
    .io_tensor_rd_0_data_bits_8_15(tensorLoad_1_io_tensor_rd_0_data_bits_8_15),
    .io_tensor_rd_0_data_bits_9_0(tensorLoad_1_io_tensor_rd_0_data_bits_9_0),
    .io_tensor_rd_0_data_bits_9_1(tensorLoad_1_io_tensor_rd_0_data_bits_9_1),
    .io_tensor_rd_0_data_bits_9_2(tensorLoad_1_io_tensor_rd_0_data_bits_9_2),
    .io_tensor_rd_0_data_bits_9_3(tensorLoad_1_io_tensor_rd_0_data_bits_9_3),
    .io_tensor_rd_0_data_bits_9_4(tensorLoad_1_io_tensor_rd_0_data_bits_9_4),
    .io_tensor_rd_0_data_bits_9_5(tensorLoad_1_io_tensor_rd_0_data_bits_9_5),
    .io_tensor_rd_0_data_bits_9_6(tensorLoad_1_io_tensor_rd_0_data_bits_9_6),
    .io_tensor_rd_0_data_bits_9_7(tensorLoad_1_io_tensor_rd_0_data_bits_9_7),
    .io_tensor_rd_0_data_bits_9_8(tensorLoad_1_io_tensor_rd_0_data_bits_9_8),
    .io_tensor_rd_0_data_bits_9_9(tensorLoad_1_io_tensor_rd_0_data_bits_9_9),
    .io_tensor_rd_0_data_bits_9_10(tensorLoad_1_io_tensor_rd_0_data_bits_9_10),
    .io_tensor_rd_0_data_bits_9_11(tensorLoad_1_io_tensor_rd_0_data_bits_9_11),
    .io_tensor_rd_0_data_bits_9_12(tensorLoad_1_io_tensor_rd_0_data_bits_9_12),
    .io_tensor_rd_0_data_bits_9_13(tensorLoad_1_io_tensor_rd_0_data_bits_9_13),
    .io_tensor_rd_0_data_bits_9_14(tensorLoad_1_io_tensor_rd_0_data_bits_9_14),
    .io_tensor_rd_0_data_bits_9_15(tensorLoad_1_io_tensor_rd_0_data_bits_9_15),
    .io_tensor_rd_0_data_bits_10_0(tensorLoad_1_io_tensor_rd_0_data_bits_10_0),
    .io_tensor_rd_0_data_bits_10_1(tensorLoad_1_io_tensor_rd_0_data_bits_10_1),
    .io_tensor_rd_0_data_bits_10_2(tensorLoad_1_io_tensor_rd_0_data_bits_10_2),
    .io_tensor_rd_0_data_bits_10_3(tensorLoad_1_io_tensor_rd_0_data_bits_10_3),
    .io_tensor_rd_0_data_bits_10_4(tensorLoad_1_io_tensor_rd_0_data_bits_10_4),
    .io_tensor_rd_0_data_bits_10_5(tensorLoad_1_io_tensor_rd_0_data_bits_10_5),
    .io_tensor_rd_0_data_bits_10_6(tensorLoad_1_io_tensor_rd_0_data_bits_10_6),
    .io_tensor_rd_0_data_bits_10_7(tensorLoad_1_io_tensor_rd_0_data_bits_10_7),
    .io_tensor_rd_0_data_bits_10_8(tensorLoad_1_io_tensor_rd_0_data_bits_10_8),
    .io_tensor_rd_0_data_bits_10_9(tensorLoad_1_io_tensor_rd_0_data_bits_10_9),
    .io_tensor_rd_0_data_bits_10_10(tensorLoad_1_io_tensor_rd_0_data_bits_10_10),
    .io_tensor_rd_0_data_bits_10_11(tensorLoad_1_io_tensor_rd_0_data_bits_10_11),
    .io_tensor_rd_0_data_bits_10_12(tensorLoad_1_io_tensor_rd_0_data_bits_10_12),
    .io_tensor_rd_0_data_bits_10_13(tensorLoad_1_io_tensor_rd_0_data_bits_10_13),
    .io_tensor_rd_0_data_bits_10_14(tensorLoad_1_io_tensor_rd_0_data_bits_10_14),
    .io_tensor_rd_0_data_bits_10_15(tensorLoad_1_io_tensor_rd_0_data_bits_10_15),
    .io_tensor_rd_0_data_bits_11_0(tensorLoad_1_io_tensor_rd_0_data_bits_11_0),
    .io_tensor_rd_0_data_bits_11_1(tensorLoad_1_io_tensor_rd_0_data_bits_11_1),
    .io_tensor_rd_0_data_bits_11_2(tensorLoad_1_io_tensor_rd_0_data_bits_11_2),
    .io_tensor_rd_0_data_bits_11_3(tensorLoad_1_io_tensor_rd_0_data_bits_11_3),
    .io_tensor_rd_0_data_bits_11_4(tensorLoad_1_io_tensor_rd_0_data_bits_11_4),
    .io_tensor_rd_0_data_bits_11_5(tensorLoad_1_io_tensor_rd_0_data_bits_11_5),
    .io_tensor_rd_0_data_bits_11_6(tensorLoad_1_io_tensor_rd_0_data_bits_11_6),
    .io_tensor_rd_0_data_bits_11_7(tensorLoad_1_io_tensor_rd_0_data_bits_11_7),
    .io_tensor_rd_0_data_bits_11_8(tensorLoad_1_io_tensor_rd_0_data_bits_11_8),
    .io_tensor_rd_0_data_bits_11_9(tensorLoad_1_io_tensor_rd_0_data_bits_11_9),
    .io_tensor_rd_0_data_bits_11_10(tensorLoad_1_io_tensor_rd_0_data_bits_11_10),
    .io_tensor_rd_0_data_bits_11_11(tensorLoad_1_io_tensor_rd_0_data_bits_11_11),
    .io_tensor_rd_0_data_bits_11_12(tensorLoad_1_io_tensor_rd_0_data_bits_11_12),
    .io_tensor_rd_0_data_bits_11_13(tensorLoad_1_io_tensor_rd_0_data_bits_11_13),
    .io_tensor_rd_0_data_bits_11_14(tensorLoad_1_io_tensor_rd_0_data_bits_11_14),
    .io_tensor_rd_0_data_bits_11_15(tensorLoad_1_io_tensor_rd_0_data_bits_11_15),
    .io_tensor_rd_0_data_bits_12_0(tensorLoad_1_io_tensor_rd_0_data_bits_12_0),
    .io_tensor_rd_0_data_bits_12_1(tensorLoad_1_io_tensor_rd_0_data_bits_12_1),
    .io_tensor_rd_0_data_bits_12_2(tensorLoad_1_io_tensor_rd_0_data_bits_12_2),
    .io_tensor_rd_0_data_bits_12_3(tensorLoad_1_io_tensor_rd_0_data_bits_12_3),
    .io_tensor_rd_0_data_bits_12_4(tensorLoad_1_io_tensor_rd_0_data_bits_12_4),
    .io_tensor_rd_0_data_bits_12_5(tensorLoad_1_io_tensor_rd_0_data_bits_12_5),
    .io_tensor_rd_0_data_bits_12_6(tensorLoad_1_io_tensor_rd_0_data_bits_12_6),
    .io_tensor_rd_0_data_bits_12_7(tensorLoad_1_io_tensor_rd_0_data_bits_12_7),
    .io_tensor_rd_0_data_bits_12_8(tensorLoad_1_io_tensor_rd_0_data_bits_12_8),
    .io_tensor_rd_0_data_bits_12_9(tensorLoad_1_io_tensor_rd_0_data_bits_12_9),
    .io_tensor_rd_0_data_bits_12_10(tensorLoad_1_io_tensor_rd_0_data_bits_12_10),
    .io_tensor_rd_0_data_bits_12_11(tensorLoad_1_io_tensor_rd_0_data_bits_12_11),
    .io_tensor_rd_0_data_bits_12_12(tensorLoad_1_io_tensor_rd_0_data_bits_12_12),
    .io_tensor_rd_0_data_bits_12_13(tensorLoad_1_io_tensor_rd_0_data_bits_12_13),
    .io_tensor_rd_0_data_bits_12_14(tensorLoad_1_io_tensor_rd_0_data_bits_12_14),
    .io_tensor_rd_0_data_bits_12_15(tensorLoad_1_io_tensor_rd_0_data_bits_12_15),
    .io_tensor_rd_0_data_bits_13_0(tensorLoad_1_io_tensor_rd_0_data_bits_13_0),
    .io_tensor_rd_0_data_bits_13_1(tensorLoad_1_io_tensor_rd_0_data_bits_13_1),
    .io_tensor_rd_0_data_bits_13_2(tensorLoad_1_io_tensor_rd_0_data_bits_13_2),
    .io_tensor_rd_0_data_bits_13_3(tensorLoad_1_io_tensor_rd_0_data_bits_13_3),
    .io_tensor_rd_0_data_bits_13_4(tensorLoad_1_io_tensor_rd_0_data_bits_13_4),
    .io_tensor_rd_0_data_bits_13_5(tensorLoad_1_io_tensor_rd_0_data_bits_13_5),
    .io_tensor_rd_0_data_bits_13_6(tensorLoad_1_io_tensor_rd_0_data_bits_13_6),
    .io_tensor_rd_0_data_bits_13_7(tensorLoad_1_io_tensor_rd_0_data_bits_13_7),
    .io_tensor_rd_0_data_bits_13_8(tensorLoad_1_io_tensor_rd_0_data_bits_13_8),
    .io_tensor_rd_0_data_bits_13_9(tensorLoad_1_io_tensor_rd_0_data_bits_13_9),
    .io_tensor_rd_0_data_bits_13_10(tensorLoad_1_io_tensor_rd_0_data_bits_13_10),
    .io_tensor_rd_0_data_bits_13_11(tensorLoad_1_io_tensor_rd_0_data_bits_13_11),
    .io_tensor_rd_0_data_bits_13_12(tensorLoad_1_io_tensor_rd_0_data_bits_13_12),
    .io_tensor_rd_0_data_bits_13_13(tensorLoad_1_io_tensor_rd_0_data_bits_13_13),
    .io_tensor_rd_0_data_bits_13_14(tensorLoad_1_io_tensor_rd_0_data_bits_13_14),
    .io_tensor_rd_0_data_bits_13_15(tensorLoad_1_io_tensor_rd_0_data_bits_13_15),
    .io_tensor_rd_0_data_bits_14_0(tensorLoad_1_io_tensor_rd_0_data_bits_14_0),
    .io_tensor_rd_0_data_bits_14_1(tensorLoad_1_io_tensor_rd_0_data_bits_14_1),
    .io_tensor_rd_0_data_bits_14_2(tensorLoad_1_io_tensor_rd_0_data_bits_14_2),
    .io_tensor_rd_0_data_bits_14_3(tensorLoad_1_io_tensor_rd_0_data_bits_14_3),
    .io_tensor_rd_0_data_bits_14_4(tensorLoad_1_io_tensor_rd_0_data_bits_14_4),
    .io_tensor_rd_0_data_bits_14_5(tensorLoad_1_io_tensor_rd_0_data_bits_14_5),
    .io_tensor_rd_0_data_bits_14_6(tensorLoad_1_io_tensor_rd_0_data_bits_14_6),
    .io_tensor_rd_0_data_bits_14_7(tensorLoad_1_io_tensor_rd_0_data_bits_14_7),
    .io_tensor_rd_0_data_bits_14_8(tensorLoad_1_io_tensor_rd_0_data_bits_14_8),
    .io_tensor_rd_0_data_bits_14_9(tensorLoad_1_io_tensor_rd_0_data_bits_14_9),
    .io_tensor_rd_0_data_bits_14_10(tensorLoad_1_io_tensor_rd_0_data_bits_14_10),
    .io_tensor_rd_0_data_bits_14_11(tensorLoad_1_io_tensor_rd_0_data_bits_14_11),
    .io_tensor_rd_0_data_bits_14_12(tensorLoad_1_io_tensor_rd_0_data_bits_14_12),
    .io_tensor_rd_0_data_bits_14_13(tensorLoad_1_io_tensor_rd_0_data_bits_14_13),
    .io_tensor_rd_0_data_bits_14_14(tensorLoad_1_io_tensor_rd_0_data_bits_14_14),
    .io_tensor_rd_0_data_bits_14_15(tensorLoad_1_io_tensor_rd_0_data_bits_14_15),
    .io_tensor_rd_0_data_bits_15_0(tensorLoad_1_io_tensor_rd_0_data_bits_15_0),
    .io_tensor_rd_0_data_bits_15_1(tensorLoad_1_io_tensor_rd_0_data_bits_15_1),
    .io_tensor_rd_0_data_bits_15_2(tensorLoad_1_io_tensor_rd_0_data_bits_15_2),
    .io_tensor_rd_0_data_bits_15_3(tensorLoad_1_io_tensor_rd_0_data_bits_15_3),
    .io_tensor_rd_0_data_bits_15_4(tensorLoad_1_io_tensor_rd_0_data_bits_15_4),
    .io_tensor_rd_0_data_bits_15_5(tensorLoad_1_io_tensor_rd_0_data_bits_15_5),
    .io_tensor_rd_0_data_bits_15_6(tensorLoad_1_io_tensor_rd_0_data_bits_15_6),
    .io_tensor_rd_0_data_bits_15_7(tensorLoad_1_io_tensor_rd_0_data_bits_15_7),
    .io_tensor_rd_0_data_bits_15_8(tensorLoad_1_io_tensor_rd_0_data_bits_15_8),
    .io_tensor_rd_0_data_bits_15_9(tensorLoad_1_io_tensor_rd_0_data_bits_15_9),
    .io_tensor_rd_0_data_bits_15_10(tensorLoad_1_io_tensor_rd_0_data_bits_15_10),
    .io_tensor_rd_0_data_bits_15_11(tensorLoad_1_io_tensor_rd_0_data_bits_15_11),
    .io_tensor_rd_0_data_bits_15_12(tensorLoad_1_io_tensor_rd_0_data_bits_15_12),
    .io_tensor_rd_0_data_bits_15_13(tensorLoad_1_io_tensor_rd_0_data_bits_15_13),
    .io_tensor_rd_0_data_bits_15_14(tensorLoad_1_io_tensor_rd_0_data_bits_15_14),
    .io_tensor_rd_0_data_bits_15_15(tensorLoad_1_io_tensor_rd_0_data_bits_15_15),
    .io_tensor_rd_0_data_bits_16_0(tensorLoad_1_io_tensor_rd_0_data_bits_16_0),
    .io_tensor_rd_0_data_bits_16_1(tensorLoad_1_io_tensor_rd_0_data_bits_16_1),
    .io_tensor_rd_0_data_bits_16_2(tensorLoad_1_io_tensor_rd_0_data_bits_16_2),
    .io_tensor_rd_0_data_bits_16_3(tensorLoad_1_io_tensor_rd_0_data_bits_16_3),
    .io_tensor_rd_0_data_bits_16_4(tensorLoad_1_io_tensor_rd_0_data_bits_16_4),
    .io_tensor_rd_0_data_bits_16_5(tensorLoad_1_io_tensor_rd_0_data_bits_16_5),
    .io_tensor_rd_0_data_bits_16_6(tensorLoad_1_io_tensor_rd_0_data_bits_16_6),
    .io_tensor_rd_0_data_bits_16_7(tensorLoad_1_io_tensor_rd_0_data_bits_16_7),
    .io_tensor_rd_0_data_bits_16_8(tensorLoad_1_io_tensor_rd_0_data_bits_16_8),
    .io_tensor_rd_0_data_bits_16_9(tensorLoad_1_io_tensor_rd_0_data_bits_16_9),
    .io_tensor_rd_0_data_bits_16_10(tensorLoad_1_io_tensor_rd_0_data_bits_16_10),
    .io_tensor_rd_0_data_bits_16_11(tensorLoad_1_io_tensor_rd_0_data_bits_16_11),
    .io_tensor_rd_0_data_bits_16_12(tensorLoad_1_io_tensor_rd_0_data_bits_16_12),
    .io_tensor_rd_0_data_bits_16_13(tensorLoad_1_io_tensor_rd_0_data_bits_16_13),
    .io_tensor_rd_0_data_bits_16_14(tensorLoad_1_io_tensor_rd_0_data_bits_16_14),
    .io_tensor_rd_0_data_bits_16_15(tensorLoad_1_io_tensor_rd_0_data_bits_16_15),
    .io_tensor_rd_0_data_bits_17_0(tensorLoad_1_io_tensor_rd_0_data_bits_17_0),
    .io_tensor_rd_0_data_bits_17_1(tensorLoad_1_io_tensor_rd_0_data_bits_17_1),
    .io_tensor_rd_0_data_bits_17_2(tensorLoad_1_io_tensor_rd_0_data_bits_17_2),
    .io_tensor_rd_0_data_bits_17_3(tensorLoad_1_io_tensor_rd_0_data_bits_17_3),
    .io_tensor_rd_0_data_bits_17_4(tensorLoad_1_io_tensor_rd_0_data_bits_17_4),
    .io_tensor_rd_0_data_bits_17_5(tensorLoad_1_io_tensor_rd_0_data_bits_17_5),
    .io_tensor_rd_0_data_bits_17_6(tensorLoad_1_io_tensor_rd_0_data_bits_17_6),
    .io_tensor_rd_0_data_bits_17_7(tensorLoad_1_io_tensor_rd_0_data_bits_17_7),
    .io_tensor_rd_0_data_bits_17_8(tensorLoad_1_io_tensor_rd_0_data_bits_17_8),
    .io_tensor_rd_0_data_bits_17_9(tensorLoad_1_io_tensor_rd_0_data_bits_17_9),
    .io_tensor_rd_0_data_bits_17_10(tensorLoad_1_io_tensor_rd_0_data_bits_17_10),
    .io_tensor_rd_0_data_bits_17_11(tensorLoad_1_io_tensor_rd_0_data_bits_17_11),
    .io_tensor_rd_0_data_bits_17_12(tensorLoad_1_io_tensor_rd_0_data_bits_17_12),
    .io_tensor_rd_0_data_bits_17_13(tensorLoad_1_io_tensor_rd_0_data_bits_17_13),
    .io_tensor_rd_0_data_bits_17_14(tensorLoad_1_io_tensor_rd_0_data_bits_17_14),
    .io_tensor_rd_0_data_bits_17_15(tensorLoad_1_io_tensor_rd_0_data_bits_17_15),
    .io_tensor_rd_0_data_bits_18_0(tensorLoad_1_io_tensor_rd_0_data_bits_18_0),
    .io_tensor_rd_0_data_bits_18_1(tensorLoad_1_io_tensor_rd_0_data_bits_18_1),
    .io_tensor_rd_0_data_bits_18_2(tensorLoad_1_io_tensor_rd_0_data_bits_18_2),
    .io_tensor_rd_0_data_bits_18_3(tensorLoad_1_io_tensor_rd_0_data_bits_18_3),
    .io_tensor_rd_0_data_bits_18_4(tensorLoad_1_io_tensor_rd_0_data_bits_18_4),
    .io_tensor_rd_0_data_bits_18_5(tensorLoad_1_io_tensor_rd_0_data_bits_18_5),
    .io_tensor_rd_0_data_bits_18_6(tensorLoad_1_io_tensor_rd_0_data_bits_18_6),
    .io_tensor_rd_0_data_bits_18_7(tensorLoad_1_io_tensor_rd_0_data_bits_18_7),
    .io_tensor_rd_0_data_bits_18_8(tensorLoad_1_io_tensor_rd_0_data_bits_18_8),
    .io_tensor_rd_0_data_bits_18_9(tensorLoad_1_io_tensor_rd_0_data_bits_18_9),
    .io_tensor_rd_0_data_bits_18_10(tensorLoad_1_io_tensor_rd_0_data_bits_18_10),
    .io_tensor_rd_0_data_bits_18_11(tensorLoad_1_io_tensor_rd_0_data_bits_18_11),
    .io_tensor_rd_0_data_bits_18_12(tensorLoad_1_io_tensor_rd_0_data_bits_18_12),
    .io_tensor_rd_0_data_bits_18_13(tensorLoad_1_io_tensor_rd_0_data_bits_18_13),
    .io_tensor_rd_0_data_bits_18_14(tensorLoad_1_io_tensor_rd_0_data_bits_18_14),
    .io_tensor_rd_0_data_bits_18_15(tensorLoad_1_io_tensor_rd_0_data_bits_18_15),
    .io_tensor_rd_0_data_bits_19_0(tensorLoad_1_io_tensor_rd_0_data_bits_19_0),
    .io_tensor_rd_0_data_bits_19_1(tensorLoad_1_io_tensor_rd_0_data_bits_19_1),
    .io_tensor_rd_0_data_bits_19_2(tensorLoad_1_io_tensor_rd_0_data_bits_19_2),
    .io_tensor_rd_0_data_bits_19_3(tensorLoad_1_io_tensor_rd_0_data_bits_19_3),
    .io_tensor_rd_0_data_bits_19_4(tensorLoad_1_io_tensor_rd_0_data_bits_19_4),
    .io_tensor_rd_0_data_bits_19_5(tensorLoad_1_io_tensor_rd_0_data_bits_19_5),
    .io_tensor_rd_0_data_bits_19_6(tensorLoad_1_io_tensor_rd_0_data_bits_19_6),
    .io_tensor_rd_0_data_bits_19_7(tensorLoad_1_io_tensor_rd_0_data_bits_19_7),
    .io_tensor_rd_0_data_bits_19_8(tensorLoad_1_io_tensor_rd_0_data_bits_19_8),
    .io_tensor_rd_0_data_bits_19_9(tensorLoad_1_io_tensor_rd_0_data_bits_19_9),
    .io_tensor_rd_0_data_bits_19_10(tensorLoad_1_io_tensor_rd_0_data_bits_19_10),
    .io_tensor_rd_0_data_bits_19_11(tensorLoad_1_io_tensor_rd_0_data_bits_19_11),
    .io_tensor_rd_0_data_bits_19_12(tensorLoad_1_io_tensor_rd_0_data_bits_19_12),
    .io_tensor_rd_0_data_bits_19_13(tensorLoad_1_io_tensor_rd_0_data_bits_19_13),
    .io_tensor_rd_0_data_bits_19_14(tensorLoad_1_io_tensor_rd_0_data_bits_19_14),
    .io_tensor_rd_0_data_bits_19_15(tensorLoad_1_io_tensor_rd_0_data_bits_19_15),
    .io_tensor_rd_0_data_bits_20_0(tensorLoad_1_io_tensor_rd_0_data_bits_20_0),
    .io_tensor_rd_0_data_bits_20_1(tensorLoad_1_io_tensor_rd_0_data_bits_20_1),
    .io_tensor_rd_0_data_bits_20_2(tensorLoad_1_io_tensor_rd_0_data_bits_20_2),
    .io_tensor_rd_0_data_bits_20_3(tensorLoad_1_io_tensor_rd_0_data_bits_20_3),
    .io_tensor_rd_0_data_bits_20_4(tensorLoad_1_io_tensor_rd_0_data_bits_20_4),
    .io_tensor_rd_0_data_bits_20_5(tensorLoad_1_io_tensor_rd_0_data_bits_20_5),
    .io_tensor_rd_0_data_bits_20_6(tensorLoad_1_io_tensor_rd_0_data_bits_20_6),
    .io_tensor_rd_0_data_bits_20_7(tensorLoad_1_io_tensor_rd_0_data_bits_20_7),
    .io_tensor_rd_0_data_bits_20_8(tensorLoad_1_io_tensor_rd_0_data_bits_20_8),
    .io_tensor_rd_0_data_bits_20_9(tensorLoad_1_io_tensor_rd_0_data_bits_20_9),
    .io_tensor_rd_0_data_bits_20_10(tensorLoad_1_io_tensor_rd_0_data_bits_20_10),
    .io_tensor_rd_0_data_bits_20_11(tensorLoad_1_io_tensor_rd_0_data_bits_20_11),
    .io_tensor_rd_0_data_bits_20_12(tensorLoad_1_io_tensor_rd_0_data_bits_20_12),
    .io_tensor_rd_0_data_bits_20_13(tensorLoad_1_io_tensor_rd_0_data_bits_20_13),
    .io_tensor_rd_0_data_bits_20_14(tensorLoad_1_io_tensor_rd_0_data_bits_20_14),
    .io_tensor_rd_0_data_bits_20_15(tensorLoad_1_io_tensor_rd_0_data_bits_20_15),
    .io_tensor_rd_0_data_bits_21_0(tensorLoad_1_io_tensor_rd_0_data_bits_21_0),
    .io_tensor_rd_0_data_bits_21_1(tensorLoad_1_io_tensor_rd_0_data_bits_21_1),
    .io_tensor_rd_0_data_bits_21_2(tensorLoad_1_io_tensor_rd_0_data_bits_21_2),
    .io_tensor_rd_0_data_bits_21_3(tensorLoad_1_io_tensor_rd_0_data_bits_21_3),
    .io_tensor_rd_0_data_bits_21_4(tensorLoad_1_io_tensor_rd_0_data_bits_21_4),
    .io_tensor_rd_0_data_bits_21_5(tensorLoad_1_io_tensor_rd_0_data_bits_21_5),
    .io_tensor_rd_0_data_bits_21_6(tensorLoad_1_io_tensor_rd_0_data_bits_21_6),
    .io_tensor_rd_0_data_bits_21_7(tensorLoad_1_io_tensor_rd_0_data_bits_21_7),
    .io_tensor_rd_0_data_bits_21_8(tensorLoad_1_io_tensor_rd_0_data_bits_21_8),
    .io_tensor_rd_0_data_bits_21_9(tensorLoad_1_io_tensor_rd_0_data_bits_21_9),
    .io_tensor_rd_0_data_bits_21_10(tensorLoad_1_io_tensor_rd_0_data_bits_21_10),
    .io_tensor_rd_0_data_bits_21_11(tensorLoad_1_io_tensor_rd_0_data_bits_21_11),
    .io_tensor_rd_0_data_bits_21_12(tensorLoad_1_io_tensor_rd_0_data_bits_21_12),
    .io_tensor_rd_0_data_bits_21_13(tensorLoad_1_io_tensor_rd_0_data_bits_21_13),
    .io_tensor_rd_0_data_bits_21_14(tensorLoad_1_io_tensor_rd_0_data_bits_21_14),
    .io_tensor_rd_0_data_bits_21_15(tensorLoad_1_io_tensor_rd_0_data_bits_21_15),
    .io_tensor_rd_0_data_bits_22_0(tensorLoad_1_io_tensor_rd_0_data_bits_22_0),
    .io_tensor_rd_0_data_bits_22_1(tensorLoad_1_io_tensor_rd_0_data_bits_22_1),
    .io_tensor_rd_0_data_bits_22_2(tensorLoad_1_io_tensor_rd_0_data_bits_22_2),
    .io_tensor_rd_0_data_bits_22_3(tensorLoad_1_io_tensor_rd_0_data_bits_22_3),
    .io_tensor_rd_0_data_bits_22_4(tensorLoad_1_io_tensor_rd_0_data_bits_22_4),
    .io_tensor_rd_0_data_bits_22_5(tensorLoad_1_io_tensor_rd_0_data_bits_22_5),
    .io_tensor_rd_0_data_bits_22_6(tensorLoad_1_io_tensor_rd_0_data_bits_22_6),
    .io_tensor_rd_0_data_bits_22_7(tensorLoad_1_io_tensor_rd_0_data_bits_22_7),
    .io_tensor_rd_0_data_bits_22_8(tensorLoad_1_io_tensor_rd_0_data_bits_22_8),
    .io_tensor_rd_0_data_bits_22_9(tensorLoad_1_io_tensor_rd_0_data_bits_22_9),
    .io_tensor_rd_0_data_bits_22_10(tensorLoad_1_io_tensor_rd_0_data_bits_22_10),
    .io_tensor_rd_0_data_bits_22_11(tensorLoad_1_io_tensor_rd_0_data_bits_22_11),
    .io_tensor_rd_0_data_bits_22_12(tensorLoad_1_io_tensor_rd_0_data_bits_22_12),
    .io_tensor_rd_0_data_bits_22_13(tensorLoad_1_io_tensor_rd_0_data_bits_22_13),
    .io_tensor_rd_0_data_bits_22_14(tensorLoad_1_io_tensor_rd_0_data_bits_22_14),
    .io_tensor_rd_0_data_bits_22_15(tensorLoad_1_io_tensor_rd_0_data_bits_22_15),
    .io_tensor_rd_0_data_bits_23_0(tensorLoad_1_io_tensor_rd_0_data_bits_23_0),
    .io_tensor_rd_0_data_bits_23_1(tensorLoad_1_io_tensor_rd_0_data_bits_23_1),
    .io_tensor_rd_0_data_bits_23_2(tensorLoad_1_io_tensor_rd_0_data_bits_23_2),
    .io_tensor_rd_0_data_bits_23_3(tensorLoad_1_io_tensor_rd_0_data_bits_23_3),
    .io_tensor_rd_0_data_bits_23_4(tensorLoad_1_io_tensor_rd_0_data_bits_23_4),
    .io_tensor_rd_0_data_bits_23_5(tensorLoad_1_io_tensor_rd_0_data_bits_23_5),
    .io_tensor_rd_0_data_bits_23_6(tensorLoad_1_io_tensor_rd_0_data_bits_23_6),
    .io_tensor_rd_0_data_bits_23_7(tensorLoad_1_io_tensor_rd_0_data_bits_23_7),
    .io_tensor_rd_0_data_bits_23_8(tensorLoad_1_io_tensor_rd_0_data_bits_23_8),
    .io_tensor_rd_0_data_bits_23_9(tensorLoad_1_io_tensor_rd_0_data_bits_23_9),
    .io_tensor_rd_0_data_bits_23_10(tensorLoad_1_io_tensor_rd_0_data_bits_23_10),
    .io_tensor_rd_0_data_bits_23_11(tensorLoad_1_io_tensor_rd_0_data_bits_23_11),
    .io_tensor_rd_0_data_bits_23_12(tensorLoad_1_io_tensor_rd_0_data_bits_23_12),
    .io_tensor_rd_0_data_bits_23_13(tensorLoad_1_io_tensor_rd_0_data_bits_23_13),
    .io_tensor_rd_0_data_bits_23_14(tensorLoad_1_io_tensor_rd_0_data_bits_23_14),
    .io_tensor_rd_0_data_bits_23_15(tensorLoad_1_io_tensor_rd_0_data_bits_23_15),
    .io_tensor_rd_0_data_bits_24_0(tensorLoad_1_io_tensor_rd_0_data_bits_24_0),
    .io_tensor_rd_0_data_bits_24_1(tensorLoad_1_io_tensor_rd_0_data_bits_24_1),
    .io_tensor_rd_0_data_bits_24_2(tensorLoad_1_io_tensor_rd_0_data_bits_24_2),
    .io_tensor_rd_0_data_bits_24_3(tensorLoad_1_io_tensor_rd_0_data_bits_24_3),
    .io_tensor_rd_0_data_bits_24_4(tensorLoad_1_io_tensor_rd_0_data_bits_24_4),
    .io_tensor_rd_0_data_bits_24_5(tensorLoad_1_io_tensor_rd_0_data_bits_24_5),
    .io_tensor_rd_0_data_bits_24_6(tensorLoad_1_io_tensor_rd_0_data_bits_24_6),
    .io_tensor_rd_0_data_bits_24_7(tensorLoad_1_io_tensor_rd_0_data_bits_24_7),
    .io_tensor_rd_0_data_bits_24_8(tensorLoad_1_io_tensor_rd_0_data_bits_24_8),
    .io_tensor_rd_0_data_bits_24_9(tensorLoad_1_io_tensor_rd_0_data_bits_24_9),
    .io_tensor_rd_0_data_bits_24_10(tensorLoad_1_io_tensor_rd_0_data_bits_24_10),
    .io_tensor_rd_0_data_bits_24_11(tensorLoad_1_io_tensor_rd_0_data_bits_24_11),
    .io_tensor_rd_0_data_bits_24_12(tensorLoad_1_io_tensor_rd_0_data_bits_24_12),
    .io_tensor_rd_0_data_bits_24_13(tensorLoad_1_io_tensor_rd_0_data_bits_24_13),
    .io_tensor_rd_0_data_bits_24_14(tensorLoad_1_io_tensor_rd_0_data_bits_24_14),
    .io_tensor_rd_0_data_bits_24_15(tensorLoad_1_io_tensor_rd_0_data_bits_24_15),
    .io_tensor_rd_0_data_bits_25_0(tensorLoad_1_io_tensor_rd_0_data_bits_25_0),
    .io_tensor_rd_0_data_bits_25_1(tensorLoad_1_io_tensor_rd_0_data_bits_25_1),
    .io_tensor_rd_0_data_bits_25_2(tensorLoad_1_io_tensor_rd_0_data_bits_25_2),
    .io_tensor_rd_0_data_bits_25_3(tensorLoad_1_io_tensor_rd_0_data_bits_25_3),
    .io_tensor_rd_0_data_bits_25_4(tensorLoad_1_io_tensor_rd_0_data_bits_25_4),
    .io_tensor_rd_0_data_bits_25_5(tensorLoad_1_io_tensor_rd_0_data_bits_25_5),
    .io_tensor_rd_0_data_bits_25_6(tensorLoad_1_io_tensor_rd_0_data_bits_25_6),
    .io_tensor_rd_0_data_bits_25_7(tensorLoad_1_io_tensor_rd_0_data_bits_25_7),
    .io_tensor_rd_0_data_bits_25_8(tensorLoad_1_io_tensor_rd_0_data_bits_25_8),
    .io_tensor_rd_0_data_bits_25_9(tensorLoad_1_io_tensor_rd_0_data_bits_25_9),
    .io_tensor_rd_0_data_bits_25_10(tensorLoad_1_io_tensor_rd_0_data_bits_25_10),
    .io_tensor_rd_0_data_bits_25_11(tensorLoad_1_io_tensor_rd_0_data_bits_25_11),
    .io_tensor_rd_0_data_bits_25_12(tensorLoad_1_io_tensor_rd_0_data_bits_25_12),
    .io_tensor_rd_0_data_bits_25_13(tensorLoad_1_io_tensor_rd_0_data_bits_25_13),
    .io_tensor_rd_0_data_bits_25_14(tensorLoad_1_io_tensor_rd_0_data_bits_25_14),
    .io_tensor_rd_0_data_bits_25_15(tensorLoad_1_io_tensor_rd_0_data_bits_25_15),
    .io_tensor_rd_0_data_bits_26_0(tensorLoad_1_io_tensor_rd_0_data_bits_26_0),
    .io_tensor_rd_0_data_bits_26_1(tensorLoad_1_io_tensor_rd_0_data_bits_26_1),
    .io_tensor_rd_0_data_bits_26_2(tensorLoad_1_io_tensor_rd_0_data_bits_26_2),
    .io_tensor_rd_0_data_bits_26_3(tensorLoad_1_io_tensor_rd_0_data_bits_26_3),
    .io_tensor_rd_0_data_bits_26_4(tensorLoad_1_io_tensor_rd_0_data_bits_26_4),
    .io_tensor_rd_0_data_bits_26_5(tensorLoad_1_io_tensor_rd_0_data_bits_26_5),
    .io_tensor_rd_0_data_bits_26_6(tensorLoad_1_io_tensor_rd_0_data_bits_26_6),
    .io_tensor_rd_0_data_bits_26_7(tensorLoad_1_io_tensor_rd_0_data_bits_26_7),
    .io_tensor_rd_0_data_bits_26_8(tensorLoad_1_io_tensor_rd_0_data_bits_26_8),
    .io_tensor_rd_0_data_bits_26_9(tensorLoad_1_io_tensor_rd_0_data_bits_26_9),
    .io_tensor_rd_0_data_bits_26_10(tensorLoad_1_io_tensor_rd_0_data_bits_26_10),
    .io_tensor_rd_0_data_bits_26_11(tensorLoad_1_io_tensor_rd_0_data_bits_26_11),
    .io_tensor_rd_0_data_bits_26_12(tensorLoad_1_io_tensor_rd_0_data_bits_26_12),
    .io_tensor_rd_0_data_bits_26_13(tensorLoad_1_io_tensor_rd_0_data_bits_26_13),
    .io_tensor_rd_0_data_bits_26_14(tensorLoad_1_io_tensor_rd_0_data_bits_26_14),
    .io_tensor_rd_0_data_bits_26_15(tensorLoad_1_io_tensor_rd_0_data_bits_26_15),
    .io_tensor_rd_0_data_bits_27_0(tensorLoad_1_io_tensor_rd_0_data_bits_27_0),
    .io_tensor_rd_0_data_bits_27_1(tensorLoad_1_io_tensor_rd_0_data_bits_27_1),
    .io_tensor_rd_0_data_bits_27_2(tensorLoad_1_io_tensor_rd_0_data_bits_27_2),
    .io_tensor_rd_0_data_bits_27_3(tensorLoad_1_io_tensor_rd_0_data_bits_27_3),
    .io_tensor_rd_0_data_bits_27_4(tensorLoad_1_io_tensor_rd_0_data_bits_27_4),
    .io_tensor_rd_0_data_bits_27_5(tensorLoad_1_io_tensor_rd_0_data_bits_27_5),
    .io_tensor_rd_0_data_bits_27_6(tensorLoad_1_io_tensor_rd_0_data_bits_27_6),
    .io_tensor_rd_0_data_bits_27_7(tensorLoad_1_io_tensor_rd_0_data_bits_27_7),
    .io_tensor_rd_0_data_bits_27_8(tensorLoad_1_io_tensor_rd_0_data_bits_27_8),
    .io_tensor_rd_0_data_bits_27_9(tensorLoad_1_io_tensor_rd_0_data_bits_27_9),
    .io_tensor_rd_0_data_bits_27_10(tensorLoad_1_io_tensor_rd_0_data_bits_27_10),
    .io_tensor_rd_0_data_bits_27_11(tensorLoad_1_io_tensor_rd_0_data_bits_27_11),
    .io_tensor_rd_0_data_bits_27_12(tensorLoad_1_io_tensor_rd_0_data_bits_27_12),
    .io_tensor_rd_0_data_bits_27_13(tensorLoad_1_io_tensor_rd_0_data_bits_27_13),
    .io_tensor_rd_0_data_bits_27_14(tensorLoad_1_io_tensor_rd_0_data_bits_27_14),
    .io_tensor_rd_0_data_bits_27_15(tensorLoad_1_io_tensor_rd_0_data_bits_27_15),
    .io_tensor_rd_0_data_bits_28_0(tensorLoad_1_io_tensor_rd_0_data_bits_28_0),
    .io_tensor_rd_0_data_bits_28_1(tensorLoad_1_io_tensor_rd_0_data_bits_28_1),
    .io_tensor_rd_0_data_bits_28_2(tensorLoad_1_io_tensor_rd_0_data_bits_28_2),
    .io_tensor_rd_0_data_bits_28_3(tensorLoad_1_io_tensor_rd_0_data_bits_28_3),
    .io_tensor_rd_0_data_bits_28_4(tensorLoad_1_io_tensor_rd_0_data_bits_28_4),
    .io_tensor_rd_0_data_bits_28_5(tensorLoad_1_io_tensor_rd_0_data_bits_28_5),
    .io_tensor_rd_0_data_bits_28_6(tensorLoad_1_io_tensor_rd_0_data_bits_28_6),
    .io_tensor_rd_0_data_bits_28_7(tensorLoad_1_io_tensor_rd_0_data_bits_28_7),
    .io_tensor_rd_0_data_bits_28_8(tensorLoad_1_io_tensor_rd_0_data_bits_28_8),
    .io_tensor_rd_0_data_bits_28_9(tensorLoad_1_io_tensor_rd_0_data_bits_28_9),
    .io_tensor_rd_0_data_bits_28_10(tensorLoad_1_io_tensor_rd_0_data_bits_28_10),
    .io_tensor_rd_0_data_bits_28_11(tensorLoad_1_io_tensor_rd_0_data_bits_28_11),
    .io_tensor_rd_0_data_bits_28_12(tensorLoad_1_io_tensor_rd_0_data_bits_28_12),
    .io_tensor_rd_0_data_bits_28_13(tensorLoad_1_io_tensor_rd_0_data_bits_28_13),
    .io_tensor_rd_0_data_bits_28_14(tensorLoad_1_io_tensor_rd_0_data_bits_28_14),
    .io_tensor_rd_0_data_bits_28_15(tensorLoad_1_io_tensor_rd_0_data_bits_28_15),
    .io_tensor_rd_0_data_bits_29_0(tensorLoad_1_io_tensor_rd_0_data_bits_29_0),
    .io_tensor_rd_0_data_bits_29_1(tensorLoad_1_io_tensor_rd_0_data_bits_29_1),
    .io_tensor_rd_0_data_bits_29_2(tensorLoad_1_io_tensor_rd_0_data_bits_29_2),
    .io_tensor_rd_0_data_bits_29_3(tensorLoad_1_io_tensor_rd_0_data_bits_29_3),
    .io_tensor_rd_0_data_bits_29_4(tensorLoad_1_io_tensor_rd_0_data_bits_29_4),
    .io_tensor_rd_0_data_bits_29_5(tensorLoad_1_io_tensor_rd_0_data_bits_29_5),
    .io_tensor_rd_0_data_bits_29_6(tensorLoad_1_io_tensor_rd_0_data_bits_29_6),
    .io_tensor_rd_0_data_bits_29_7(tensorLoad_1_io_tensor_rd_0_data_bits_29_7),
    .io_tensor_rd_0_data_bits_29_8(tensorLoad_1_io_tensor_rd_0_data_bits_29_8),
    .io_tensor_rd_0_data_bits_29_9(tensorLoad_1_io_tensor_rd_0_data_bits_29_9),
    .io_tensor_rd_0_data_bits_29_10(tensorLoad_1_io_tensor_rd_0_data_bits_29_10),
    .io_tensor_rd_0_data_bits_29_11(tensorLoad_1_io_tensor_rd_0_data_bits_29_11),
    .io_tensor_rd_0_data_bits_29_12(tensorLoad_1_io_tensor_rd_0_data_bits_29_12),
    .io_tensor_rd_0_data_bits_29_13(tensorLoad_1_io_tensor_rd_0_data_bits_29_13),
    .io_tensor_rd_0_data_bits_29_14(tensorLoad_1_io_tensor_rd_0_data_bits_29_14),
    .io_tensor_rd_0_data_bits_29_15(tensorLoad_1_io_tensor_rd_0_data_bits_29_15),
    .io_tensor_rd_0_data_bits_30_0(tensorLoad_1_io_tensor_rd_0_data_bits_30_0),
    .io_tensor_rd_0_data_bits_30_1(tensorLoad_1_io_tensor_rd_0_data_bits_30_1),
    .io_tensor_rd_0_data_bits_30_2(tensorLoad_1_io_tensor_rd_0_data_bits_30_2),
    .io_tensor_rd_0_data_bits_30_3(tensorLoad_1_io_tensor_rd_0_data_bits_30_3),
    .io_tensor_rd_0_data_bits_30_4(tensorLoad_1_io_tensor_rd_0_data_bits_30_4),
    .io_tensor_rd_0_data_bits_30_5(tensorLoad_1_io_tensor_rd_0_data_bits_30_5),
    .io_tensor_rd_0_data_bits_30_6(tensorLoad_1_io_tensor_rd_0_data_bits_30_6),
    .io_tensor_rd_0_data_bits_30_7(tensorLoad_1_io_tensor_rd_0_data_bits_30_7),
    .io_tensor_rd_0_data_bits_30_8(tensorLoad_1_io_tensor_rd_0_data_bits_30_8),
    .io_tensor_rd_0_data_bits_30_9(tensorLoad_1_io_tensor_rd_0_data_bits_30_9),
    .io_tensor_rd_0_data_bits_30_10(tensorLoad_1_io_tensor_rd_0_data_bits_30_10),
    .io_tensor_rd_0_data_bits_30_11(tensorLoad_1_io_tensor_rd_0_data_bits_30_11),
    .io_tensor_rd_0_data_bits_30_12(tensorLoad_1_io_tensor_rd_0_data_bits_30_12),
    .io_tensor_rd_0_data_bits_30_13(tensorLoad_1_io_tensor_rd_0_data_bits_30_13),
    .io_tensor_rd_0_data_bits_30_14(tensorLoad_1_io_tensor_rd_0_data_bits_30_14),
    .io_tensor_rd_0_data_bits_30_15(tensorLoad_1_io_tensor_rd_0_data_bits_30_15),
    .io_tensor_rd_0_data_bits_31_0(tensorLoad_1_io_tensor_rd_0_data_bits_31_0),
    .io_tensor_rd_0_data_bits_31_1(tensorLoad_1_io_tensor_rd_0_data_bits_31_1),
    .io_tensor_rd_0_data_bits_31_2(tensorLoad_1_io_tensor_rd_0_data_bits_31_2),
    .io_tensor_rd_0_data_bits_31_3(tensorLoad_1_io_tensor_rd_0_data_bits_31_3),
    .io_tensor_rd_0_data_bits_31_4(tensorLoad_1_io_tensor_rd_0_data_bits_31_4),
    .io_tensor_rd_0_data_bits_31_5(tensorLoad_1_io_tensor_rd_0_data_bits_31_5),
    .io_tensor_rd_0_data_bits_31_6(tensorLoad_1_io_tensor_rd_0_data_bits_31_6),
    .io_tensor_rd_0_data_bits_31_7(tensorLoad_1_io_tensor_rd_0_data_bits_31_7),
    .io_tensor_rd_0_data_bits_31_8(tensorLoad_1_io_tensor_rd_0_data_bits_31_8),
    .io_tensor_rd_0_data_bits_31_9(tensorLoad_1_io_tensor_rd_0_data_bits_31_9),
    .io_tensor_rd_0_data_bits_31_10(tensorLoad_1_io_tensor_rd_0_data_bits_31_10),
    .io_tensor_rd_0_data_bits_31_11(tensorLoad_1_io_tensor_rd_0_data_bits_31_11),
    .io_tensor_rd_0_data_bits_31_12(tensorLoad_1_io_tensor_rd_0_data_bits_31_12),
    .io_tensor_rd_0_data_bits_31_13(tensorLoad_1_io_tensor_rd_0_data_bits_31_13),
    .io_tensor_rd_0_data_bits_31_14(tensorLoad_1_io_tensor_rd_0_data_bits_31_14),
    .io_tensor_rd_0_data_bits_31_15(tensorLoad_1_io_tensor_rd_0_data_bits_31_15)
  );
  assign io_o_post = dec_io_push_next & _inst_q_io_deq_ready_T_3; // @[Load.scala 104:33]
  assign io_inst_ready = inst_q_io_enq_ready; // @[Load.scala 85:17]
  assign io_vme_rd_0_cmd_valid = tensorLoad_0_io_vme_rd_cmd_valid; // @[Load.scala 98:18]
  assign io_vme_rd_0_cmd_bits_addr = tensorLoad_0_io_vme_rd_cmd_bits_addr; // @[Load.scala 98:18]
  assign io_vme_rd_0_cmd_bits_len = tensorLoad_0_io_vme_rd_cmd_bits_len; // @[Load.scala 98:18]
  assign io_vme_rd_0_cmd_bits_tag = tensorLoad_0_io_vme_rd_cmd_bits_tag; // @[Load.scala 98:18]
  assign io_vme_rd_1_cmd_valid = tensorLoad_1_io_vme_rd_cmd_valid; // @[Load.scala 98:18]
  assign io_vme_rd_1_cmd_bits_addr = tensorLoad_1_io_vme_rd_cmd_bits_addr; // @[Load.scala 98:18]
  assign io_vme_rd_1_cmd_bits_len = tensorLoad_1_io_vme_rd_cmd_bits_len; // @[Load.scala 98:18]
  assign io_vme_rd_1_cmd_bits_tag = tensorLoad_1_io_vme_rd_cmd_bits_tag; // @[Load.scala 98:18]
  assign io_inp_rd_0_data_valid = tensorLoad_0_io_tensor_rd_0_data_valid; // @[Load.scala 97:29]
  assign io_inp_rd_0_data_bits_0_0 = tensorLoad_0_io_tensor_rd_0_data_bits_0_0; // @[Load.scala 97:29]
  assign io_inp_rd_0_data_bits_0_1 = tensorLoad_0_io_tensor_rd_0_data_bits_0_1; // @[Load.scala 97:29]
  assign io_inp_rd_0_data_bits_0_2 = tensorLoad_0_io_tensor_rd_0_data_bits_0_2; // @[Load.scala 97:29]
  assign io_inp_rd_0_data_bits_0_3 = tensorLoad_0_io_tensor_rd_0_data_bits_0_3; // @[Load.scala 97:29]
  assign io_inp_rd_0_data_bits_0_4 = tensorLoad_0_io_tensor_rd_0_data_bits_0_4; // @[Load.scala 97:29]
  assign io_inp_rd_0_data_bits_0_5 = tensorLoad_0_io_tensor_rd_0_data_bits_0_5; // @[Load.scala 97:29]
  assign io_inp_rd_0_data_bits_0_6 = tensorLoad_0_io_tensor_rd_0_data_bits_0_6; // @[Load.scala 97:29]
  assign io_inp_rd_0_data_bits_0_7 = tensorLoad_0_io_tensor_rd_0_data_bits_0_7; // @[Load.scala 97:29]
  assign io_inp_rd_0_data_bits_0_8 = tensorLoad_0_io_tensor_rd_0_data_bits_0_8; // @[Load.scala 97:29]
  assign io_inp_rd_0_data_bits_0_9 = tensorLoad_0_io_tensor_rd_0_data_bits_0_9; // @[Load.scala 97:29]
  assign io_inp_rd_0_data_bits_0_10 = tensorLoad_0_io_tensor_rd_0_data_bits_0_10; // @[Load.scala 97:29]
  assign io_inp_rd_0_data_bits_0_11 = tensorLoad_0_io_tensor_rd_0_data_bits_0_11; // @[Load.scala 97:29]
  assign io_inp_rd_0_data_bits_0_12 = tensorLoad_0_io_tensor_rd_0_data_bits_0_12; // @[Load.scala 97:29]
  assign io_inp_rd_0_data_bits_0_13 = tensorLoad_0_io_tensor_rd_0_data_bits_0_13; // @[Load.scala 97:29]
  assign io_inp_rd_0_data_bits_0_14 = tensorLoad_0_io_tensor_rd_0_data_bits_0_14; // @[Load.scala 97:29]
  assign io_inp_rd_0_data_bits_0_15 = tensorLoad_0_io_tensor_rd_0_data_bits_0_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_valid = tensorLoad_1_io_tensor_rd_0_data_valid; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_0_0 = tensorLoad_1_io_tensor_rd_0_data_bits_0_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_0_1 = tensorLoad_1_io_tensor_rd_0_data_bits_0_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_0_2 = tensorLoad_1_io_tensor_rd_0_data_bits_0_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_0_3 = tensorLoad_1_io_tensor_rd_0_data_bits_0_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_0_4 = tensorLoad_1_io_tensor_rd_0_data_bits_0_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_0_5 = tensorLoad_1_io_tensor_rd_0_data_bits_0_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_0_6 = tensorLoad_1_io_tensor_rd_0_data_bits_0_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_0_7 = tensorLoad_1_io_tensor_rd_0_data_bits_0_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_0_8 = tensorLoad_1_io_tensor_rd_0_data_bits_0_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_0_9 = tensorLoad_1_io_tensor_rd_0_data_bits_0_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_0_10 = tensorLoad_1_io_tensor_rd_0_data_bits_0_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_0_11 = tensorLoad_1_io_tensor_rd_0_data_bits_0_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_0_12 = tensorLoad_1_io_tensor_rd_0_data_bits_0_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_0_13 = tensorLoad_1_io_tensor_rd_0_data_bits_0_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_0_14 = tensorLoad_1_io_tensor_rd_0_data_bits_0_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_0_15 = tensorLoad_1_io_tensor_rd_0_data_bits_0_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_1_0 = tensorLoad_1_io_tensor_rd_0_data_bits_1_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_1_1 = tensorLoad_1_io_tensor_rd_0_data_bits_1_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_1_2 = tensorLoad_1_io_tensor_rd_0_data_bits_1_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_1_3 = tensorLoad_1_io_tensor_rd_0_data_bits_1_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_1_4 = tensorLoad_1_io_tensor_rd_0_data_bits_1_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_1_5 = tensorLoad_1_io_tensor_rd_0_data_bits_1_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_1_6 = tensorLoad_1_io_tensor_rd_0_data_bits_1_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_1_7 = tensorLoad_1_io_tensor_rd_0_data_bits_1_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_1_8 = tensorLoad_1_io_tensor_rd_0_data_bits_1_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_1_9 = tensorLoad_1_io_tensor_rd_0_data_bits_1_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_1_10 = tensorLoad_1_io_tensor_rd_0_data_bits_1_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_1_11 = tensorLoad_1_io_tensor_rd_0_data_bits_1_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_1_12 = tensorLoad_1_io_tensor_rd_0_data_bits_1_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_1_13 = tensorLoad_1_io_tensor_rd_0_data_bits_1_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_1_14 = tensorLoad_1_io_tensor_rd_0_data_bits_1_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_1_15 = tensorLoad_1_io_tensor_rd_0_data_bits_1_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_2_0 = tensorLoad_1_io_tensor_rd_0_data_bits_2_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_2_1 = tensorLoad_1_io_tensor_rd_0_data_bits_2_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_2_2 = tensorLoad_1_io_tensor_rd_0_data_bits_2_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_2_3 = tensorLoad_1_io_tensor_rd_0_data_bits_2_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_2_4 = tensorLoad_1_io_tensor_rd_0_data_bits_2_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_2_5 = tensorLoad_1_io_tensor_rd_0_data_bits_2_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_2_6 = tensorLoad_1_io_tensor_rd_0_data_bits_2_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_2_7 = tensorLoad_1_io_tensor_rd_0_data_bits_2_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_2_8 = tensorLoad_1_io_tensor_rd_0_data_bits_2_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_2_9 = tensorLoad_1_io_tensor_rd_0_data_bits_2_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_2_10 = tensorLoad_1_io_tensor_rd_0_data_bits_2_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_2_11 = tensorLoad_1_io_tensor_rd_0_data_bits_2_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_2_12 = tensorLoad_1_io_tensor_rd_0_data_bits_2_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_2_13 = tensorLoad_1_io_tensor_rd_0_data_bits_2_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_2_14 = tensorLoad_1_io_tensor_rd_0_data_bits_2_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_2_15 = tensorLoad_1_io_tensor_rd_0_data_bits_2_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_3_0 = tensorLoad_1_io_tensor_rd_0_data_bits_3_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_3_1 = tensorLoad_1_io_tensor_rd_0_data_bits_3_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_3_2 = tensorLoad_1_io_tensor_rd_0_data_bits_3_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_3_3 = tensorLoad_1_io_tensor_rd_0_data_bits_3_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_3_4 = tensorLoad_1_io_tensor_rd_0_data_bits_3_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_3_5 = tensorLoad_1_io_tensor_rd_0_data_bits_3_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_3_6 = tensorLoad_1_io_tensor_rd_0_data_bits_3_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_3_7 = tensorLoad_1_io_tensor_rd_0_data_bits_3_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_3_8 = tensorLoad_1_io_tensor_rd_0_data_bits_3_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_3_9 = tensorLoad_1_io_tensor_rd_0_data_bits_3_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_3_10 = tensorLoad_1_io_tensor_rd_0_data_bits_3_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_3_11 = tensorLoad_1_io_tensor_rd_0_data_bits_3_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_3_12 = tensorLoad_1_io_tensor_rd_0_data_bits_3_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_3_13 = tensorLoad_1_io_tensor_rd_0_data_bits_3_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_3_14 = tensorLoad_1_io_tensor_rd_0_data_bits_3_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_3_15 = tensorLoad_1_io_tensor_rd_0_data_bits_3_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_4_0 = tensorLoad_1_io_tensor_rd_0_data_bits_4_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_4_1 = tensorLoad_1_io_tensor_rd_0_data_bits_4_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_4_2 = tensorLoad_1_io_tensor_rd_0_data_bits_4_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_4_3 = tensorLoad_1_io_tensor_rd_0_data_bits_4_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_4_4 = tensorLoad_1_io_tensor_rd_0_data_bits_4_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_4_5 = tensorLoad_1_io_tensor_rd_0_data_bits_4_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_4_6 = tensorLoad_1_io_tensor_rd_0_data_bits_4_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_4_7 = tensorLoad_1_io_tensor_rd_0_data_bits_4_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_4_8 = tensorLoad_1_io_tensor_rd_0_data_bits_4_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_4_9 = tensorLoad_1_io_tensor_rd_0_data_bits_4_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_4_10 = tensorLoad_1_io_tensor_rd_0_data_bits_4_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_4_11 = tensorLoad_1_io_tensor_rd_0_data_bits_4_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_4_12 = tensorLoad_1_io_tensor_rd_0_data_bits_4_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_4_13 = tensorLoad_1_io_tensor_rd_0_data_bits_4_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_4_14 = tensorLoad_1_io_tensor_rd_0_data_bits_4_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_4_15 = tensorLoad_1_io_tensor_rd_0_data_bits_4_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_5_0 = tensorLoad_1_io_tensor_rd_0_data_bits_5_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_5_1 = tensorLoad_1_io_tensor_rd_0_data_bits_5_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_5_2 = tensorLoad_1_io_tensor_rd_0_data_bits_5_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_5_3 = tensorLoad_1_io_tensor_rd_0_data_bits_5_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_5_4 = tensorLoad_1_io_tensor_rd_0_data_bits_5_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_5_5 = tensorLoad_1_io_tensor_rd_0_data_bits_5_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_5_6 = tensorLoad_1_io_tensor_rd_0_data_bits_5_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_5_7 = tensorLoad_1_io_tensor_rd_0_data_bits_5_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_5_8 = tensorLoad_1_io_tensor_rd_0_data_bits_5_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_5_9 = tensorLoad_1_io_tensor_rd_0_data_bits_5_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_5_10 = tensorLoad_1_io_tensor_rd_0_data_bits_5_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_5_11 = tensorLoad_1_io_tensor_rd_0_data_bits_5_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_5_12 = tensorLoad_1_io_tensor_rd_0_data_bits_5_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_5_13 = tensorLoad_1_io_tensor_rd_0_data_bits_5_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_5_14 = tensorLoad_1_io_tensor_rd_0_data_bits_5_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_5_15 = tensorLoad_1_io_tensor_rd_0_data_bits_5_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_6_0 = tensorLoad_1_io_tensor_rd_0_data_bits_6_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_6_1 = tensorLoad_1_io_tensor_rd_0_data_bits_6_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_6_2 = tensorLoad_1_io_tensor_rd_0_data_bits_6_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_6_3 = tensorLoad_1_io_tensor_rd_0_data_bits_6_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_6_4 = tensorLoad_1_io_tensor_rd_0_data_bits_6_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_6_5 = tensorLoad_1_io_tensor_rd_0_data_bits_6_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_6_6 = tensorLoad_1_io_tensor_rd_0_data_bits_6_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_6_7 = tensorLoad_1_io_tensor_rd_0_data_bits_6_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_6_8 = tensorLoad_1_io_tensor_rd_0_data_bits_6_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_6_9 = tensorLoad_1_io_tensor_rd_0_data_bits_6_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_6_10 = tensorLoad_1_io_tensor_rd_0_data_bits_6_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_6_11 = tensorLoad_1_io_tensor_rd_0_data_bits_6_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_6_12 = tensorLoad_1_io_tensor_rd_0_data_bits_6_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_6_13 = tensorLoad_1_io_tensor_rd_0_data_bits_6_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_6_14 = tensorLoad_1_io_tensor_rd_0_data_bits_6_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_6_15 = tensorLoad_1_io_tensor_rd_0_data_bits_6_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_7_0 = tensorLoad_1_io_tensor_rd_0_data_bits_7_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_7_1 = tensorLoad_1_io_tensor_rd_0_data_bits_7_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_7_2 = tensorLoad_1_io_tensor_rd_0_data_bits_7_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_7_3 = tensorLoad_1_io_tensor_rd_0_data_bits_7_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_7_4 = tensorLoad_1_io_tensor_rd_0_data_bits_7_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_7_5 = tensorLoad_1_io_tensor_rd_0_data_bits_7_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_7_6 = tensorLoad_1_io_tensor_rd_0_data_bits_7_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_7_7 = tensorLoad_1_io_tensor_rd_0_data_bits_7_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_7_8 = tensorLoad_1_io_tensor_rd_0_data_bits_7_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_7_9 = tensorLoad_1_io_tensor_rd_0_data_bits_7_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_7_10 = tensorLoad_1_io_tensor_rd_0_data_bits_7_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_7_11 = tensorLoad_1_io_tensor_rd_0_data_bits_7_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_7_12 = tensorLoad_1_io_tensor_rd_0_data_bits_7_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_7_13 = tensorLoad_1_io_tensor_rd_0_data_bits_7_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_7_14 = tensorLoad_1_io_tensor_rd_0_data_bits_7_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_7_15 = tensorLoad_1_io_tensor_rd_0_data_bits_7_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_8_0 = tensorLoad_1_io_tensor_rd_0_data_bits_8_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_8_1 = tensorLoad_1_io_tensor_rd_0_data_bits_8_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_8_2 = tensorLoad_1_io_tensor_rd_0_data_bits_8_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_8_3 = tensorLoad_1_io_tensor_rd_0_data_bits_8_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_8_4 = tensorLoad_1_io_tensor_rd_0_data_bits_8_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_8_5 = tensorLoad_1_io_tensor_rd_0_data_bits_8_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_8_6 = tensorLoad_1_io_tensor_rd_0_data_bits_8_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_8_7 = tensorLoad_1_io_tensor_rd_0_data_bits_8_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_8_8 = tensorLoad_1_io_tensor_rd_0_data_bits_8_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_8_9 = tensorLoad_1_io_tensor_rd_0_data_bits_8_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_8_10 = tensorLoad_1_io_tensor_rd_0_data_bits_8_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_8_11 = tensorLoad_1_io_tensor_rd_0_data_bits_8_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_8_12 = tensorLoad_1_io_tensor_rd_0_data_bits_8_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_8_13 = tensorLoad_1_io_tensor_rd_0_data_bits_8_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_8_14 = tensorLoad_1_io_tensor_rd_0_data_bits_8_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_8_15 = tensorLoad_1_io_tensor_rd_0_data_bits_8_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_9_0 = tensorLoad_1_io_tensor_rd_0_data_bits_9_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_9_1 = tensorLoad_1_io_tensor_rd_0_data_bits_9_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_9_2 = tensorLoad_1_io_tensor_rd_0_data_bits_9_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_9_3 = tensorLoad_1_io_tensor_rd_0_data_bits_9_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_9_4 = tensorLoad_1_io_tensor_rd_0_data_bits_9_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_9_5 = tensorLoad_1_io_tensor_rd_0_data_bits_9_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_9_6 = tensorLoad_1_io_tensor_rd_0_data_bits_9_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_9_7 = tensorLoad_1_io_tensor_rd_0_data_bits_9_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_9_8 = tensorLoad_1_io_tensor_rd_0_data_bits_9_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_9_9 = tensorLoad_1_io_tensor_rd_0_data_bits_9_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_9_10 = tensorLoad_1_io_tensor_rd_0_data_bits_9_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_9_11 = tensorLoad_1_io_tensor_rd_0_data_bits_9_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_9_12 = tensorLoad_1_io_tensor_rd_0_data_bits_9_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_9_13 = tensorLoad_1_io_tensor_rd_0_data_bits_9_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_9_14 = tensorLoad_1_io_tensor_rd_0_data_bits_9_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_9_15 = tensorLoad_1_io_tensor_rd_0_data_bits_9_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_10_0 = tensorLoad_1_io_tensor_rd_0_data_bits_10_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_10_1 = tensorLoad_1_io_tensor_rd_0_data_bits_10_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_10_2 = tensorLoad_1_io_tensor_rd_0_data_bits_10_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_10_3 = tensorLoad_1_io_tensor_rd_0_data_bits_10_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_10_4 = tensorLoad_1_io_tensor_rd_0_data_bits_10_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_10_5 = tensorLoad_1_io_tensor_rd_0_data_bits_10_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_10_6 = tensorLoad_1_io_tensor_rd_0_data_bits_10_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_10_7 = tensorLoad_1_io_tensor_rd_0_data_bits_10_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_10_8 = tensorLoad_1_io_tensor_rd_0_data_bits_10_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_10_9 = tensorLoad_1_io_tensor_rd_0_data_bits_10_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_10_10 = tensorLoad_1_io_tensor_rd_0_data_bits_10_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_10_11 = tensorLoad_1_io_tensor_rd_0_data_bits_10_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_10_12 = tensorLoad_1_io_tensor_rd_0_data_bits_10_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_10_13 = tensorLoad_1_io_tensor_rd_0_data_bits_10_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_10_14 = tensorLoad_1_io_tensor_rd_0_data_bits_10_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_10_15 = tensorLoad_1_io_tensor_rd_0_data_bits_10_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_11_0 = tensorLoad_1_io_tensor_rd_0_data_bits_11_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_11_1 = tensorLoad_1_io_tensor_rd_0_data_bits_11_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_11_2 = tensorLoad_1_io_tensor_rd_0_data_bits_11_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_11_3 = tensorLoad_1_io_tensor_rd_0_data_bits_11_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_11_4 = tensorLoad_1_io_tensor_rd_0_data_bits_11_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_11_5 = tensorLoad_1_io_tensor_rd_0_data_bits_11_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_11_6 = tensorLoad_1_io_tensor_rd_0_data_bits_11_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_11_7 = tensorLoad_1_io_tensor_rd_0_data_bits_11_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_11_8 = tensorLoad_1_io_tensor_rd_0_data_bits_11_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_11_9 = tensorLoad_1_io_tensor_rd_0_data_bits_11_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_11_10 = tensorLoad_1_io_tensor_rd_0_data_bits_11_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_11_11 = tensorLoad_1_io_tensor_rd_0_data_bits_11_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_11_12 = tensorLoad_1_io_tensor_rd_0_data_bits_11_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_11_13 = tensorLoad_1_io_tensor_rd_0_data_bits_11_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_11_14 = tensorLoad_1_io_tensor_rd_0_data_bits_11_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_11_15 = tensorLoad_1_io_tensor_rd_0_data_bits_11_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_12_0 = tensorLoad_1_io_tensor_rd_0_data_bits_12_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_12_1 = tensorLoad_1_io_tensor_rd_0_data_bits_12_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_12_2 = tensorLoad_1_io_tensor_rd_0_data_bits_12_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_12_3 = tensorLoad_1_io_tensor_rd_0_data_bits_12_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_12_4 = tensorLoad_1_io_tensor_rd_0_data_bits_12_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_12_5 = tensorLoad_1_io_tensor_rd_0_data_bits_12_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_12_6 = tensorLoad_1_io_tensor_rd_0_data_bits_12_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_12_7 = tensorLoad_1_io_tensor_rd_0_data_bits_12_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_12_8 = tensorLoad_1_io_tensor_rd_0_data_bits_12_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_12_9 = tensorLoad_1_io_tensor_rd_0_data_bits_12_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_12_10 = tensorLoad_1_io_tensor_rd_0_data_bits_12_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_12_11 = tensorLoad_1_io_tensor_rd_0_data_bits_12_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_12_12 = tensorLoad_1_io_tensor_rd_0_data_bits_12_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_12_13 = tensorLoad_1_io_tensor_rd_0_data_bits_12_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_12_14 = tensorLoad_1_io_tensor_rd_0_data_bits_12_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_12_15 = tensorLoad_1_io_tensor_rd_0_data_bits_12_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_13_0 = tensorLoad_1_io_tensor_rd_0_data_bits_13_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_13_1 = tensorLoad_1_io_tensor_rd_0_data_bits_13_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_13_2 = tensorLoad_1_io_tensor_rd_0_data_bits_13_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_13_3 = tensorLoad_1_io_tensor_rd_0_data_bits_13_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_13_4 = tensorLoad_1_io_tensor_rd_0_data_bits_13_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_13_5 = tensorLoad_1_io_tensor_rd_0_data_bits_13_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_13_6 = tensorLoad_1_io_tensor_rd_0_data_bits_13_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_13_7 = tensorLoad_1_io_tensor_rd_0_data_bits_13_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_13_8 = tensorLoad_1_io_tensor_rd_0_data_bits_13_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_13_9 = tensorLoad_1_io_tensor_rd_0_data_bits_13_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_13_10 = tensorLoad_1_io_tensor_rd_0_data_bits_13_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_13_11 = tensorLoad_1_io_tensor_rd_0_data_bits_13_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_13_12 = tensorLoad_1_io_tensor_rd_0_data_bits_13_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_13_13 = tensorLoad_1_io_tensor_rd_0_data_bits_13_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_13_14 = tensorLoad_1_io_tensor_rd_0_data_bits_13_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_13_15 = tensorLoad_1_io_tensor_rd_0_data_bits_13_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_14_0 = tensorLoad_1_io_tensor_rd_0_data_bits_14_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_14_1 = tensorLoad_1_io_tensor_rd_0_data_bits_14_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_14_2 = tensorLoad_1_io_tensor_rd_0_data_bits_14_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_14_3 = tensorLoad_1_io_tensor_rd_0_data_bits_14_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_14_4 = tensorLoad_1_io_tensor_rd_0_data_bits_14_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_14_5 = tensorLoad_1_io_tensor_rd_0_data_bits_14_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_14_6 = tensorLoad_1_io_tensor_rd_0_data_bits_14_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_14_7 = tensorLoad_1_io_tensor_rd_0_data_bits_14_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_14_8 = tensorLoad_1_io_tensor_rd_0_data_bits_14_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_14_9 = tensorLoad_1_io_tensor_rd_0_data_bits_14_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_14_10 = tensorLoad_1_io_tensor_rd_0_data_bits_14_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_14_11 = tensorLoad_1_io_tensor_rd_0_data_bits_14_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_14_12 = tensorLoad_1_io_tensor_rd_0_data_bits_14_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_14_13 = tensorLoad_1_io_tensor_rd_0_data_bits_14_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_14_14 = tensorLoad_1_io_tensor_rd_0_data_bits_14_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_14_15 = tensorLoad_1_io_tensor_rd_0_data_bits_14_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_15_0 = tensorLoad_1_io_tensor_rd_0_data_bits_15_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_15_1 = tensorLoad_1_io_tensor_rd_0_data_bits_15_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_15_2 = tensorLoad_1_io_tensor_rd_0_data_bits_15_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_15_3 = tensorLoad_1_io_tensor_rd_0_data_bits_15_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_15_4 = tensorLoad_1_io_tensor_rd_0_data_bits_15_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_15_5 = tensorLoad_1_io_tensor_rd_0_data_bits_15_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_15_6 = tensorLoad_1_io_tensor_rd_0_data_bits_15_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_15_7 = tensorLoad_1_io_tensor_rd_0_data_bits_15_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_15_8 = tensorLoad_1_io_tensor_rd_0_data_bits_15_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_15_9 = tensorLoad_1_io_tensor_rd_0_data_bits_15_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_15_10 = tensorLoad_1_io_tensor_rd_0_data_bits_15_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_15_11 = tensorLoad_1_io_tensor_rd_0_data_bits_15_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_15_12 = tensorLoad_1_io_tensor_rd_0_data_bits_15_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_15_13 = tensorLoad_1_io_tensor_rd_0_data_bits_15_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_15_14 = tensorLoad_1_io_tensor_rd_0_data_bits_15_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_15_15 = tensorLoad_1_io_tensor_rd_0_data_bits_15_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_16_0 = tensorLoad_1_io_tensor_rd_0_data_bits_16_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_16_1 = tensorLoad_1_io_tensor_rd_0_data_bits_16_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_16_2 = tensorLoad_1_io_tensor_rd_0_data_bits_16_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_16_3 = tensorLoad_1_io_tensor_rd_0_data_bits_16_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_16_4 = tensorLoad_1_io_tensor_rd_0_data_bits_16_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_16_5 = tensorLoad_1_io_tensor_rd_0_data_bits_16_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_16_6 = tensorLoad_1_io_tensor_rd_0_data_bits_16_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_16_7 = tensorLoad_1_io_tensor_rd_0_data_bits_16_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_16_8 = tensorLoad_1_io_tensor_rd_0_data_bits_16_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_16_9 = tensorLoad_1_io_tensor_rd_0_data_bits_16_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_16_10 = tensorLoad_1_io_tensor_rd_0_data_bits_16_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_16_11 = tensorLoad_1_io_tensor_rd_0_data_bits_16_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_16_12 = tensorLoad_1_io_tensor_rd_0_data_bits_16_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_16_13 = tensorLoad_1_io_tensor_rd_0_data_bits_16_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_16_14 = tensorLoad_1_io_tensor_rd_0_data_bits_16_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_16_15 = tensorLoad_1_io_tensor_rd_0_data_bits_16_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_17_0 = tensorLoad_1_io_tensor_rd_0_data_bits_17_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_17_1 = tensorLoad_1_io_tensor_rd_0_data_bits_17_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_17_2 = tensorLoad_1_io_tensor_rd_0_data_bits_17_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_17_3 = tensorLoad_1_io_tensor_rd_0_data_bits_17_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_17_4 = tensorLoad_1_io_tensor_rd_0_data_bits_17_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_17_5 = tensorLoad_1_io_tensor_rd_0_data_bits_17_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_17_6 = tensorLoad_1_io_tensor_rd_0_data_bits_17_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_17_7 = tensorLoad_1_io_tensor_rd_0_data_bits_17_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_17_8 = tensorLoad_1_io_tensor_rd_0_data_bits_17_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_17_9 = tensorLoad_1_io_tensor_rd_0_data_bits_17_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_17_10 = tensorLoad_1_io_tensor_rd_0_data_bits_17_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_17_11 = tensorLoad_1_io_tensor_rd_0_data_bits_17_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_17_12 = tensorLoad_1_io_tensor_rd_0_data_bits_17_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_17_13 = tensorLoad_1_io_tensor_rd_0_data_bits_17_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_17_14 = tensorLoad_1_io_tensor_rd_0_data_bits_17_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_17_15 = tensorLoad_1_io_tensor_rd_0_data_bits_17_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_18_0 = tensorLoad_1_io_tensor_rd_0_data_bits_18_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_18_1 = tensorLoad_1_io_tensor_rd_0_data_bits_18_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_18_2 = tensorLoad_1_io_tensor_rd_0_data_bits_18_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_18_3 = tensorLoad_1_io_tensor_rd_0_data_bits_18_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_18_4 = tensorLoad_1_io_tensor_rd_0_data_bits_18_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_18_5 = tensorLoad_1_io_tensor_rd_0_data_bits_18_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_18_6 = tensorLoad_1_io_tensor_rd_0_data_bits_18_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_18_7 = tensorLoad_1_io_tensor_rd_0_data_bits_18_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_18_8 = tensorLoad_1_io_tensor_rd_0_data_bits_18_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_18_9 = tensorLoad_1_io_tensor_rd_0_data_bits_18_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_18_10 = tensorLoad_1_io_tensor_rd_0_data_bits_18_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_18_11 = tensorLoad_1_io_tensor_rd_0_data_bits_18_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_18_12 = tensorLoad_1_io_tensor_rd_0_data_bits_18_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_18_13 = tensorLoad_1_io_tensor_rd_0_data_bits_18_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_18_14 = tensorLoad_1_io_tensor_rd_0_data_bits_18_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_18_15 = tensorLoad_1_io_tensor_rd_0_data_bits_18_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_19_0 = tensorLoad_1_io_tensor_rd_0_data_bits_19_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_19_1 = tensorLoad_1_io_tensor_rd_0_data_bits_19_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_19_2 = tensorLoad_1_io_tensor_rd_0_data_bits_19_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_19_3 = tensorLoad_1_io_tensor_rd_0_data_bits_19_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_19_4 = tensorLoad_1_io_tensor_rd_0_data_bits_19_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_19_5 = tensorLoad_1_io_tensor_rd_0_data_bits_19_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_19_6 = tensorLoad_1_io_tensor_rd_0_data_bits_19_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_19_7 = tensorLoad_1_io_tensor_rd_0_data_bits_19_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_19_8 = tensorLoad_1_io_tensor_rd_0_data_bits_19_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_19_9 = tensorLoad_1_io_tensor_rd_0_data_bits_19_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_19_10 = tensorLoad_1_io_tensor_rd_0_data_bits_19_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_19_11 = tensorLoad_1_io_tensor_rd_0_data_bits_19_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_19_12 = tensorLoad_1_io_tensor_rd_0_data_bits_19_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_19_13 = tensorLoad_1_io_tensor_rd_0_data_bits_19_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_19_14 = tensorLoad_1_io_tensor_rd_0_data_bits_19_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_19_15 = tensorLoad_1_io_tensor_rd_0_data_bits_19_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_20_0 = tensorLoad_1_io_tensor_rd_0_data_bits_20_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_20_1 = tensorLoad_1_io_tensor_rd_0_data_bits_20_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_20_2 = tensorLoad_1_io_tensor_rd_0_data_bits_20_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_20_3 = tensorLoad_1_io_tensor_rd_0_data_bits_20_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_20_4 = tensorLoad_1_io_tensor_rd_0_data_bits_20_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_20_5 = tensorLoad_1_io_tensor_rd_0_data_bits_20_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_20_6 = tensorLoad_1_io_tensor_rd_0_data_bits_20_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_20_7 = tensorLoad_1_io_tensor_rd_0_data_bits_20_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_20_8 = tensorLoad_1_io_tensor_rd_0_data_bits_20_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_20_9 = tensorLoad_1_io_tensor_rd_0_data_bits_20_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_20_10 = tensorLoad_1_io_tensor_rd_0_data_bits_20_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_20_11 = tensorLoad_1_io_tensor_rd_0_data_bits_20_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_20_12 = tensorLoad_1_io_tensor_rd_0_data_bits_20_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_20_13 = tensorLoad_1_io_tensor_rd_0_data_bits_20_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_20_14 = tensorLoad_1_io_tensor_rd_0_data_bits_20_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_20_15 = tensorLoad_1_io_tensor_rd_0_data_bits_20_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_21_0 = tensorLoad_1_io_tensor_rd_0_data_bits_21_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_21_1 = tensorLoad_1_io_tensor_rd_0_data_bits_21_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_21_2 = tensorLoad_1_io_tensor_rd_0_data_bits_21_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_21_3 = tensorLoad_1_io_tensor_rd_0_data_bits_21_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_21_4 = tensorLoad_1_io_tensor_rd_0_data_bits_21_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_21_5 = tensorLoad_1_io_tensor_rd_0_data_bits_21_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_21_6 = tensorLoad_1_io_tensor_rd_0_data_bits_21_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_21_7 = tensorLoad_1_io_tensor_rd_0_data_bits_21_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_21_8 = tensorLoad_1_io_tensor_rd_0_data_bits_21_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_21_9 = tensorLoad_1_io_tensor_rd_0_data_bits_21_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_21_10 = tensorLoad_1_io_tensor_rd_0_data_bits_21_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_21_11 = tensorLoad_1_io_tensor_rd_0_data_bits_21_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_21_12 = tensorLoad_1_io_tensor_rd_0_data_bits_21_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_21_13 = tensorLoad_1_io_tensor_rd_0_data_bits_21_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_21_14 = tensorLoad_1_io_tensor_rd_0_data_bits_21_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_21_15 = tensorLoad_1_io_tensor_rd_0_data_bits_21_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_22_0 = tensorLoad_1_io_tensor_rd_0_data_bits_22_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_22_1 = tensorLoad_1_io_tensor_rd_0_data_bits_22_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_22_2 = tensorLoad_1_io_tensor_rd_0_data_bits_22_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_22_3 = tensorLoad_1_io_tensor_rd_0_data_bits_22_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_22_4 = tensorLoad_1_io_tensor_rd_0_data_bits_22_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_22_5 = tensorLoad_1_io_tensor_rd_0_data_bits_22_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_22_6 = tensorLoad_1_io_tensor_rd_0_data_bits_22_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_22_7 = tensorLoad_1_io_tensor_rd_0_data_bits_22_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_22_8 = tensorLoad_1_io_tensor_rd_0_data_bits_22_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_22_9 = tensorLoad_1_io_tensor_rd_0_data_bits_22_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_22_10 = tensorLoad_1_io_tensor_rd_0_data_bits_22_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_22_11 = tensorLoad_1_io_tensor_rd_0_data_bits_22_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_22_12 = tensorLoad_1_io_tensor_rd_0_data_bits_22_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_22_13 = tensorLoad_1_io_tensor_rd_0_data_bits_22_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_22_14 = tensorLoad_1_io_tensor_rd_0_data_bits_22_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_22_15 = tensorLoad_1_io_tensor_rd_0_data_bits_22_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_23_0 = tensorLoad_1_io_tensor_rd_0_data_bits_23_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_23_1 = tensorLoad_1_io_tensor_rd_0_data_bits_23_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_23_2 = tensorLoad_1_io_tensor_rd_0_data_bits_23_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_23_3 = tensorLoad_1_io_tensor_rd_0_data_bits_23_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_23_4 = tensorLoad_1_io_tensor_rd_0_data_bits_23_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_23_5 = tensorLoad_1_io_tensor_rd_0_data_bits_23_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_23_6 = tensorLoad_1_io_tensor_rd_0_data_bits_23_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_23_7 = tensorLoad_1_io_tensor_rd_0_data_bits_23_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_23_8 = tensorLoad_1_io_tensor_rd_0_data_bits_23_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_23_9 = tensorLoad_1_io_tensor_rd_0_data_bits_23_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_23_10 = tensorLoad_1_io_tensor_rd_0_data_bits_23_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_23_11 = tensorLoad_1_io_tensor_rd_0_data_bits_23_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_23_12 = tensorLoad_1_io_tensor_rd_0_data_bits_23_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_23_13 = tensorLoad_1_io_tensor_rd_0_data_bits_23_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_23_14 = tensorLoad_1_io_tensor_rd_0_data_bits_23_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_23_15 = tensorLoad_1_io_tensor_rd_0_data_bits_23_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_24_0 = tensorLoad_1_io_tensor_rd_0_data_bits_24_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_24_1 = tensorLoad_1_io_tensor_rd_0_data_bits_24_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_24_2 = tensorLoad_1_io_tensor_rd_0_data_bits_24_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_24_3 = tensorLoad_1_io_tensor_rd_0_data_bits_24_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_24_4 = tensorLoad_1_io_tensor_rd_0_data_bits_24_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_24_5 = tensorLoad_1_io_tensor_rd_0_data_bits_24_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_24_6 = tensorLoad_1_io_tensor_rd_0_data_bits_24_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_24_7 = tensorLoad_1_io_tensor_rd_0_data_bits_24_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_24_8 = tensorLoad_1_io_tensor_rd_0_data_bits_24_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_24_9 = tensorLoad_1_io_tensor_rd_0_data_bits_24_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_24_10 = tensorLoad_1_io_tensor_rd_0_data_bits_24_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_24_11 = tensorLoad_1_io_tensor_rd_0_data_bits_24_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_24_12 = tensorLoad_1_io_tensor_rd_0_data_bits_24_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_24_13 = tensorLoad_1_io_tensor_rd_0_data_bits_24_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_24_14 = tensorLoad_1_io_tensor_rd_0_data_bits_24_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_24_15 = tensorLoad_1_io_tensor_rd_0_data_bits_24_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_25_0 = tensorLoad_1_io_tensor_rd_0_data_bits_25_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_25_1 = tensorLoad_1_io_tensor_rd_0_data_bits_25_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_25_2 = tensorLoad_1_io_tensor_rd_0_data_bits_25_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_25_3 = tensorLoad_1_io_tensor_rd_0_data_bits_25_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_25_4 = tensorLoad_1_io_tensor_rd_0_data_bits_25_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_25_5 = tensorLoad_1_io_tensor_rd_0_data_bits_25_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_25_6 = tensorLoad_1_io_tensor_rd_0_data_bits_25_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_25_7 = tensorLoad_1_io_tensor_rd_0_data_bits_25_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_25_8 = tensorLoad_1_io_tensor_rd_0_data_bits_25_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_25_9 = tensorLoad_1_io_tensor_rd_0_data_bits_25_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_25_10 = tensorLoad_1_io_tensor_rd_0_data_bits_25_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_25_11 = tensorLoad_1_io_tensor_rd_0_data_bits_25_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_25_12 = tensorLoad_1_io_tensor_rd_0_data_bits_25_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_25_13 = tensorLoad_1_io_tensor_rd_0_data_bits_25_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_25_14 = tensorLoad_1_io_tensor_rd_0_data_bits_25_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_25_15 = tensorLoad_1_io_tensor_rd_0_data_bits_25_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_26_0 = tensorLoad_1_io_tensor_rd_0_data_bits_26_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_26_1 = tensorLoad_1_io_tensor_rd_0_data_bits_26_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_26_2 = tensorLoad_1_io_tensor_rd_0_data_bits_26_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_26_3 = tensorLoad_1_io_tensor_rd_0_data_bits_26_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_26_4 = tensorLoad_1_io_tensor_rd_0_data_bits_26_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_26_5 = tensorLoad_1_io_tensor_rd_0_data_bits_26_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_26_6 = tensorLoad_1_io_tensor_rd_0_data_bits_26_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_26_7 = tensorLoad_1_io_tensor_rd_0_data_bits_26_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_26_8 = tensorLoad_1_io_tensor_rd_0_data_bits_26_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_26_9 = tensorLoad_1_io_tensor_rd_0_data_bits_26_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_26_10 = tensorLoad_1_io_tensor_rd_0_data_bits_26_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_26_11 = tensorLoad_1_io_tensor_rd_0_data_bits_26_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_26_12 = tensorLoad_1_io_tensor_rd_0_data_bits_26_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_26_13 = tensorLoad_1_io_tensor_rd_0_data_bits_26_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_26_14 = tensorLoad_1_io_tensor_rd_0_data_bits_26_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_26_15 = tensorLoad_1_io_tensor_rd_0_data_bits_26_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_27_0 = tensorLoad_1_io_tensor_rd_0_data_bits_27_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_27_1 = tensorLoad_1_io_tensor_rd_0_data_bits_27_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_27_2 = tensorLoad_1_io_tensor_rd_0_data_bits_27_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_27_3 = tensorLoad_1_io_tensor_rd_0_data_bits_27_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_27_4 = tensorLoad_1_io_tensor_rd_0_data_bits_27_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_27_5 = tensorLoad_1_io_tensor_rd_0_data_bits_27_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_27_6 = tensorLoad_1_io_tensor_rd_0_data_bits_27_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_27_7 = tensorLoad_1_io_tensor_rd_0_data_bits_27_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_27_8 = tensorLoad_1_io_tensor_rd_0_data_bits_27_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_27_9 = tensorLoad_1_io_tensor_rd_0_data_bits_27_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_27_10 = tensorLoad_1_io_tensor_rd_0_data_bits_27_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_27_11 = tensorLoad_1_io_tensor_rd_0_data_bits_27_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_27_12 = tensorLoad_1_io_tensor_rd_0_data_bits_27_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_27_13 = tensorLoad_1_io_tensor_rd_0_data_bits_27_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_27_14 = tensorLoad_1_io_tensor_rd_0_data_bits_27_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_27_15 = tensorLoad_1_io_tensor_rd_0_data_bits_27_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_28_0 = tensorLoad_1_io_tensor_rd_0_data_bits_28_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_28_1 = tensorLoad_1_io_tensor_rd_0_data_bits_28_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_28_2 = tensorLoad_1_io_tensor_rd_0_data_bits_28_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_28_3 = tensorLoad_1_io_tensor_rd_0_data_bits_28_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_28_4 = tensorLoad_1_io_tensor_rd_0_data_bits_28_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_28_5 = tensorLoad_1_io_tensor_rd_0_data_bits_28_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_28_6 = tensorLoad_1_io_tensor_rd_0_data_bits_28_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_28_7 = tensorLoad_1_io_tensor_rd_0_data_bits_28_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_28_8 = tensorLoad_1_io_tensor_rd_0_data_bits_28_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_28_9 = tensorLoad_1_io_tensor_rd_0_data_bits_28_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_28_10 = tensorLoad_1_io_tensor_rd_0_data_bits_28_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_28_11 = tensorLoad_1_io_tensor_rd_0_data_bits_28_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_28_12 = tensorLoad_1_io_tensor_rd_0_data_bits_28_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_28_13 = tensorLoad_1_io_tensor_rd_0_data_bits_28_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_28_14 = tensorLoad_1_io_tensor_rd_0_data_bits_28_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_28_15 = tensorLoad_1_io_tensor_rd_0_data_bits_28_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_29_0 = tensorLoad_1_io_tensor_rd_0_data_bits_29_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_29_1 = tensorLoad_1_io_tensor_rd_0_data_bits_29_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_29_2 = tensorLoad_1_io_tensor_rd_0_data_bits_29_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_29_3 = tensorLoad_1_io_tensor_rd_0_data_bits_29_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_29_4 = tensorLoad_1_io_tensor_rd_0_data_bits_29_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_29_5 = tensorLoad_1_io_tensor_rd_0_data_bits_29_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_29_6 = tensorLoad_1_io_tensor_rd_0_data_bits_29_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_29_7 = tensorLoad_1_io_tensor_rd_0_data_bits_29_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_29_8 = tensorLoad_1_io_tensor_rd_0_data_bits_29_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_29_9 = tensorLoad_1_io_tensor_rd_0_data_bits_29_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_29_10 = tensorLoad_1_io_tensor_rd_0_data_bits_29_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_29_11 = tensorLoad_1_io_tensor_rd_0_data_bits_29_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_29_12 = tensorLoad_1_io_tensor_rd_0_data_bits_29_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_29_13 = tensorLoad_1_io_tensor_rd_0_data_bits_29_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_29_14 = tensorLoad_1_io_tensor_rd_0_data_bits_29_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_29_15 = tensorLoad_1_io_tensor_rd_0_data_bits_29_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_30_0 = tensorLoad_1_io_tensor_rd_0_data_bits_30_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_30_1 = tensorLoad_1_io_tensor_rd_0_data_bits_30_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_30_2 = tensorLoad_1_io_tensor_rd_0_data_bits_30_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_30_3 = tensorLoad_1_io_tensor_rd_0_data_bits_30_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_30_4 = tensorLoad_1_io_tensor_rd_0_data_bits_30_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_30_5 = tensorLoad_1_io_tensor_rd_0_data_bits_30_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_30_6 = tensorLoad_1_io_tensor_rd_0_data_bits_30_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_30_7 = tensorLoad_1_io_tensor_rd_0_data_bits_30_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_30_8 = tensorLoad_1_io_tensor_rd_0_data_bits_30_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_30_9 = tensorLoad_1_io_tensor_rd_0_data_bits_30_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_30_10 = tensorLoad_1_io_tensor_rd_0_data_bits_30_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_30_11 = tensorLoad_1_io_tensor_rd_0_data_bits_30_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_30_12 = tensorLoad_1_io_tensor_rd_0_data_bits_30_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_30_13 = tensorLoad_1_io_tensor_rd_0_data_bits_30_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_30_14 = tensorLoad_1_io_tensor_rd_0_data_bits_30_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_30_15 = tensorLoad_1_io_tensor_rd_0_data_bits_30_15; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_31_0 = tensorLoad_1_io_tensor_rd_0_data_bits_31_0; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_31_1 = tensorLoad_1_io_tensor_rd_0_data_bits_31_1; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_31_2 = tensorLoad_1_io_tensor_rd_0_data_bits_31_2; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_31_3 = tensorLoad_1_io_tensor_rd_0_data_bits_31_3; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_31_4 = tensorLoad_1_io_tensor_rd_0_data_bits_31_4; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_31_5 = tensorLoad_1_io_tensor_rd_0_data_bits_31_5; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_31_6 = tensorLoad_1_io_tensor_rd_0_data_bits_31_6; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_31_7 = tensorLoad_1_io_tensor_rd_0_data_bits_31_7; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_31_8 = tensorLoad_1_io_tensor_rd_0_data_bits_31_8; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_31_9 = tensorLoad_1_io_tensor_rd_0_data_bits_31_9; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_31_10 = tensorLoad_1_io_tensor_rd_0_data_bits_31_10; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_31_11 = tensorLoad_1_io_tensor_rd_0_data_bits_31_11; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_31_12 = tensorLoad_1_io_tensor_rd_0_data_bits_31_12; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_31_13 = tensorLoad_1_io_tensor_rd_0_data_bits_31_13; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_31_14 = tensorLoad_1_io_tensor_rd_0_data_bits_31_14; // @[Load.scala 97:29]
  assign io_wgt_rd_0_data_bits_31_15 = tensorLoad_1_io_tensor_rd_0_data_bits_31_15; // @[Load.scala 97:29]
  assign s_clock = clock;
  assign s_reset = reset;
  assign s_io_spost = io_i_post; // @[Load.scala 102:14]
  assign s_io_swait = dec_io_pop_next & _tensorLoad_0_io_start_T_1; // @[Load.scala 103:33]
  assign inst_q_clock = clock;
  assign inst_q_reset = reset;
  assign inst_q_io_enq_valid = io_inst_valid; // @[Load.scala 85:17]
  assign inst_q_io_enq_bits = io_inst_bits; // @[Load.scala 85:17]
  assign inst_q_io_deq_ready = state == 2'h2 & done | state == 2'h1; // @[Load.scala 86:50]
  assign dec_io_inst = inst_q_io_deq_bits; // @[Load.scala 53:15]
  assign tensorLoad_0_clock = clock;
  assign tensorLoad_0_reset = reset;
  assign tensorLoad_0_io_start = state == 2'h0 & start & dec_io_isInput; // @[Load.scala 94:55]
  assign tensorLoad_0_io_inst = inst_q_io_deq_bits; // @[Load.scala 95:27]
  assign tensorLoad_0_io_baddr = io_inp_baddr; // @[Load.scala 96:28]
  assign tensorLoad_0_io_vme_rd_cmd_ready = io_vme_rd_0_cmd_ready; // @[Load.scala 98:18]
  assign tensorLoad_0_io_vme_rd_data_valid = io_vme_rd_0_data_valid; // @[Load.scala 98:18]
  assign tensorLoad_0_io_vme_rd_data_bits_data = io_vme_rd_0_data_bits_data; // @[Load.scala 98:18]
  assign tensorLoad_0_io_vme_rd_data_bits_tag = io_vme_rd_0_data_bits_tag; // @[Load.scala 98:18]
  assign tensorLoad_0_io_tensor_rd_0_idx_valid = io_inp_rd_0_idx_valid; // @[Load.scala 97:29]
  assign tensorLoad_0_io_tensor_rd_0_idx_bits = io_inp_rd_0_idx_bits; // @[Load.scala 97:29]
  assign tensorLoad_1_clock = clock;
  assign tensorLoad_1_reset = reset;
  assign tensorLoad_1_io_start = state == 2'h0 & start & dec_io_isWeight; // @[Load.scala 94:55]
  assign tensorLoad_1_io_inst = inst_q_io_deq_bits; // @[Load.scala 95:27]
  assign tensorLoad_1_io_baddr = io_wgt_baddr; // @[Load.scala 96:28]
  assign tensorLoad_1_io_vme_rd_cmd_ready = io_vme_rd_1_cmd_ready; // @[Load.scala 98:18]
  assign tensorLoad_1_io_vme_rd_data_valid = io_vme_rd_1_data_valid; // @[Load.scala 98:18]
  assign tensorLoad_1_io_vme_rd_data_bits_data = io_vme_rd_1_data_bits_data; // @[Load.scala 98:18]
  assign tensorLoad_1_io_vme_rd_data_bits_tag = io_vme_rd_1_data_bits_tag; // @[Load.scala 98:18]
  assign tensorLoad_1_io_tensor_rd_0_idx_valid = io_wgt_rd_0_idx_valid; // @[Load.scala 97:29]
  assign tensorLoad_1_io_tensor_rd_0_idx_bits = io_wgt_rd_0_idx_bits; // @[Load.scala 97:29]
  always @(posedge clock) begin
    if (reset) begin // @[Load.scala 47:22]
      state <= 2'h0; // @[Load.scala 47:22]
    end else if (2'h0 == state) begin // @[Load.scala 64:17]
      if (start) begin // @[Load.scala 66:19]
        if (dec_io_isSync) begin // @[Load.scala 67:29]
          state <= 2'h1; // @[Load.scala 68:17]
        end else begin
          state <= _GEN_0;
        end
      end
    end else if (2'h1 == state) begin // @[Load.scala 64:17]
      state <= 2'h0; // @[Load.scala 75:13]
    end else if (2'h2 == state) begin // @[Load.scala 64:17]
      state <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module GenVMECmdWide(
  input         clock,
  input         reset,
  input         io_start,
  input         io_isBusy,
  input         io_updateState,
  input  [31:0] io_baddr,
  output        io_vmeCmd_valid,
  output [31:0] io_vmeCmd_bits_addr,
  output [3:0]  io_vmeCmd_bits_len,
  output [20:0] io_vmeCmd_bits_tag,
  output [4:0]  io_readLen,
  output        io_done,
  input  [15:0] io_ysize,
  input  [15:0] io_xsize,
  input  [15:0] io_xstride,
  input  [31:0] io_dram_offset,
  input  [15:0] io_sram_offset,
  input  [3:0]  io_xpad_0,
  input  [3:0]  io_xpad_1,
  input  [3:0]  io_ypad_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] dramLineIdx; // @[TensorLoadWideVME.scala 501:24]
  wire [15:0] _dramLineIdx_T_1 = dramLineIdx + 16'h1; // @[TensorLoadWideVME.scala 505:32]
  reg [14:0] clReadIdx; // @[TensorLoadWideVME.scala 591:22]
  wire [17:0] rdLineBytes = {io_xsize, 2'h0}; // @[TensorLoadWideVME.scala 552:30]
  reg [31:0] rdLineElemBeginAddr; // @[TensorLoadWideVME.scala 520:32]
  wire [31:0] _GEN_0 = rdLineElemBeginAddr % 32'h8; // @[TensorLoadWideVME.scala 562:51]
  wire [3:0] rd1stPulseOffsetBytes = _GEN_0[3:0]; // @[TensorLoadWideVME.scala 562:51]
  wire [17:0] _GEN_30 = {{14'd0}, rd1stPulseOffsetBytes}; // @[TensorLoadWideVME.scala 570:22]
  wire [17:0] _rdLineClNb_T_1 = rdLineBytes + _GEN_30; // @[TensorLoadWideVME.scala 570:22]
  wire [17:0] _GEN_1 = _rdLineClNb_T_1 % 18'h8; // @[TensorLoadWideVME.scala 570:47]
  wire [3:0] _rdLineClNb_T_2 = _GEN_1[3:0]; // @[TensorLoadWideVME.scala 570:47]
  wire [14:0] rdLineClNbTmp = _rdLineClNb_T_1[17:3]; // @[TensorLoadWideVME.scala 568:61]
  wire [14:0] _rdLineClNb_T_5 = rdLineClNbTmp + 15'h1; // @[TensorLoadWideVME.scala 570:97]
  wire [14:0] rdLineClNb = _rdLineClNb_T_2 == 4'h0 ? rdLineClNbTmp : _rdLineClNb_T_5; // @[TensorLoadWideVME.scala 570:8]
  wire  newReadRow = clReadIdx == 15'h0; // @[TensorLoadWideVME.scala 592:30]
  wire [14:0] clRemained = rdLineClNb - clReadIdx; // @[TensorLoadWideVME.scala 642:31]
  wire [31:0] rdLineClBeginAddr = rdLineElemBeginAddr & 32'hfffffff8; // @[TensorLoadWideVME.scala 521:47]
  wire [31:0] _GEN_2 = rdLineClBeginAddr % 32'h80; // @[TensorLoadWideVME.scala 557:62]
  wire [7:0] _rdLen1stMaxTransBytes_T = _GEN_2[7:0]; // @[TensorLoadWideVME.scala 557:62]
  wire [7:0] rdLen1stMaxTransBytes = 8'h80 - _rdLen1stMaxTransBytes_T; // @[TensorLoadWideVME.scala 557:42]
  wire [4:0] rdLen1stMaxTransClNb = rdLen1stMaxTransBytes[7:3]; // @[TensorLoadWideVME.scala 559:52]
  wire [14:0] _GEN_32 = {{10'd0}, rdLen1stMaxTransClNb}; // @[TensorLoadWideVME.scala 644:21]
  wire [14:0] _GEN_16 = clRemained < _GEN_32 ? clRemained : {{10'd0}, rdLen1stMaxTransClNb}; // @[TensorLoadWideVME.scala 644:45 645:13 647:13]
  wire [14:0] _GEN_17 = clRemained < 15'h10 ? clRemained : 15'h10; // @[TensorLoadWideVME.scala 650:36 651:13 653:13]
  wire [14:0] _GEN_18 = newReadRow ? _GEN_16 : _GEN_17; // @[TensorLoadWideVME.scala 643:21]
  wire [4:0] rdLen = _GEN_18[4:0]; // @[TensorLoadWideVME.scala 537:19]
  wire [14:0] _GEN_33 = {{10'd0}, rdLen}; // @[TensorLoadWideVME.scala 635:34]
  wire [14:0] _T_28 = rdLineClNb - _GEN_33; // @[TensorLoadWideVME.scala 635:34]
  wire  _T_29 = clReadIdx == _T_28; // @[TensorLoadWideVME.scala 635:19]
  wire [15:0] _T_31 = io_ysize - 16'h1; // @[TensorLoadWideVME.scala 635:72]
  wire  stride = clReadIdx == _T_28 & dramLineIdx != _T_31 & io_updateState; // @[TensorLoadWideVME.scala 635:79]
  wire [33:0] _dramInitialAddr_T = {io_dram_offset, 2'h0}; // @[TensorLoadWideVME.scala 512:41]
  wire [31:0] dramInitialAddr = _dramInitialAddr_T[31:0]; // @[TensorLoadWideVME.scala 512:{73,73}]
  wire [31:0] xferElemInitAddr = io_baddr | dramInitialAddr; // @[TensorLoadWideVME.scala 513:35]
  wire [31:0] xferClInitAddr = xferElemInitAddr & 32'hfffffff8; // @[TensorLoadWideVME.scala 519:41]
  wire [17:0] _nextLineBeginElemAddr_T = {io_xstride, 2'h0}; // @[TensorLoadWideVME.scala 523:65]
  wire [31:0] _GEN_34 = {{14'd0}, _nextLineBeginElemAddr_T}; // @[TensorLoadWideVME.scala 523:51]
  wire [31:0] nextLineBeginElemAddr = rdLineElemBeginAddr + _GEN_34; // @[TensorLoadWideVME.scala 523:51]
  wire [31:0] nextLineBeginClAddr = nextLineBeginElemAddr & 32'hfffffff8; // @[TensorLoadWideVME.scala 524:51]
  reg [31:0] rdLineAddr; // @[TensorLoadWideVME.scala 538:23]
  wire [7:0] _rdLineAddr_T = {rdLen, 3'h0}; // @[TensorLoadWideVME.scala 545:41]
  wire [31:0] _GEN_35 = {{24'd0}, _rdLineAddr_T}; // @[TensorLoadWideVME.scala 545:32]
  wire [31:0] _rdLineAddr_T_2 = rdLineAddr + _GEN_35; // @[TensorLoadWideVME.scala 545:32]
  wire  _T_3 = ~reset; // @[TensorLoadWideVME.scala 563:9]
  wire [31:0] _GEN_36 = {{14'd0}, rdLineBytes}; // @[TensorLoadWideVME.scala 573:48]
  wire [31:0] _rdLastPulseBytes_T_1 = rdLineElemBeginAddr + _GEN_36; // @[TensorLoadWideVME.scala 573:48]
  wire [31:0] _GEN_3 = _rdLastPulseBytes_T_1 % 32'h8; // @[TensorLoadWideVME.scala 573:63]
  wire [3:0] rdLastPulseBytes = _GEN_3[3:0]; // @[TensorLoadWideVME.scala 573:63]
  wire [1:0] rdLastPulseTensNb = rdLastPulseBytes[3:2] == 2'h0 ? 2'h2 : rdLastPulseBytes[3:2]; // @[TensorLoadWideVME.scala 578:28]
  reg [6:0] rdCmdStartIdx; // @[TensorLoadWideVME.scala 588:26]
  reg  commandsDone; // @[TensorLoadWideVME.scala 589:29]
  wire [14:0] nextClIdx = clReadIdx + _GEN_33; // @[TensorLoadWideVME.scala 600:31]
  wire  _GEN_7 = nextClIdx == rdLineClNb & dramLineIdx == _T_31 | commandsDone; // @[TensorLoadWideVME.scala 595:16 602:71 603:20]
  wire  _GEN_9 = io_updateState ? _GEN_7 : commandsDone; // @[TensorLoadWideVME.scala 595:16 599:31]
  wire  _GEN_11 = io_start | stride ? 1'h0 : _GEN_9; // @[TensorLoadWideVME.scala 596:29 598:18]
  wire [1:0] rdCmd1stPluseOffsetTensNb = newReadRow ? rd1stPulseOffsetBytes[3:2] : 2'h0; // @[TensorLoadWideVME.scala 619:20 621:31 624:31]
  wire [1:0] rdCmdLastPluseTensNb = _T_29 ? rdLastPulseTensNb : 2'h2; // @[TensorLoadWideVME.scala 626:43 628:26 631:26]
  wire [15:0] _GEN_40 = {{12'd0}, io_xpad_0}; // @[TensorLoadWideVME.scala 657:29]
  wire [15:0] _totalWidth_T_1 = io_xsize + _GEN_40; // @[TensorLoadWideVME.scala 657:29]
  wire [15:0] _GEN_41 = {{12'd0}, io_xpad_1}; // @[TensorLoadWideVME.scala 657:41]
  wire [15:0] totalWidth = _totalWidth_T_1 + _GEN_41; // @[TensorLoadWideVME.scala 657:41]
  reg [19:0] currentRowIdx; // @[TensorLoadWideVME.scala 661:26]
  wire [19:0] _GEN_42 = {{16'd0}, io_ypad_0}; // @[TensorLoadWideVME.scala 663:39]
  wire [15:0] _GEN_43 = {{12'd0}, io_ypad_0}; // @[TensorLoadWideVME.scala 664:31]
  wire [15:0] _rdCmdStartIdxValid_T_2 = io_ysize + _GEN_43; // @[TensorLoadWideVME.scala 664:31]
  wire [19:0] _GEN_44 = {{4'd0}, _rdCmdStartIdxValid_T_2}; // @[TensorLoadWideVME.scala 664:19]
  wire  _rdCmdStartIdxValid_T_3 = currentRowIdx < _GEN_44; // @[TensorLoadWideVME.scala 664:19]
  wire  _rdCmdStartIdxValid_T_4 = currentRowIdx >= _GEN_42 & _rdCmdStartIdxValid_T_3; // @[TensorLoadWideVME.scala 663:52]
  wire  _rdCmdStartIdxValid_T_5 = _rdCmdStartIdxValid_T_4 & io_isBusy; // @[TensorLoadWideVME.scala 664:44]
  wire  _rdCmdStartIdxValid_T_6 = ~commandsDone; // @[TensorLoadWideVME.scala 666:5]
  wire  rdCmdStartIdxValid = _rdCmdStartIdxValid_T_5 & _rdCmdStartIdxValid_T_6; // @[TensorLoadWideVME.scala 665:15]
  wire [15:0] _rdCmdStartIdx_T_1 = io_sram_offset + _GEN_40; // @[TensorLoadWideVME.scala 669:37]
  wire [15:0] _GEN_47 = {{9'd0}, rdCmdStartIdx}; // @[TensorLoadWideVME.scala 671:36]
  wire [15:0] _rdCmdStartIdx_T_3 = _GEN_47 + totalWidth; // @[TensorLoadWideVME.scala 671:36]
  wire [19:0] _currentRowIdx_T_1 = currentRowIdx + 20'h1; // @[TensorLoadWideVME.scala 672:36]
  wire [15:0] _GEN_19 = io_isBusy & (currentRowIdx < _GEN_42 | stride) ? _rdCmdStartIdx_T_3 : {{9'd0}, rdCmdStartIdx}; // @[TensorLoadWideVME.scala 670:67 671:19 588:26]
  wire [15:0] _GEN_22 = io_start ? _rdCmdStartIdx_T_1 : _GEN_19; // @[TensorLoadWideVME.scala 667:19 669:19]
  wire  startIssueCmdRead = newReadRow & rdCmdStartIdxValid; // @[TensorLoadWideVME.scala 675:19]
  reg [6:0] rdCmdDestElemIdxNext; // @[TensorLoadWideVME.scala 688:33]
  wire [5:0] _rdCmdTransactionTensNb_T = {rdLen, 1'h0}; // @[TensorLoadWideVME.scala 694:39]
  wire [5:0] _GEN_48 = {{4'd0}, rdCmd1stPluseOffsetTensNb}; // @[TensorLoadWideVME.scala 694:71]
  wire [5:0] rdCmdTransactionTensNb = _rdCmdTransactionTensNb_T - _GEN_48; // @[TensorLoadWideVME.scala 694:71]
  wire [6:0] _GEN_49 = {{1'd0}, rdCmdTransactionTensNb}; // @[TensorLoadWideVME.scala 700:44]
  wire [6:0] _rdCmdDestElemIdxNext_T_1 = rdCmdStartIdx + _GEN_49; // @[TensorLoadWideVME.scala 700:44]
  wire [6:0] _rdCmdDestElemIdxNext_T_3 = rdCmdDestElemIdxNext + _GEN_49; // @[TensorLoadWideVME.scala 703:51]
  wire [6:0] _GEN_25 = startIssueCmdRead ? rdCmdStartIdx : rdCmdDestElemIdxNext; // @[TensorLoadWideVME.scala 690:20 698:29 699:24]
  wire [6:0] rdCmdDestElemIdx = rdCmdStartIdxValid ? _GEN_25 : rdCmdDestElemIdxNext; // @[TensorLoadWideVME.scala 690:20 696:28]
  wire [4:0] _io_vmeCmd_bits_len_T_1 = rdLen - 5'h1; // @[TensorLoadWideVME.scala 716:31]
  wire [31:0] _GEN_4 = rdLineAddr % 32'h80; // @[TensorLoadWideVME.scala 717:87]
  wire [7:0] _T_49 = _GEN_4[7:0]; // @[TensorLoadWideVME.scala 717:87]
  wire [7:0] _T_51 = 8'h80 - _T_49; // @[TensorLoadWideVME.scala 717:74]
  wire [10:0] _io_vmeCmd_bits_tag_T_1 = {rdCmdDestElemIdx,rdCmd1stPluseOffsetTensNb,rdCmdLastPluseTensNb}; // @[Cat.scala 31:58]
  assign io_vmeCmd_valid = _rdCmdStartIdxValid_T_5 & _rdCmdStartIdxValid_T_6; // @[TensorLoadWideVME.scala 665:15]
  assign io_vmeCmd_bits_addr = rdLineAddr; // @[TensorLoadWideVME.scala 715:23]
  assign io_vmeCmd_bits_len = _io_vmeCmd_bits_len_T_1[3:0]; // @[TensorLoadWideVME.scala 716:22]
  assign io_vmeCmd_bits_tag = {{10'd0}, _io_vmeCmd_bits_tag_T_1}; // @[TensorLoadWideVME.scala 721:22]
  assign io_readLen = _GEN_18[4:0]; // @[TensorLoadWideVME.scala 537:19]
  assign io_done = commandsDone; // @[TensorLoadWideVME.scala 726:11]
  always @(posedge clock) begin
    if (io_start) begin // @[TensorLoadWideVME.scala 502:19]
      dramLineIdx <= 16'h0; // @[TensorLoadWideVME.scala 503:17]
    end else if (stride) begin // @[TensorLoadWideVME.scala 504:23]
      dramLineIdx <= _dramLineIdx_T_1; // @[TensorLoadWideVME.scala 505:17]
    end
    if (io_start | stride) begin // @[TensorLoadWideVME.scala 596:29]
      clReadIdx <= 15'h0; // @[TensorLoadWideVME.scala 597:15]
    end else if (io_updateState) begin // @[TensorLoadWideVME.scala 599:31]
      clReadIdx <= nextClIdx; // @[TensorLoadWideVME.scala 601:15]
    end
    if (io_start) begin // @[TensorLoadWideVME.scala 525:19]
      rdLineElemBeginAddr <= xferElemInitAddr; // @[TensorLoadWideVME.scala 526:25]
    end else if (stride) begin // @[TensorLoadWideVME.scala 527:23]
      rdLineElemBeginAddr <= nextLineBeginElemAddr; // @[TensorLoadWideVME.scala 528:25]
    end
    if (io_start) begin // @[TensorLoadWideVME.scala 539:19]
      rdLineAddr <= xferClInitAddr; // @[TensorLoadWideVME.scala 540:16]
    end else if (io_updateState) begin // @[TensorLoadWideVME.scala 541:31]
      if (stride) begin // @[TensorLoadWideVME.scala 542:18]
        rdLineAddr <= nextLineBeginClAddr; // @[TensorLoadWideVME.scala 543:18]
      end else begin
        rdLineAddr <= _rdLineAddr_T_2; // @[TensorLoadWideVME.scala 545:18]
      end
    end
    rdCmdStartIdx <= _GEN_22[6:0];
    commandsDone <= reset | _GEN_11; // @[TensorLoadWideVME.scala 589:{29,29}]
    if (io_start) begin // @[TensorLoadWideVME.scala 667:19]
      currentRowIdx <= 20'h0; // @[TensorLoadWideVME.scala 668:19]
    end else if (io_isBusy & (currentRowIdx < _GEN_42 | stride)) begin // @[TensorLoadWideVME.scala 670:67]
      currentRowIdx <= _currentRowIdx_T_1; // @[TensorLoadWideVME.scala 672:19]
    end
    if (rdCmdStartIdxValid) begin // @[TensorLoadWideVME.scala 696:28]
      if (startIssueCmdRead) begin // @[TensorLoadWideVME.scala 698:29]
        rdCmdDestElemIdxNext <= _rdCmdDestElemIdxNext_T_1; // @[TensorLoadWideVME.scala 700:27]
      end else if (io_updateState) begin // @[TensorLoadWideVME.scala 701:33]
        rdCmdDestElemIdxNext <= _rdCmdDestElemIdxNext_T_3; // @[TensorLoadWideVME.scala 703:27]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(rd1stPulseOffsetBytes[3:2] <= 2'h2)) begin
          $fwrite(32'h80000002,
            "Assertion failed: -F- Expecting the number of tensors to skip in CL\n    at TensorLoadWideVME.scala:563 assert(rd1stPulseOffsetBytes >> log2Ceil(elemBytes) <= tp.clSizeRatio.U,\n"
            ); // @[TensorLoadWideVME.scala 563:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~(rdLastPulseBytes[3:2] <= 2'h2)) begin
          $fwrite(32'h80000002,
            "Assertion failed: -F- Expecting the number of active tensors in CL\n    at TensorLoadWideVME.scala:574 assert(rdLastPulseBytes >> log2Ceil(elemBytes) <= (clBytes/elemBytes).U,\n"
            ); // @[TensorLoadWideVME.scala 574:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~(~io_isBusy | rdLineClNb >= clReadIdx)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorLoadWideVME.scala:641 assert(!io.isBusy || rdLineClNb >= clReadIdx)// define how many cachelines to read at this cycle\n"
            ); // @[TensorLoadWideVME.scala 641:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~(~io_vmeCmd_valid | _rdLineAddr_T <= _T_51)) begin
          $fwrite(32'h80000002,
            "Assertion failed: -F- uop DRAM page alignment failure. DRAM address + len overlaps mp.lenBits*memBlockSize alignment %x %x\n    at TensorLoadWideVME.scala:717 assert(!io.vmeCmd.valid || ((rdLen << log2Ceil(clBytes)) <= maxTrBytes - rdLineAddr %% maxTrBytes),\n"
            ,rdLineAddr,rdLen); // @[TensorLoadWideVME.scala 717:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dramLineIdx = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  clReadIdx = _RAND_1[14:0];
  _RAND_2 = {1{`RANDOM}};
  rdLineElemBeginAddr = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  rdLineAddr = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  rdCmdStartIdx = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  commandsDone = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  currentRowIdx = _RAND_6[19:0];
  _RAND_7 = {1{`RANDOM}};
  rdCmdDestElemIdxNext = _RAND_7[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(rd1stPulseOffsetBytes[3:2] <= 2'h2); // @[TensorLoadWideVME.scala 563:9]
    end
    //
    if (_T_3) begin
      assert(rdLastPulseBytes[3:2] <= 2'h2); // @[TensorLoadWideVME.scala 574:9]
    end
    //
    if (_T_3) begin
      assert(~io_isBusy | rdLineClNb >= clReadIdx); // @[TensorLoadWideVME.scala 641:9]
    end
    //
    if (_T_3) begin
      assert(~io_vmeCmd_valid | _rdLineAddr_T <= _T_51); // @[TensorLoadWideVME.scala 717:9]
    end
  end
endmodule
module GenVMECmdWideTL(
  input          clock,
  input          reset,
  input          io_start,
  input          io_isBusy,
  input  [127:0] io_inst,
  input  [31:0]  io_baddr,
  input          io_vmeCmd_ready,
  output         io_vmeCmd_valid,
  output [31:0]  io_vmeCmd_bits_addr,
  output [3:0]   io_vmeCmd_bits_len,
  output [20:0]  io_vmeCmd_bits_tag,
  output [4:0]   io_readLen,
  output         io_done
);
  wire  cmdGen_clock; // @[TensorLoadWideVME.scala 746:23]
  wire  cmdGen_reset; // @[TensorLoadWideVME.scala 746:23]
  wire  cmdGen_io_start; // @[TensorLoadWideVME.scala 746:23]
  wire  cmdGen_io_isBusy; // @[TensorLoadWideVME.scala 746:23]
  wire  cmdGen_io_updateState; // @[TensorLoadWideVME.scala 746:23]
  wire [31:0] cmdGen_io_baddr; // @[TensorLoadWideVME.scala 746:23]
  wire  cmdGen_io_vmeCmd_valid; // @[TensorLoadWideVME.scala 746:23]
  wire [31:0] cmdGen_io_vmeCmd_bits_addr; // @[TensorLoadWideVME.scala 746:23]
  wire [3:0] cmdGen_io_vmeCmd_bits_len; // @[TensorLoadWideVME.scala 746:23]
  wire [20:0] cmdGen_io_vmeCmd_bits_tag; // @[TensorLoadWideVME.scala 746:23]
  wire [4:0] cmdGen_io_readLen; // @[TensorLoadWideVME.scala 746:23]
  wire  cmdGen_io_done; // @[TensorLoadWideVME.scala 746:23]
  wire [15:0] cmdGen_io_ysize; // @[TensorLoadWideVME.scala 746:23]
  wire [15:0] cmdGen_io_xsize; // @[TensorLoadWideVME.scala 746:23]
  wire [15:0] cmdGen_io_xstride; // @[TensorLoadWideVME.scala 746:23]
  wire [31:0] cmdGen_io_dram_offset; // @[TensorLoadWideVME.scala 746:23]
  wire [15:0] cmdGen_io_sram_offset; // @[TensorLoadWideVME.scala 746:23]
  wire [3:0] cmdGen_io_xpad_0; // @[TensorLoadWideVME.scala 746:23]
  wire [3:0] cmdGen_io_xpad_1; // @[TensorLoadWideVME.scala 746:23]
  wire [3:0] cmdGen_io_ypad_0; // @[TensorLoadWideVME.scala 746:23]
  GenVMECmdWide cmdGen ( // @[TensorLoadWideVME.scala 746:23]
    .clock(cmdGen_clock),
    .reset(cmdGen_reset),
    .io_start(cmdGen_io_start),
    .io_isBusy(cmdGen_io_isBusy),
    .io_updateState(cmdGen_io_updateState),
    .io_baddr(cmdGen_io_baddr),
    .io_vmeCmd_valid(cmdGen_io_vmeCmd_valid),
    .io_vmeCmd_bits_addr(cmdGen_io_vmeCmd_bits_addr),
    .io_vmeCmd_bits_len(cmdGen_io_vmeCmd_bits_len),
    .io_vmeCmd_bits_tag(cmdGen_io_vmeCmd_bits_tag),
    .io_readLen(cmdGen_io_readLen),
    .io_done(cmdGen_io_done),
    .io_ysize(cmdGen_io_ysize),
    .io_xsize(cmdGen_io_xsize),
    .io_xstride(cmdGen_io_xstride),
    .io_dram_offset(cmdGen_io_dram_offset),
    .io_sram_offset(cmdGen_io_sram_offset),
    .io_xpad_0(cmdGen_io_xpad_0),
    .io_xpad_1(cmdGen_io_xpad_1),
    .io_ypad_0(cmdGen_io_ypad_0)
  );
  assign io_vmeCmd_valid = cmdGen_io_vmeCmd_valid; // @[TensorLoadWideVME.scala 751:13]
  assign io_vmeCmd_bits_addr = cmdGen_io_vmeCmd_bits_addr; // @[TensorLoadWideVME.scala 751:13]
  assign io_vmeCmd_bits_len = cmdGen_io_vmeCmd_bits_len; // @[TensorLoadWideVME.scala 751:13]
  assign io_vmeCmd_bits_tag = cmdGen_io_vmeCmd_bits_tag; // @[TensorLoadWideVME.scala 751:13]
  assign io_readLen = cmdGen_io_readLen; // @[TensorLoadWideVME.scala 752:14]
  assign io_done = cmdGen_io_done; // @[TensorLoadWideVME.scala 753:11]
  assign cmdGen_clock = clock;
  assign cmdGen_reset = reset;
  assign cmdGen_io_start = io_start; // @[TensorLoadWideVME.scala 748:19]
  assign cmdGen_io_isBusy = io_isBusy; // @[TensorLoadWideVME.scala 749:20]
  assign cmdGen_io_updateState = io_vmeCmd_ready & io_vmeCmd_valid; // @[Decoupled.scala 50:35]
  assign cmdGen_io_baddr = io_baddr; // @[TensorLoadWideVME.scala 750:19]
  assign cmdGen_io_ysize = io_inst[79:64]; // @[TensorLoadWideVME.scala 744:29]
  assign cmdGen_io_xsize = io_inst[95:80]; // @[TensorLoadWideVME.scala 744:29]
  assign cmdGen_io_xstride = io_inst[111:96]; // @[TensorLoadWideVME.scala 744:29]
  assign cmdGen_io_dram_offset = io_inst[57:26]; // @[TensorLoadWideVME.scala 744:29]
  assign cmdGen_io_sram_offset = io_inst[25:10]; // @[TensorLoadWideVME.scala 744:29]
  assign cmdGen_io_xpad_0 = io_inst[123:120]; // @[TensorLoadWideVME.scala 744:29]
  assign cmdGen_io_xpad_1 = io_inst[127:124]; // @[TensorLoadWideVME.scala 744:29]
  assign cmdGen_io_ypad_0 = io_inst[115:112]; // @[TensorLoadWideVME.scala 744:29]
endmodule
module ReadVMEDataWide(
  input         clock,
  input         reset,
  input         io_start,
  output        io_vmeData_ready,
  input         io_vmeData_valid,
  input  [63:0] io_vmeData_bits_data,
  input  [20:0] io_vmeData_bits_tag,
  input         io_vmeData_bits_last,
  output [6:0]  io_destIdx_0,
  output [6:0]  io_destIdx_1,
  output [31:0] io_destData_0,
  output [31:0] io_destData_1,
  output        io_destMask_0,
  output        io_destMask_1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [20:0] vmeTagDecodeLast; // @[TensorLoadWideVME.scala 352:29]
  wire [16:0] rdDataElemIdx = io_vmeData_bits_tag[20:4]; // @[TensorLoadWideVME.scala 356:35]
  wire [1:0] rdFstOffsetNb = io_vmeData_bits_tag[3:2]; // @[TensorLoadWideVME.scala 360:35]
  wire [1:0] rdLstNb = io_vmeData_bits_tag[1:0]; // @[TensorLoadWideVME.scala 366:31]
  wire [1:0] _wrMask1st_T_1 = 2'h2 - rdFstOffsetNb; // @[TensorLoadWideVME.scala 374:32]
  wire  _wrMask1st_T_2 = 2'h0 < _wrMask1st_T_1; // @[TensorLoadWideVME.scala 374:13]
  wire  _wrMask1st_T_5 = 2'h1 < _wrMask1st_T_1; // @[TensorLoadWideVME.scala 374:13]
  wire [1:0] _wrMask1st_T_6 = {_wrMask1st_T_5,_wrMask1st_T_2}; // @[TensorLoadWideVME.scala 375:8]
  wire [1:0] wrMask1st = {_wrMask1st_T_6[0],_wrMask1st_T_6[1]}; // @[Cat.scala 31:58]
  wire  _wrMaskLast_T = 2'h0 < rdLstNb; // @[TensorLoadWideVME.scala 381:13]
  wire  _wrMaskLast_T_1 = 2'h1 < rdLstNb; // @[TensorLoadWideVME.scala 381:13]
  wire [1:0] wrMaskLast = {_wrMaskLast_T_1,_wrMaskLast_T}; // @[TensorLoadWideVME.scala 382:8]
  reg [6:0] rdDataElemDestIdxNext; // @[TensorLoadWideVME.scala 385:34]
  wire  _T_1 = io_vmeData_ready & io_vmeData_valid; // @[Decoupled.scala 50:35]
  reg  vmeTagDecodeLastValidNext; // @[TensorLoadWideVME.scala 390:42]
  wire  _T_3 = io_vmeData_bits_tag != vmeTagDecodeLast; // @[TensorLoadWideVME.scala 421:29]
  wire  _T_4 = vmeTagDecodeLastValidNext & _T_3; // @[TensorLoadWideVME.scala 420:34]
  wire  _T_5 = ~vmeTagDecodeLastValidNext | _T_4; // @[TensorLoadWideVME.scala 419:34]
  wire [16:0] _GEN_4 = _T_5 ? rdDataElemIdx : {{10'd0}, rdDataElemDestIdxNext}; // @[TensorLoadWideVME.scala 421:59 425:25 430:25]
  wire [6:0] rdDataElemDestIdx = _GEN_4[6:0]; // @[TensorLoadWideVME.scala 384:31]
  wire [5:0] rdDataClDestIdx = rdDataElemDestIdx[6:1]; // @[TensorLoadWideVME.scala 386:43]
  wire [6:0] _GEN_1 = rdDataElemDestIdx % 7'h2; // @[TensorLoadWideVME.scala 387:48]
  wire [1:0] rdDataDestElemOffset = _GEN_1[1:0]; // @[TensorLoadWideVME.scala 387:48]
  wire  _GEN_0 = _T_1 | vmeTagDecodeLastValidNext; // @[TensorLoadWideVME.scala 395:31 396:27 398:27]
  wire  isFirstPulse = _T_1 & _T_5; // @[TensorLoadWideVME.scala 416:16 417:25]
  wire  _wmaskSel_T = isFirstPulse & io_vmeData_bits_last; // @[TensorLoadWideVME.scala 405:20]
  wire [1:0] _wmaskSel_T_1 = wrMask1st & wrMaskLast; // @[TensorLoadWideVME.scala 406:17]
  wire [1:0] _wmaskSel_T_2 = io_vmeData_bits_last ? wrMaskLast : 2'h3; // @[TensorLoadWideVME.scala 410:12]
  wire [1:0] _wmaskSel_T_3 = isFirstPulse ? wrMask1st : _wmaskSel_T_2; // @[TensorLoadWideVME.scala 407:10]
  wire [1:0] wmaskSel = _wmaskSel_T ? _wmaskSel_T_1 : _wmaskSel_T_3; // @[TensorLoadWideVME.scala 404:8]
  wire [1:0] wmask = _T_1 ? wmaskSel : 2'h0; // @[TensorLoadWideVME.scala 414:18]
  wire [1:0] _rdDataElemDestIdxNext_T_2 = wmask[0] + wmask[1]; // @[Bitwise.scala 48:55]
  wire [16:0] _GEN_10 = {{15'd0}, _rdDataElemDestIdxNext_T_2}; // @[TensorLoadWideVME.scala 427:46]
  wire [16:0] _rdDataElemDestIdxNext_T_5 = rdDataElemIdx + _GEN_10; // @[TensorLoadWideVME.scala 427:46]
  wire [6:0] _GEN_11 = {{5'd0}, _rdDataElemDestIdxNext_T_2}; // @[TensorLoadWideVME.scala 429:54]
  wire [6:0] _rdDataElemDestIdxNext_T_11 = rdDataElemDestIdxNext + _GEN_11; // @[TensorLoadWideVME.scala 429:54]
  wire [16:0] _GEN_5 = _T_5 ? _rdDataElemDestIdxNext_T_5 : {{10'd0}, _rdDataElemDestIdxNext_T_11}; // @[TensorLoadWideVME.scala 421:59 427:29 429:29]
  wire [16:0] _GEN_9 = _T_1 ? _GEN_5 : {{10'd0}, rdDataElemDestIdxNext}; // @[TensorLoadWideVME.scala 417:25 385:34]
  wire [31:0] srcData_0 = io_vmeData_bits_data[31:0]; // @[TensorLoadWideVME.scala 435:47]
  wire [31:0] srcData_1 = io_vmeData_bits_data[63:32]; // @[TensorLoadWideVME.scala 435:47]
  wire [1:0] _srcOffset_0_T = isFirstPulse ? rdFstOffsetNb : 2'h0; // @[TensorLoadWideVME.scala 441:30]
  wire [2:0] _srcOffset_0_T_1 = {{1'd0}, _srcOffset_0_T}; // @[TensorLoadWideVME.scala 441:25]
  wire [1:0] srcOffset_0 = _srcOffset_0_T_1[1:0]; // @[TensorLoadWideVME.scala 441:25]
  wire [1:0] _srcIdx_0_T_1 = srcOffset_0 - rdDataDestElemOffset; // @[TensorLoadWideVME.scala 442:31]
  wire  srcIdx_0 = _srcIdx_0_T_1[0]; // @[TensorLoadWideVME.scala 437:20 442:15]
  wire [1:0] srcIdxOH = 2'h1 << srcIdx_0; // @[OneHot.scala 57:35]
  wire [31:0] _io_destData_0_T_2 = srcIdxOH[0] ? srcData_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_destData_0_T_3 = srcIdxOH[1] ? srcData_1 : 32'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_destMask_0_T = srcIdxOH & wmask; // @[Mux.scala 30:47]
  wire  incrIdx = srcOffset_0 >= rdDataDestElemOffset ? 1'h0 : 1'h1; // @[TensorLoadWideVME.scala 451:10]
  wire [5:0] _GEN_12 = {{5'd0}, incrIdx}; // @[TensorLoadWideVME.scala 453:38]
  wire [5:0] _io_destIdx_0_T_1 = rdDataClDestIdx + _GEN_12; // @[TensorLoadWideVME.scala 453:38]
  wire [1:0] srcOffset_1 = 2'h1 + _srcOffset_0_T; // @[TensorLoadWideVME.scala 441:25]
  wire [1:0] _srcIdx_1_T_1 = srcOffset_1 - rdDataDestElemOffset; // @[TensorLoadWideVME.scala 442:31]
  wire  srcIdx_1 = _srcIdx_1_T_1[0]; // @[TensorLoadWideVME.scala 437:20 442:15]
  wire [1:0] srcIdxOH_1 = 2'h1 << srcIdx_1; // @[OneHot.scala 57:35]
  wire [31:0] _io_destData_1_T_2 = srcIdxOH_1[0] ? srcData_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _io_destData_1_T_3 = srcIdxOH_1[1] ? srcData_1 : 32'h0; // @[Mux.scala 27:73]
  wire [1:0] _io_destMask_1_T = srcIdxOH_1 & wmask; // @[Mux.scala 30:47]
  wire  incrIdx_1 = srcOffset_1 >= rdDataDestElemOffset ? 1'h0 : 1'h1; // @[TensorLoadWideVME.scala 451:10]
  wire [5:0] _GEN_13 = {{5'd0}, incrIdx_1}; // @[TensorLoadWideVME.scala 453:38]
  wire [5:0] _io_destIdx_1_T_1 = rdDataClDestIdx + _GEN_13; // @[TensorLoadWideVME.scala 453:38]
  assign io_vmeData_ready = 1'h1; // @[TensorLoadWideVME.scala 344:20]
  assign io_destIdx_0 = {{1'd0}, _io_destIdx_0_T_1}; // @[TensorLoadWideVME.scala 453:19]
  assign io_destIdx_1 = {{1'd0}, _io_destIdx_1_T_1}; // @[TensorLoadWideVME.scala 453:19]
  assign io_destData_0 = _io_destData_0_T_2 | _io_destData_0_T_3; // @[Mux.scala 27:73]
  assign io_destData_1 = _io_destData_1_T_2 | _io_destData_1_T_3; // @[Mux.scala 27:73]
  assign io_destMask_0 = |_io_destMask_0_T; // @[Mux.scala 30:53]
  assign io_destMask_1 = |_io_destMask_1_T; // @[Mux.scala 30:53]
  always @(posedge clock) begin
    if (_T_1) begin // @[TensorLoadWideVME.scala 417:25]
      if (_T_5) begin // @[TensorLoadWideVME.scala 421:59]
        vmeTagDecodeLast <= io_vmeData_bits_tag; // @[TensorLoadWideVME.scala 423:24]
      end
    end
    rdDataElemDestIdxNext <= _GEN_9[6:0];
    if (reset) begin // @[TensorLoadWideVME.scala 390:42]
      vmeTagDecodeLastValidNext <= 1'h0; // @[TensorLoadWideVME.scala 390:42]
    end else if (io_start) begin // @[TensorLoadWideVME.scala 393:18]
      vmeTagDecodeLastValidNext <= 1'h0; // @[TensorLoadWideVME.scala 394:27]
    end else begin
      vmeTagDecodeLastValidNext <= _GEN_0;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~io_vmeData_valid | rdLstNb > 2'h0)) begin
          $fwrite(32'h80000002,
            "Assertion failed: -F- Expecting some elements to read\n    at TensorLoadWideVME.scala:367 assert(!io.vmeData.valid || readNb > 0.U,\"-F- Expecting some elements to read\")\n"
            ); // @[TensorLoadWideVME.scala 367:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  vmeTagDecodeLast = _RAND_0[20:0];
  _RAND_1 = {1{`RANDOM}};
  rdDataElemDestIdxNext = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  vmeTagDecodeLastValidNext = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~io_vmeData_valid | rdLstNb > 2'h0); // @[TensorLoadWideVME.scala 367:11]
    end
  end
endmodule
module TensorLoadWideVME(
  input          clock,
  input          reset,
  input          io_start,
  output         io_done,
  input  [127:0] io_inst,
  input  [31:0]  io_baddr,
  input          io_vme_rd_cmd_ready,
  output         io_vme_rd_cmd_valid,
  output [31:0]  io_vme_rd_cmd_bits_addr,
  output [3:0]   io_vme_rd_cmd_bits_len,
  output [20:0]  io_vme_rd_cmd_bits_tag,
  output         io_vme_rd_data_ready,
  input          io_vme_rd_data_valid,
  input  [63:0]  io_vme_rd_data_bits_data,
  input  [20:0]  io_vme_rd_data_bits_tag,
  input          io_vme_rd_data_bits_last,
  input          io_tensor_rd_0_idx_valid,
  input  [6:0]   io_tensor_rd_0_idx_bits,
  output         io_tensor_rd_0_data_valid,
  output [31:0]  io_tensor_rd_0_data_bits_0_0
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  vmeCmd_clock; // @[TensorLoadWideVME.scala 105:23]
  wire  vmeCmd_reset; // @[TensorLoadWideVME.scala 105:23]
  wire  vmeCmd_io_start; // @[TensorLoadWideVME.scala 105:23]
  wire  vmeCmd_io_isBusy; // @[TensorLoadWideVME.scala 105:23]
  wire [127:0] vmeCmd_io_inst; // @[TensorLoadWideVME.scala 105:23]
  wire [31:0] vmeCmd_io_baddr; // @[TensorLoadWideVME.scala 105:23]
  wire  vmeCmd_io_vmeCmd_ready; // @[TensorLoadWideVME.scala 105:23]
  wire  vmeCmd_io_vmeCmd_valid; // @[TensorLoadWideVME.scala 105:23]
  wire [31:0] vmeCmd_io_vmeCmd_bits_addr; // @[TensorLoadWideVME.scala 105:23]
  wire [3:0] vmeCmd_io_vmeCmd_bits_len; // @[TensorLoadWideVME.scala 105:23]
  wire [20:0] vmeCmd_io_vmeCmd_bits_tag; // @[TensorLoadWideVME.scala 105:23]
  wire [4:0] vmeCmd_io_readLen; // @[TensorLoadWideVME.scala 105:23]
  wire  vmeCmd_io_done; // @[TensorLoadWideVME.scala 105:23]
  wire  readData_clock; // @[TensorLoadWideVME.scala 150:24]
  wire  readData_reset; // @[TensorLoadWideVME.scala 150:24]
  wire  readData_io_start; // @[TensorLoadWideVME.scala 150:24]
  wire  readData_io_vmeData_ready; // @[TensorLoadWideVME.scala 150:24]
  wire  readData_io_vmeData_valid; // @[TensorLoadWideVME.scala 150:24]
  wire [63:0] readData_io_vmeData_bits_data; // @[TensorLoadWideVME.scala 150:24]
  wire [20:0] readData_io_vmeData_bits_tag; // @[TensorLoadWideVME.scala 150:24]
  wire  readData_io_vmeData_bits_last; // @[TensorLoadWideVME.scala 150:24]
  wire [6:0] readData_io_destIdx_0; // @[TensorLoadWideVME.scala 150:24]
  wire [6:0] readData_io_destIdx_1; // @[TensorLoadWideVME.scala 150:24]
  wire [31:0] readData_io_destData_0; // @[TensorLoadWideVME.scala 150:24]
  wire [31:0] readData_io_destData_1; // @[TensorLoadWideVME.scala 150:24]
  wire  readData_io_destMask_0; // @[TensorLoadWideVME.scala 150:24]
  wire  readData_io_destMask_1; // @[TensorLoadWideVME.scala 150:24]
  wire  fillPadding_clock; // @[TensorLoadWideVME.scala 166:27]
  wire  fillPadding_reset; // @[TensorLoadWideVME.scala 166:27]
  wire  fillPadding_io_canWriteMem; // @[TensorLoadWideVME.scala 166:27]
  wire [127:0] fillPadding_io_inst; // @[TensorLoadWideVME.scala 166:27]
  wire  fillPadding_io_tensorIdx_valid; // @[TensorLoadWideVME.scala 166:27]
  wire [6:0] fillPadding_io_tensorIdx_bits; // @[TensorLoadWideVME.scala 166:27]
  wire  fillPadding_io_start; // @[TensorLoadWideVME.scala 166:27]
  wire  fillPadding_io_done; // @[TensorLoadWideVME.scala 166:27]
  reg [31:0] tensorFile_0 [0:63]; // @[TensorLoadWideVME.scala 193:16]
  wire  tensorFile_0_rdataVec_MPORT_en; // @[TensorLoadWideVME.scala 193:16]
  wire [5:0] tensorFile_0_rdataVec_MPORT_addr; // @[TensorLoadWideVME.scala 193:16]
  wire [31:0] tensorFile_0_rdataVec_MPORT_data; // @[TensorLoadWideVME.scala 193:16]
  wire [31:0] tensorFile_0_MPORT_data; // @[TensorLoadWideVME.scala 193:16]
  wire [5:0] tensorFile_0_MPORT_addr; // @[TensorLoadWideVME.scala 193:16]
  wire  tensorFile_0_MPORT_mask; // @[TensorLoadWideVME.scala 193:16]
  wire  tensorFile_0_MPORT_en; // @[TensorLoadWideVME.scala 193:16]
  reg  tensorFile_0_rdataVec_MPORT_en_pipe_0;
  reg [5:0] tensorFile_0_rdataVec_MPORT_addr_pipe_0;
  reg [31:0] tensorFile_1 [0:63]; // @[TensorLoadWideVME.scala 193:16]
  wire  tensorFile_1_rdataVec_MPORT_1_en; // @[TensorLoadWideVME.scala 193:16]
  wire [5:0] tensorFile_1_rdataVec_MPORT_1_addr; // @[TensorLoadWideVME.scala 193:16]
  wire [31:0] tensorFile_1_rdataVec_MPORT_1_data; // @[TensorLoadWideVME.scala 193:16]
  wire [31:0] tensorFile_1_MPORT_1_data; // @[TensorLoadWideVME.scala 193:16]
  wire [5:0] tensorFile_1_MPORT_1_addr; // @[TensorLoadWideVME.scala 193:16]
  wire  tensorFile_1_MPORT_1_mask; // @[TensorLoadWideVME.scala 193:16]
  wire  tensorFile_1_MPORT_1_en; // @[TensorLoadWideVME.scala 193:16]
  reg  tensorFile_1_rdataVec_MPORT_1_en_pipe_0;
  reg [5:0] tensorFile_1_rdataVec_MPORT_1_addr_pipe_0;
  reg  state; // @[TensorLoadWideVME.scala 84:22]
  reg [6:0] clInFlight; // @[TensorLoadWideVME.scala 132:23]
  wire  loadDone = clInFlight == 7'h0 & vmeCmd_io_done & state; // @[TensorLoadWideVME.scala 315:53]
  wire  localDone = loadDone & fillPadding_io_done; // @[TensorLoadWideVME.scala 316:25]
  wire  _GEN_0 = localDone ? 1'h0 : state; // @[TensorLoadWideVME.scala 90:25 91:11 84:22]
  wire  _GEN_1 = io_start | _GEN_0; // @[TensorLoadWideVME.scala 88:18 89:11]
  wire  vmeDataFirePipe = io_vme_rd_data_valid & io_vme_rd_data_ready; // @[TensorLoadWideVME.scala 100:42]
  wire  _T = io_vme_rd_cmd_ready & io_vme_rd_cmd_valid; // @[Decoupled.scala 50:35]
  wire  _T_1 = state & _T; // @[TensorLoadWideVME.scala 135:21]
  wire  _T_3 = state & _T & ~vmeDataFirePipe; // @[TensorLoadWideVME.scala 135:43]
  wire [6:0] _GEN_26 = {{2'd0}, vmeCmd_io_readLen}; // @[TensorLoadWideVME.scala 136:30]
  wire [6:0] _clInFlight_T_1 = clInFlight + _GEN_26; // @[TensorLoadWideVME.scala 136:30]
  wire  _T_6 = _T_1 & vmeDataFirePipe; // @[TensorLoadWideVME.scala 137:43]
  wire [6:0] _clInFlight_T_5 = _clInFlight_T_1 - 7'h1; // @[TensorLoadWideVME.scala 138:40]
  wire  _T_10 = state & ~_T & vmeDataFirePipe; // @[TensorLoadWideVME.scala 139:44]
  wire  _T_13 = ~reset; // @[TensorLoadWideVME.scala 140:11]
  wire [6:0] _clInFlight_T_7 = clInFlight - 7'h1; // @[TensorLoadWideVME.scala 141:30]
  wire [5:0] zpDestIdx = fillPadding_io_tensorIdx_bits[6:1]; // @[TensorLoadWideVME.scala 172:49]
  wire [1:0] zpDestMask = 2'h1 << fillPadding_io_tensorIdx_bits[0]; // @[OneHot.scala 57:35]
  wire  _wmask_0_T = ~state; // @[TensorLoadWideVME.scala 223:33]
  wire  _wmask_0_T_3 = vmeDataFirePipe & readData_io_destMask_0; // @[TensorLoadWideVME.scala 228:18]
  wire  _wmask_0_T_4 = fillPadding_io_tensorIdx_valid ? zpDestMask[0] : _wmask_0_T_3; // @[TensorLoadWideVME.scala 225:16]
  wire  _wmask_1_T_3 = vmeDataFirePipe & readData_io_destMask_1; // @[TensorLoadWideVME.scala 228:18]
  wire  _wmask_1_T_4 = fillPadding_io_tensorIdx_valid ? zpDestMask[1] : _wmask_1_T_3; // @[TensorLoadWideVME.scala 225:16]
  wire [31:0] _wdata_0_WIRE_2 = readData_io_destData_0;
  wire [31:0] _wdata_0_T_2 = fillPadding_io_tensorIdx_valid ? 32'h0 : _wdata_0_WIRE_2; // @[TensorLoadWideVME.scala 243:12]
  wire [31:0] _wdata_1_WIRE_2 = readData_io_destData_1;
  wire [31:0] _wdata_1_T_2 = fillPadding_io_tensorIdx_valid ? 32'h0 : _wdata_1_WIRE_2; // @[TensorLoadWideVME.scala 243:12]
  wire [6:0] _widx_0_T_1 = fillPadding_io_tensorIdx_valid ? {{1'd0}, zpDestIdx} : readData_io_destIdx_0; // @[TensorLoadWideVME.scala 259:16]
  wire [6:0] widx_0 = _wmask_0_T ? 7'h0 : _widx_0_T_1; // @[TensorLoadWideVME.scala 256:14]
  wire [6:0] _widx_1_T_1 = fillPadding_io_tensorIdx_valid ? {{1'd0}, zpDestIdx} : readData_io_destIdx_1; // @[TensorLoadWideVME.scala 259:16]
  wire [6:0] widx_1 = _wmask_0_T ? 7'h0 : _widx_1_T_1; // @[TensorLoadWideVME.scala 256:14]
  wire [1:0] _rMask_T_1 = 2'h1 << io_tensor_rd_0_idx_bits[0]; // @[OneHot.scala 57:35]
  wire [1:0] rMask = io_tensor_rd_0_idx_valid ? _rMask_T_1 : 2'h0; // @[TensorLoadWideVME.scala 290:10]
  reg [1:0] rdata_r; // @[Reg.scala 16:16]
  wire [31:0] _rdataVec_WIRE_2_0 = tensorFile_0_rdataVec_MPORT_data; // @[TensorLoadWideVME.scala 297:{14,14}]
  wire [31:0] _rdata_T_2 = rdata_r[0] ? _rdataVec_WIRE_2_0 : 32'h0; // @[Mux.scala 27:73]
  wire [31:0] _rdataVec_WIRE_5_0 = tensorFile_1_rdataVec_MPORT_1_data; // @[TensorLoadWideVME.scala 297:{14,14}]
  wire [31:0] _rdata_T_3 = rdata_r[1] ? _rdataVec_WIRE_5_0 : 32'h0; // @[Mux.scala 27:73]
  reg  rvalid; // @[Reg.scala 28:20]
  GenVMECmdWideTL vmeCmd ( // @[TensorLoadWideVME.scala 105:23]
    .clock(vmeCmd_clock),
    .reset(vmeCmd_reset),
    .io_start(vmeCmd_io_start),
    .io_isBusy(vmeCmd_io_isBusy),
    .io_inst(vmeCmd_io_inst),
    .io_baddr(vmeCmd_io_baddr),
    .io_vmeCmd_ready(vmeCmd_io_vmeCmd_ready),
    .io_vmeCmd_valid(vmeCmd_io_vmeCmd_valid),
    .io_vmeCmd_bits_addr(vmeCmd_io_vmeCmd_bits_addr),
    .io_vmeCmd_bits_len(vmeCmd_io_vmeCmd_bits_len),
    .io_vmeCmd_bits_tag(vmeCmd_io_vmeCmd_bits_tag),
    .io_readLen(vmeCmd_io_readLen),
    .io_done(vmeCmd_io_done)
  );
  ReadVMEDataWide readData ( // @[TensorLoadWideVME.scala 150:24]
    .clock(readData_clock),
    .reset(readData_reset),
    .io_start(readData_io_start),
    .io_vmeData_ready(readData_io_vmeData_ready),
    .io_vmeData_valid(readData_io_vmeData_valid),
    .io_vmeData_bits_data(readData_io_vmeData_bits_data),
    .io_vmeData_bits_tag(readData_io_vmeData_bits_tag),
    .io_vmeData_bits_last(readData_io_vmeData_bits_last),
    .io_destIdx_0(readData_io_destIdx_0),
    .io_destIdx_1(readData_io_destIdx_1),
    .io_destData_0(readData_io_destData_0),
    .io_destData_1(readData_io_destData_1),
    .io_destMask_0(readData_io_destMask_0),
    .io_destMask_1(readData_io_destMask_1)
  );
  ZeroPadding fillPadding ( // @[TensorLoadWideVME.scala 166:27]
    .clock(fillPadding_clock),
    .reset(fillPadding_reset),
    .io_canWriteMem(fillPadding_io_canWriteMem),
    .io_inst(fillPadding_io_inst),
    .io_tensorIdx_valid(fillPadding_io_tensorIdx_valid),
    .io_tensorIdx_bits(fillPadding_io_tensorIdx_bits),
    .io_start(fillPadding_io_start),
    .io_done(fillPadding_io_done)
  );
  assign tensorFile_0_rdataVec_MPORT_en = tensorFile_0_rdataVec_MPORT_en_pipe_0;
  assign tensorFile_0_rdataVec_MPORT_addr = tensorFile_0_rdataVec_MPORT_addr_pipe_0;
  assign tensorFile_0_rdataVec_MPORT_data = tensorFile_0[tensorFile_0_rdataVec_MPORT_addr]; // @[TensorLoadWideVME.scala 193:16]
  assign tensorFile_0_MPORT_data = _wmask_0_T ? 32'h0 : _wdata_0_T_2;
  assign tensorFile_0_MPORT_addr = widx_0[5:0];
  assign tensorFile_0_MPORT_mask = 1'h1;
  assign tensorFile_0_MPORT_en = _wmask_0_T ? 1'h0 : _wmask_0_T_4;
  assign tensorFile_1_rdataVec_MPORT_1_en = tensorFile_1_rdataVec_MPORT_1_en_pipe_0;
  assign tensorFile_1_rdataVec_MPORT_1_addr = tensorFile_1_rdataVec_MPORT_1_addr_pipe_0;
  assign tensorFile_1_rdataVec_MPORT_1_data = tensorFile_1[tensorFile_1_rdataVec_MPORT_1_addr]; // @[TensorLoadWideVME.scala 193:16]
  assign tensorFile_1_MPORT_1_data = _wmask_0_T ? 32'h0 : _wdata_1_T_2;
  assign tensorFile_1_MPORT_1_addr = widx_1[5:0];
  assign tensorFile_1_MPORT_1_mask = 1'h1;
  assign tensorFile_1_MPORT_1_en = _wmask_0_T ? 1'h0 : _wmask_1_T_4;
  assign io_done = loadDone & fillPadding_io_done; // @[TensorLoadWideVME.scala 316:25]
  assign io_vme_rd_cmd_valid = vmeCmd_io_vmeCmd_valid; // @[TensorLoadWideVME.scala 110:20]
  assign io_vme_rd_cmd_bits_addr = vmeCmd_io_vmeCmd_bits_addr; // @[TensorLoadWideVME.scala 110:20]
  assign io_vme_rd_cmd_bits_len = vmeCmd_io_vmeCmd_bits_len; // @[TensorLoadWideVME.scala 110:20]
  assign io_vme_rd_cmd_bits_tag = vmeCmd_io_vmeCmd_bits_tag; // @[TensorLoadWideVME.scala 110:20]
  assign io_vme_rd_data_ready = 1'h1; // @[TensorLoadWideVME.scala 156:24]
  assign io_tensor_rd_0_data_valid = rvalid; // @[TensorLoadWideVME.scala 311:37]
  assign io_tensor_rd_0_data_bits_0_0 = _rdata_T_2 | _rdata_T_3; // @[Mux.scala 27:73]
  assign vmeCmd_clock = clock;
  assign vmeCmd_reset = reset;
  assign vmeCmd_io_start = io_start; // @[TensorLoadWideVME.scala 106:19]
  assign vmeCmd_io_isBusy = state; // @[TensorLoadWideVME.scala 86:22]
  assign vmeCmd_io_inst = io_inst; // @[TensorLoadWideVME.scala 108:18]
  assign vmeCmd_io_baddr = io_baddr; // @[TensorLoadWideVME.scala 109:19]
  assign vmeCmd_io_vmeCmd_ready = io_vme_rd_cmd_ready; // @[TensorLoadWideVME.scala 110:20]
  assign readData_clock = clock;
  assign readData_reset = reset;
  assign readData_io_start = io_start; // @[TensorLoadWideVME.scala 151:21]
  assign readData_io_vmeData_valid = io_vme_rd_data_valid; // @[TensorLoadWideVME.scala 152:29]
  assign readData_io_vmeData_bits_data = io_vme_rd_data_bits_data; // @[TensorLoadWideVME.scala 153:28]
  assign readData_io_vmeData_bits_tag = io_vme_rd_data_bits_tag; // @[TensorLoadWideVME.scala 153:28]
  assign readData_io_vmeData_bits_last = io_vme_rd_data_bits_last; // @[TensorLoadWideVME.scala 153:28]
  assign fillPadding_clock = clock;
  assign fillPadding_reset = reset;
  assign fillPadding_io_canWriteMem = ~vmeDataFirePipe; // @[TensorLoadWideVME.scala 167:33]
  assign fillPadding_io_inst = io_inst; // @[TensorLoadWideVME.scala 168:23]
  assign fillPadding_io_start = io_start; // @[TensorLoadWideVME.scala 169:24]
  always @(posedge clock) begin
    if (tensorFile_0_MPORT_en & tensorFile_0_MPORT_mask) begin
      tensorFile_0[tensorFile_0_MPORT_addr] <= tensorFile_0_MPORT_data; // @[TensorLoadWideVME.scala 193:16]
    end
    tensorFile_0_rdataVec_MPORT_en_pipe_0 <= rMask[0];
    if (rMask[0]) begin
      tensorFile_0_rdataVec_MPORT_addr_pipe_0 <= io_tensor_rd_0_idx_bits[6:1];
    end
    if (tensorFile_1_MPORT_1_en & tensorFile_1_MPORT_1_mask) begin
      tensorFile_1[tensorFile_1_MPORT_1_addr] <= tensorFile_1_MPORT_1_data; // @[TensorLoadWideVME.scala 193:16]
    end
    tensorFile_1_rdataVec_MPORT_1_en_pipe_0 <= rMask[1];
    if (rMask[1]) begin
      tensorFile_1_rdataVec_MPORT_1_addr_pipe_0 <= io_tensor_rd_0_idx_bits[6:1];
    end
    if (reset) begin // @[TensorLoadWideVME.scala 84:22]
      state <= 1'h0; // @[TensorLoadWideVME.scala 84:22]
    end else begin
      state <= _GEN_1;
    end
    if (io_start) begin // @[TensorLoadWideVME.scala 133:18]
      clInFlight <= 7'h0; // @[TensorLoadWideVME.scala 134:16]
    end else if (state & _T & ~vmeDataFirePipe) begin // @[TensorLoadWideVME.scala 135:64]
      clInFlight <= _clInFlight_T_1; // @[TensorLoadWideVME.scala 136:16]
    end else if (_T_1 & vmeDataFirePipe) begin // @[TensorLoadWideVME.scala 137:63]
      clInFlight <= _clInFlight_T_5; // @[TensorLoadWideVME.scala 138:16]
    end else if (state & ~_T & vmeDataFirePipe) begin // @[TensorLoadWideVME.scala 139:64]
      clInFlight <= _clInFlight_T_7; // @[TensorLoadWideVME.scala 141:16]
    end
    if (io_tensor_rd_0_idx_valid) begin // @[TensorLoadWideVME.scala 290:10]
      rdata_r <= _rMask_T_1;
    end else begin
      rdata_r <= 2'h0;
    end
    if (reset) begin // @[Reg.scala 28:20]
      rvalid <= 1'h0; // @[Reg.scala 28:20]
    end else begin
      rvalid <= io_tensor_rd_0_idx_valid;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~io_start & ~_T_3 & ~_T_6 & _T_10 & ~reset & ~(clInFlight > 7'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TensorLoadWideVME.scala:140 assert(clInFlight > 0.U)\n"); // @[TensorLoadWideVME.scala 140:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_0[initvar] = _RAND_0[31:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tensorFile_1[initvar] = _RAND_3[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tensorFile_0_rdataVec_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  tensorFile_0_rdataVec_MPORT_addr_pipe_0 = _RAND_2[5:0];
  _RAND_4 = {1{`RANDOM}};
  tensorFile_1_rdataVec_MPORT_1_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  tensorFile_1_rdataVec_MPORT_1_addr_pipe_0 = _RAND_5[5:0];
  _RAND_6 = {1{`RANDOM}};
  state = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  clInFlight = _RAND_7[6:0];
  _RAND_8 = {1{`RANDOM}};
  rdata_r = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  rvalid = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~io_start & ~_T_3 & ~_T_6 & _T_10 & ~reset) begin
      assert(clInFlight > 7'h0); // @[TensorLoadWideVME.scala 140:11]
    end
    //
    if (_T_13) begin
      assert(1'h1); // @[TensorLoadWideVME.scala 154:9]
    end
  end
endmodule
module TensorLoadUop(
  input          clock,
  input          reset,
  input          io_start,
  output         io_done,
  input  [127:0] io_inst,
  input  [31:0]  io_baddr,
  input          io_vme_rd_cmd_ready,
  output         io_vme_rd_cmd_valid,
  output [31:0]  io_vme_rd_cmd_bits_addr,
  output [3:0]   io_vme_rd_cmd_bits_len,
  output [20:0]  io_vme_rd_cmd_bits_tag,
  input          io_vme_rd_data_valid,
  input  [63:0]  io_vme_rd_data_bits_data,
  input  [20:0]  io_vme_rd_data_bits_tag,
  input          io_vme_rd_data_bits_last,
  input          io_tensor_rd_0_idx_valid,
  input  [6:0]   io_tensor_rd_0_idx_bits,
  output         io_tensor_rd_0_data_valid,
  output [31:0]  io_tensor_rd_0_data_bits_0_0
);
  wire  tensorLoad_clock; // @[TensorLoad.scala 65:28]
  wire  tensorLoad_reset; // @[TensorLoad.scala 65:28]
  wire  tensorLoad_io_start; // @[TensorLoad.scala 65:28]
  wire  tensorLoad_io_done; // @[TensorLoad.scala 65:28]
  wire [127:0] tensorLoad_io_inst; // @[TensorLoad.scala 65:28]
  wire [31:0] tensorLoad_io_baddr; // @[TensorLoad.scala 65:28]
  wire  tensorLoad_io_vme_rd_cmd_ready; // @[TensorLoad.scala 65:28]
  wire  tensorLoad_io_vme_rd_cmd_valid; // @[TensorLoad.scala 65:28]
  wire [31:0] tensorLoad_io_vme_rd_cmd_bits_addr; // @[TensorLoad.scala 65:28]
  wire [3:0] tensorLoad_io_vme_rd_cmd_bits_len; // @[TensorLoad.scala 65:28]
  wire [20:0] tensorLoad_io_vme_rd_cmd_bits_tag; // @[TensorLoad.scala 65:28]
  wire  tensorLoad_io_vme_rd_data_ready; // @[TensorLoad.scala 65:28]
  wire  tensorLoad_io_vme_rd_data_valid; // @[TensorLoad.scala 65:28]
  wire [63:0] tensorLoad_io_vme_rd_data_bits_data; // @[TensorLoad.scala 65:28]
  wire [20:0] tensorLoad_io_vme_rd_data_bits_tag; // @[TensorLoad.scala 65:28]
  wire  tensorLoad_io_vme_rd_data_bits_last; // @[TensorLoad.scala 65:28]
  wire  tensorLoad_io_tensor_rd_0_idx_valid; // @[TensorLoad.scala 65:28]
  wire [6:0] tensorLoad_io_tensor_rd_0_idx_bits; // @[TensorLoad.scala 65:28]
  wire  tensorLoad_io_tensor_rd_0_data_valid; // @[TensorLoad.scala 65:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_0; // @[TensorLoad.scala 65:28]
  TensorLoadWideVME tensorLoad ( // @[TensorLoad.scala 65:28]
    .clock(tensorLoad_clock),
    .reset(tensorLoad_reset),
    .io_start(tensorLoad_io_start),
    .io_done(tensorLoad_io_done),
    .io_inst(tensorLoad_io_inst),
    .io_baddr(tensorLoad_io_baddr),
    .io_vme_rd_cmd_ready(tensorLoad_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(tensorLoad_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(tensorLoad_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(tensorLoad_io_vme_rd_cmd_bits_len),
    .io_vme_rd_cmd_bits_tag(tensorLoad_io_vme_rd_cmd_bits_tag),
    .io_vme_rd_data_ready(tensorLoad_io_vme_rd_data_ready),
    .io_vme_rd_data_valid(tensorLoad_io_vme_rd_data_valid),
    .io_vme_rd_data_bits_data(tensorLoad_io_vme_rd_data_bits_data),
    .io_vme_rd_data_bits_tag(tensorLoad_io_vme_rd_data_bits_tag),
    .io_vme_rd_data_bits_last(tensorLoad_io_vme_rd_data_bits_last),
    .io_tensor_rd_0_idx_valid(tensorLoad_io_tensor_rd_0_idx_valid),
    .io_tensor_rd_0_idx_bits(tensorLoad_io_tensor_rd_0_idx_bits),
    .io_tensor_rd_0_data_valid(tensorLoad_io_tensor_rd_0_data_valid),
    .io_tensor_rd_0_data_bits_0_0(tensorLoad_io_tensor_rd_0_data_bits_0_0)
  );
  assign io_done = tensorLoad_io_done; // @[TensorLoad.scala 66:8]
  assign io_vme_rd_cmd_valid = tensorLoad_io_vme_rd_cmd_valid; // @[TensorLoad.scala 66:8]
  assign io_vme_rd_cmd_bits_addr = tensorLoad_io_vme_rd_cmd_bits_addr; // @[TensorLoad.scala 66:8]
  assign io_vme_rd_cmd_bits_len = tensorLoad_io_vme_rd_cmd_bits_len; // @[TensorLoad.scala 66:8]
  assign io_vme_rd_cmd_bits_tag = tensorLoad_io_vme_rd_cmd_bits_tag; // @[TensorLoad.scala 66:8]
  assign io_tensor_rd_0_data_valid = tensorLoad_io_tensor_rd_0_data_valid; // @[TensorLoad.scala 66:8]
  assign io_tensor_rd_0_data_bits_0_0 = tensorLoad_io_tensor_rd_0_data_bits_0_0; // @[TensorLoad.scala 66:8]
  assign tensorLoad_clock = clock;
  assign tensorLoad_reset = reset;
  assign tensorLoad_io_start = io_start; // @[TensorLoad.scala 66:8]
  assign tensorLoad_io_inst = io_inst; // @[TensorLoad.scala 66:8]
  assign tensorLoad_io_baddr = io_baddr; // @[TensorLoad.scala 66:8]
  assign tensorLoad_io_vme_rd_cmd_ready = io_vme_rd_cmd_ready; // @[TensorLoad.scala 66:8]
  assign tensorLoad_io_vme_rd_data_valid = io_vme_rd_data_valid; // @[TensorLoad.scala 66:8]
  assign tensorLoad_io_vme_rd_data_bits_data = io_vme_rd_data_bits_data; // @[TensorLoad.scala 66:8]
  assign tensorLoad_io_vme_rd_data_bits_tag = io_vme_rd_data_bits_tag; // @[TensorLoad.scala 66:8]
  assign tensorLoad_io_vme_rd_data_bits_last = io_vme_rd_data_bits_last; // @[TensorLoad.scala 66:8]
  assign tensorLoad_io_tensor_rd_0_idx_valid = io_tensor_rd_0_idx_valid; // @[TensorLoad.scala 66:8]
  assign tensorLoad_io_tensor_rd_0_idx_bits = io_tensor_rd_0_idx_bits; // @[TensorLoad.scala 66:8]
endmodule
module LoadUopTop(
  input          clock,
  input          reset,
  input          io_start,
  output         io_done,
  input  [127:0] io_inst,
  input  [31:0]  io_baddr,
  input          io_vme_rd_cmd_ready,
  output         io_vme_rd_cmd_valid,
  output [31:0]  io_vme_rd_cmd_bits_addr,
  output [3:0]   io_vme_rd_cmd_bits_len,
  output [20:0]  io_vme_rd_cmd_bits_tag,
  input          io_vme_rd_data_valid,
  input  [63:0]  io_vme_rd_data_bits_data,
  input  [20:0]  io_vme_rd_data_bits_tag,
  input          io_vme_rd_data_bits_last,
  input          io_uop_idx_valid,
  input  [6:0]   io_uop_idx_bits,
  output         io_uop_data_valid,
  output [9:0]   io_uop_data_bits_u2,
  output [10:0]  io_uop_data_bits_u1,
  output [10:0]  io_uop_data_bits_u0
);
  wire  loadUop_clock; // @[LoadUop.scala 85:25]
  wire  loadUop_reset; // @[LoadUop.scala 85:25]
  wire  loadUop_io_start; // @[LoadUop.scala 85:25]
  wire  loadUop_io_done; // @[LoadUop.scala 85:25]
  wire [127:0] loadUop_io_inst; // @[LoadUop.scala 85:25]
  wire [31:0] loadUop_io_baddr; // @[LoadUop.scala 85:25]
  wire  loadUop_io_vme_rd_cmd_ready; // @[LoadUop.scala 85:25]
  wire  loadUop_io_vme_rd_cmd_valid; // @[LoadUop.scala 85:25]
  wire [31:0] loadUop_io_vme_rd_cmd_bits_addr; // @[LoadUop.scala 85:25]
  wire [3:0] loadUop_io_vme_rd_cmd_bits_len; // @[LoadUop.scala 85:25]
  wire [20:0] loadUop_io_vme_rd_cmd_bits_tag; // @[LoadUop.scala 85:25]
  wire  loadUop_io_vme_rd_data_valid; // @[LoadUop.scala 85:25]
  wire [63:0] loadUop_io_vme_rd_data_bits_data; // @[LoadUop.scala 85:25]
  wire [20:0] loadUop_io_vme_rd_data_bits_tag; // @[LoadUop.scala 85:25]
  wire  loadUop_io_vme_rd_data_bits_last; // @[LoadUop.scala 85:25]
  wire  loadUop_io_tensor_rd_0_idx_valid; // @[LoadUop.scala 85:25]
  wire [6:0] loadUop_io_tensor_rd_0_idx_bits; // @[LoadUop.scala 85:25]
  wire  loadUop_io_tensor_rd_0_data_valid; // @[LoadUop.scala 85:25]
  wire [31:0] loadUop_io_tensor_rd_0_data_bits_0_0; // @[LoadUop.scala 85:25]
  wire [31:0] _io_uop_data_bits_WIRE_1 = loadUop_io_tensor_rd_0_data_bits_0_0;
  TensorLoadUop loadUop ( // @[LoadUop.scala 85:25]
    .clock(loadUop_clock),
    .reset(loadUop_reset),
    .io_start(loadUop_io_start),
    .io_done(loadUop_io_done),
    .io_inst(loadUop_io_inst),
    .io_baddr(loadUop_io_baddr),
    .io_vme_rd_cmd_ready(loadUop_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(loadUop_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(loadUop_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(loadUop_io_vme_rd_cmd_bits_len),
    .io_vme_rd_cmd_bits_tag(loadUop_io_vme_rd_cmd_bits_tag),
    .io_vme_rd_data_valid(loadUop_io_vme_rd_data_valid),
    .io_vme_rd_data_bits_data(loadUop_io_vme_rd_data_bits_data),
    .io_vme_rd_data_bits_tag(loadUop_io_vme_rd_data_bits_tag),
    .io_vme_rd_data_bits_last(loadUop_io_vme_rd_data_bits_last),
    .io_tensor_rd_0_idx_valid(loadUop_io_tensor_rd_0_idx_valid),
    .io_tensor_rd_0_idx_bits(loadUop_io_tensor_rd_0_idx_bits),
    .io_tensor_rd_0_data_valid(loadUop_io_tensor_rd_0_data_valid),
    .io_tensor_rd_0_data_bits_0_0(loadUop_io_tensor_rd_0_data_bits_0_0)
  );
  assign io_done = loadUop_io_done; // @[LoadUop.scala 89:13]
  assign io_vme_rd_cmd_valid = loadUop_io_vme_rd_cmd_valid; // @[LoadUop.scala 91:23]
  assign io_vme_rd_cmd_bits_addr = loadUop_io_vme_rd_cmd_bits_addr; // @[LoadUop.scala 91:23]
  assign io_vme_rd_cmd_bits_len = loadUop_io_vme_rd_cmd_bits_len; // @[LoadUop.scala 91:23]
  assign io_vme_rd_cmd_bits_tag = loadUop_io_vme_rd_cmd_bits_tag; // @[LoadUop.scala 91:23]
  assign io_uop_data_valid = loadUop_io_tensor_rd_0_data_valid; // @[LoadUop.scala 96:23]
  assign io_uop_data_bits_u2 = _io_uop_data_bits_WIRE_1[31:22]; // @[LoadUop.scala 97:67]
  assign io_uop_data_bits_u1 = _io_uop_data_bits_WIRE_1[21:11]; // @[LoadUop.scala 97:67]
  assign io_uop_data_bits_u0 = _io_uop_data_bits_WIRE_1[10:0]; // @[LoadUop.scala 97:67]
  assign loadUop_clock = clock;
  assign loadUop_reset = reset;
  assign loadUop_io_start = io_start; // @[LoadUop.scala 88:22]
  assign loadUop_io_inst = io_inst; // @[LoadUop.scala 93:21]
  assign loadUop_io_baddr = io_baddr; // @[LoadUop.scala 90:22]
  assign loadUop_io_vme_rd_cmd_ready = io_vme_rd_cmd_ready; // @[LoadUop.scala 91:23]
  assign loadUop_io_vme_rd_data_valid = io_vme_rd_data_valid; // @[LoadUop.scala 91:23]
  assign loadUop_io_vme_rd_data_bits_data = io_vme_rd_data_bits_data; // @[LoadUop.scala 91:23]
  assign loadUop_io_vme_rd_data_bits_tag = io_vme_rd_data_bits_tag; // @[LoadUop.scala 91:23]
  assign loadUop_io_vme_rd_data_bits_last = io_vme_rd_data_bits_last; // @[LoadUop.scala 91:23]
  assign loadUop_io_tensor_rd_0_idx_valid = io_uop_idx_valid; // @[LoadUop.scala 95:33]
  assign loadUop_io_tensor_rd_0_idx_bits = io_uop_idx_bits; // @[LoadUop.scala 95:33]
endmodule
module GenVMECmd_2(
  input          clock,
  input          reset,
  input          io_start,
  input          io_isBusy,
  input  [127:0] io_inst,
  input  [31:0]  io_baddr,
  input          io_vmeCmd_ready,
  output         io_vmeCmd_valid,
  output [31:0]  io_vmeCmd_bits_addr,
  output [3:0]   io_vmeCmd_bits_len,
  output [20:0]  io_vmeCmd_bits_tag,
  output [4:0]   io_readLen,
  output         io_done
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  wire [15:0] dec_sram_offset = io_inst[25:10]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [31:0] dec_dram_offset = io_inst[57:26]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [15:0] dec_ysize = io_inst[79:64]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [15:0] dec_xsize = io_inst[95:80]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [15:0] dec_xstride = io_inst[111:96]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [3:0] dec_ypad_0 = io_inst[115:112]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [3:0] dec_xpad_0 = io_inst[123:120]; // @[TensorLoadNarrowVME.scala 566:29]
  wire [3:0] dec_xpad_1 = io_inst[127:124]; // @[TensorLoadNarrowVME.scala 566:29]
  reg [31:0] rdCmdExtAddr; // @[TensorLoadNarrowVME.scala 568:25]
  wire [38:0] _xfer_init_addr_T = {dec_dram_offset, 7'h0}; // @[TensorLoadNarrowVME.scala 573:66]
  wire [38:0] _xfer_init_addr_T_1 = 39'hffffffff & _xfer_init_addr_T; // @[TensorLoadNarrowVME.scala 573:47]
  wire [38:0] _GEN_31 = {{7'd0}, io_baddr}; // @[TensorLoadNarrowVME.scala 573:33]
  wire [38:0] xfer_init_addr = _GEN_31 | _xfer_init_addr_T_1; // @[TensorLoadNarrowVME.scala 573:33]
  wire [31:0] _GEN_0 = rdCmdExtAddr % 32'h80; // @[TensorLoadNarrowVME.scala 577:53]
  wire [7:0] _firstMaxTransfer_T = _GEN_0[7:0]; // @[TensorLoadNarrowVME.scala 577:53]
  wire [7:0] _firstMaxTransfer_T_2 = 8'h80 - _firstMaxTransfer_T; // @[TensorLoadNarrowVME.scala 577:38]
  wire [4:0] firstMaxTransfer = _firstMaxTransfer_T_2[7:3]; // @[TensorLoadNarrowVME.scala 577:67]
  reg [6:0] rdCmdStartIdx; // @[TensorLoadNarrowVME.scala 586:26]
  reg  commandsDone; // @[TensorLoadNarrowVME.scala 588:29]
  wire [19:0] blocksReadSize = {dec_xsize, 4'h0}; // @[TensorLoadNarrowVME.scala 590:35]
  reg [19:0] blocksReadNb; // @[TensorLoadNarrowVME.scala 591:25]
  reg [31:0] rdCmdExtAddrRowBegin; // @[TensorLoadNarrowVME.scala 592:33]
  reg  newReadRow; // @[TensorLoadNarrowVME.scala 593:23]
  reg [15:0] srcRowIdx; // @[TensorLoadNarrowVME.scala 596:22]
  wire [15:0] _srcRowIdx_T_1 = srcRowIdx + 16'h1; // @[TensorLoadNarrowVME.scala 600:28]
  wire [19:0] blocksRemained = blocksReadSize - blocksReadNb; // @[TensorLoadNarrowVME.scala 628:39]
  wire [19:0] _GEN_32 = {{15'd0}, firstMaxTransfer}; // @[TensorLoadNarrowVME.scala 630:25]
  wire [19:0] _GEN_8 = blocksRemained < _GEN_32 ? blocksRemained : {{15'd0}, firstMaxTransfer}; // @[TensorLoadNarrowVME.scala 630:45 631:15 633:15]
  wire [19:0] _GEN_9 = blocksRemained < 20'h10 ? blocksRemained : 20'h10; // @[TensorLoadNarrowVME.scala 636:40 637:15 639:15]
  wire [19:0] _GEN_10 = newReadRow ? _GEN_8 : _GEN_9; // @[TensorLoadNarrowVME.scala 629:21]
  wire [4:0] readLen = _GEN_10[4:0]; // @[TensorLoadNarrowVME.scala 587:21]
  wire [19:0] _GEN_33 = {{15'd0}, readLen}; // @[TensorLoadNarrowVME.scala 621:41]
  wire [19:0] _T_8 = blocksReadSize - _GEN_33; // @[TensorLoadNarrowVME.scala 621:41]
  wire [15:0] _T_11 = dec_ysize - 16'h1; // @[TensorLoadNarrowVME.scala 621:80]
  wire  _T_14 = io_vmeCmd_ready & io_vmeCmd_valid; // @[Decoupled.scala 50:35]
  wire  stride = blocksReadNb == _T_8 & srcRowIdx != _T_11 & _T_14; // @[TensorLoadNarrowVME.scala 621:87]
  wire [19:0] nextBlRNb = blocksReadNb + _GEN_33; // @[TensorLoadNarrowVME.scala 611:34]
  wire  _GEN_2 = nextBlRNb == blocksReadSize & srcRowIdx == _T_11 | commandsDone; // @[TensorLoadNarrowVME.scala 606:16 613:74 614:20]
  wire  _GEN_4 = _T_14 ? _GEN_2 : commandsDone; // @[TensorLoadNarrowVME.scala 606:16 610:31]
  wire  _GEN_6 = io_start | stride ? 1'h0 : _GEN_4; // @[TensorLoadNarrowVME.scala 607:29 609:18]
  wire  _T_20 = ~reset; // @[TensorLoadNarrowVME.scala 627:9]
  wire [15:0] _GEN_35 = {{12'd0}, dec_xpad_0}; // @[TensorLoadNarrowVME.scala 643:30]
  wire [15:0] _totalWidth_T_1 = dec_xsize + _GEN_35; // @[TensorLoadNarrowVME.scala 643:30]
  wire [15:0] _GEN_36 = {{12'd0}, dec_xpad_1}; // @[TensorLoadNarrowVME.scala 643:43]
  wire [15:0] totalWidth = _totalWidth_T_1 + _GEN_36; // @[TensorLoadNarrowVME.scala 643:43]
  reg [19:0] currentRowIdx; // @[TensorLoadNarrowVME.scala 647:26]
  wire [19:0] _GEN_37 = {{16'd0}, dec_ypad_0}; // @[TensorLoadNarrowVME.scala 649:39]
  wire [15:0] _GEN_38 = {{12'd0}, dec_ypad_0}; // @[TensorLoadNarrowVME.scala 650:32]
  wire [15:0] _rdCmdStartIdxValid_T_2 = dec_ysize + _GEN_38; // @[TensorLoadNarrowVME.scala 650:32]
  wire [19:0] _GEN_39 = {{4'd0}, _rdCmdStartIdxValid_T_2}; // @[TensorLoadNarrowVME.scala 650:19]
  wire  _rdCmdStartIdxValid_T_3 = currentRowIdx < _GEN_39; // @[TensorLoadNarrowVME.scala 650:19]
  wire  _rdCmdStartIdxValid_T_4 = currentRowIdx >= _GEN_37 & _rdCmdStartIdxValid_T_3; // @[TensorLoadNarrowVME.scala 649:53]
  wire  _rdCmdStartIdxValid_T_5 = _rdCmdStartIdxValid_T_4 & io_isBusy; // @[TensorLoadNarrowVME.scala 650:46]
  wire  _rdCmdStartIdxValid_T_6 = ~commandsDone; // @[TensorLoadNarrowVME.scala 652:5]
  wire  rdCmdStartIdxValid = _rdCmdStartIdxValid_T_5 & _rdCmdStartIdxValid_T_6; // @[TensorLoadNarrowVME.scala 651:15]
  wire [15:0] _rdCmdStartIdx_T_1 = dec_sram_offset + _GEN_35; // @[TensorLoadNarrowVME.scala 655:38]
  wire [15:0] _GEN_42 = {{9'd0}, rdCmdStartIdx}; // @[TensorLoadNarrowVME.scala 657:36]
  wire [15:0] _rdCmdStartIdx_T_3 = _GEN_42 + totalWidth; // @[TensorLoadNarrowVME.scala 657:36]
  wire [19:0] _currentRowIdx_T_1 = currentRowIdx + 20'h1; // @[TensorLoadNarrowVME.scala 658:36]
  wire [15:0] _GEN_11 = io_isBusy & (currentRowIdx < _GEN_37 | stride) ? _rdCmdStartIdx_T_3 : {{9'd0}, rdCmdStartIdx}; // @[TensorLoadNarrowVME.scala 656:68 657:19 586:26]
  wire [15:0] _GEN_14 = io_start ? _rdCmdStartIdx_T_1 : _GEN_11; // @[TensorLoadNarrowVME.scala 653:19 655:19]
  wire  startIssueCmdRead = blocksReadNb == 20'h0 & rdCmdStartIdxValid; // @[TensorLoadNarrowVME.scala 661:29]
  wire [22:0] _memRow_T = {dec_xstride, 7'h0}; // @[TensorLoadNarrowVME.scala 672:56]
  wire [31:0] _GEN_43 = {{9'd0}, _memRow_T}; // @[TensorLoadNarrowVME.scala 672:41]
  wire [31:0] memRow = rdCmdExtAddrRowBegin + _GEN_43; // @[TensorLoadNarrowVME.scala 672:41]
  wire [7:0] _rdCmdExtAddr_T = {readLen, 3'h0}; // @[TensorLoadNarrowVME.scala 679:47]
  wire [31:0] _GEN_44 = {{24'd0}, _rdCmdExtAddr_T}; // @[TensorLoadNarrowVME.scala 679:36]
  wire [31:0] _rdCmdExtAddr_T_2 = rdCmdExtAddr + _GEN_44; // @[TensorLoadNarrowVME.scala 679:36]
  wire [31:0] _GEN_16 = stride ? memRow : _rdCmdExtAddr_T_2; // @[TensorLoadNarrowVME.scala 671:18 673:20 679:20]
  wire [31:0] _GEN_17 = stride ? memRow : rdCmdExtAddrRowBegin; // @[TensorLoadNarrowVME.scala 671:18 664:24 674:28]
  wire [31:0] _GEN_19 = _T_14 ? _GEN_16 : rdCmdExtAddr; // @[TensorLoadNarrowVME.scala 670:31 682:18]
  wire [31:0] _GEN_20 = _T_14 ? _GEN_17 : rdCmdExtAddrRowBegin; // @[TensorLoadNarrowVME.scala 664:24 670:31]
  wire  _GEN_21 = _T_14 ? stride : newReadRow; // @[TensorLoadNarrowVME.scala 670:31 683:16]
  wire [38:0] _GEN_22 = io_start ? xfer_init_addr : {{7'd0}, _GEN_19}; // @[TensorLoadNarrowVME.scala 666:19 667:18]
  wire [38:0] _GEN_23 = io_start ? xfer_init_addr : {{7'd0}, _GEN_20}; // @[TensorLoadNarrowVME.scala 666:19 668:26]
  reg [10:0] rdCmdDestBlockIdxNext; // @[TensorLoadNarrowVME.scala 700:34]
  wire [10:0] _rdCmdDestBlockIdx_T = {rdCmdStartIdx, 4'h0}; // @[TensorLoadNarrowVME.scala 710:42]
  wire [10:0] _GEN_26 = startIssueCmdRead ? _rdCmdDestBlockIdx_T : rdCmdDestBlockIdxNext; // @[TensorLoadNarrowVME.scala 702:21 709:29 710:25]
  wire [10:0] rdCmdDestBlockIdx = rdCmdStartIdxValid ? _GEN_26 : rdCmdDestBlockIdxNext; // @[TensorLoadNarrowVME.scala 702:21 707:28]
  wire [10:0] _GEN_45 = {{6'd0}, readLen}; // @[TensorLoadNarrowVME.scala 711:49]
  wire [10:0] _rdCmdDestBlockIdxNext_T_1 = rdCmdDestBlockIdx + _GEN_45; // @[TensorLoadNarrowVME.scala 711:49]
  wire [10:0] _rdCmdDestBlockIdxNext_T_3 = rdCmdDestBlockIdxNext + _GEN_45; // @[TensorLoadNarrowVME.scala 714:53]
  wire [4:0] _io_vmeCmd_bits_len_T_1 = readLen - 5'h1; // @[TensorLoadNarrowVME.scala 732:33]
  assign io_vmeCmd_valid = _rdCmdStartIdxValid_T_5 & _rdCmdStartIdxValid_T_6; // @[TensorLoadNarrowVME.scala 651:15]
  assign io_vmeCmd_bits_addr = rdCmdExtAddr; // @[TensorLoadNarrowVME.scala 731:23]
  assign io_vmeCmd_bits_len = _io_vmeCmd_bits_len_T_1[3:0]; // @[TensorLoadNarrowVME.scala 732:22]
  assign io_vmeCmd_bits_tag = {{10'd0}, rdCmdDestBlockIdx}; // @[TensorLoadNarrowVME.scala 737:22]
  assign io_readLen = _GEN_10[4:0]; // @[TensorLoadNarrowVME.scala 587:21]
  assign io_done = commandsDone; // @[TensorLoadNarrowVME.scala 739:11]
  always @(posedge clock) begin
    rdCmdExtAddr <= _GEN_22[31:0];
    rdCmdStartIdx <= _GEN_14[6:0];
    commandsDone <= reset | _GEN_6; // @[TensorLoadNarrowVME.scala 588:{29,29}]
    if (io_start | stride) begin // @[TensorLoadNarrowVME.scala 607:29]
      blocksReadNb <= 20'h0; // @[TensorLoadNarrowVME.scala 608:18]
    end else if (_T_14) begin // @[TensorLoadNarrowVME.scala 610:31]
      blocksReadNb <= nextBlRNb; // @[TensorLoadNarrowVME.scala 612:18]
    end
    rdCmdExtAddrRowBegin <= _GEN_23[31:0];
    newReadRow <= io_start | _GEN_21; // @[TensorLoadNarrowVME.scala 666:19 669:16]
    if (io_start) begin // @[TensorLoadNarrowVME.scala 597:19]
      srcRowIdx <= 16'h0; // @[TensorLoadNarrowVME.scala 598:15]
    end else if (stride) begin // @[TensorLoadNarrowVME.scala 599:23]
      srcRowIdx <= _srcRowIdx_T_1; // @[TensorLoadNarrowVME.scala 600:15]
    end
    if (io_start) begin // @[TensorLoadNarrowVME.scala 653:19]
      currentRowIdx <= 20'h0; // @[TensorLoadNarrowVME.scala 654:19]
    end else if (io_isBusy & (currentRowIdx < _GEN_37 | stride)) begin // @[TensorLoadNarrowVME.scala 656:68]
      currentRowIdx <= _currentRowIdx_T_1; // @[TensorLoadNarrowVME.scala 658:19]
    end
    if (rdCmdStartIdxValid) begin // @[TensorLoadNarrowVME.scala 707:28]
      if (startIssueCmdRead) begin // @[TensorLoadNarrowVME.scala 709:29]
        rdCmdDestBlockIdxNext <= _rdCmdDestBlockIdxNext_T_1; // @[TensorLoadNarrowVME.scala 711:28]
      end else if (_T_14) begin // @[TensorLoadNarrowVME.scala 712:33]
        rdCmdDestBlockIdxNext <= _rdCmdDestBlockIdxNext_T_3; // @[TensorLoadNarrowVME.scala 714:28]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~io_isBusy | blocksReadSize >= blocksReadNb)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorLoadNarrowVME.scala:627 assert(!io.isBusy || blocksReadSize >= blocksReadNb)// define how many block to read at this cycle\n"
            ); // @[TensorLoadNarrowVME.scala 627:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_20 & ~(~io_vmeCmd_valid | _rdCmdExtAddr_T <= _firstMaxTransfer_T_2)) begin
          $fwrite(32'h80000002,
            "Assertion failed: -F- acc DRAM page alignment failure. DRAM address + len overlaps mp.lenBits*memBlockSize alignment %x %x\n    at TensorLoadNarrowVME.scala:733 assert(!io.vmeCmd.valid || ((readLen << log2Ceil(mp.dataBits/8)) <= (maxTrBytes - rdCmdExtAddr %% maxTrBytes)),\n"
            ,rdCmdExtAddr,readLen); // @[TensorLoadNarrowVME.scala 733:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rdCmdExtAddr = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  rdCmdStartIdx = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  commandsDone = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  blocksReadNb = _RAND_3[19:0];
  _RAND_4 = {1{`RANDOM}};
  rdCmdExtAddrRowBegin = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  newReadRow = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  srcRowIdx = _RAND_6[15:0];
  _RAND_7 = {1{`RANDOM}};
  currentRowIdx = _RAND_7[19:0];
  _RAND_8 = {1{`RANDOM}};
  rdCmdDestBlockIdxNext = _RAND_8[10:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~io_isBusy | blocksReadSize >= blocksReadNb); // @[TensorLoadNarrowVME.scala 627:9]
    end
    //
    if (_T_20) begin
      assert(~io_vmeCmd_valid | _rdCmdExtAddr_T <= _firstMaxTransfer_T_2); // @[TensorLoadNarrowVME.scala 733:9]
    end
  end
endmodule
module ReadVMEData_2(
  input         clock,
  input         reset,
  input         io_start,
  output        io_vmeData_ready,
  input         io_vmeData_valid,
  input  [20:0] io_vmeData_bits_tag,
  output [6:0]  io_idx,
  output [3:0]  io_col
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [20:0] vmeTagDecodeLast; // @[TensorLoadNarrowVME.scala 502:29]
  wire [16:0] rdDataIdx = io_vmeData_bits_tag[20:4]; // @[TensorLoadNarrowVME.scala 503:31]
  wire [3:0] rdDataCol = io_vmeData_bits_tag[3:0]; // @[TensorLoadNarrowVME.scala 504:65]
  reg [3:0] rdDataDestColNext; // @[TensorLoadNarrowVME.scala 505:30]
  reg [15:0] rdDataDestIdxNext; // @[TensorLoadNarrowVME.scala 506:30]
  reg  vmeTagDecodeLastValidNext; // @[TensorLoadNarrowVME.scala 509:42]
  wire  _T = io_vmeData_ready & io_vmeData_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_0 = _T | vmeTagDecodeLastValidNext; // @[TensorLoadNarrowVME.scala 514:31 515:27 517:27]
  wire  _T_3 = io_vmeData_bits_tag != vmeTagDecodeLast; // @[TensorLoadNarrowVME.scala 525:29]
  wire  _T_4 = vmeTagDecodeLastValidNext & _T_3; // @[TensorLoadNarrowVME.scala 524:34]
  wire  _T_5 = ~vmeTagDecodeLastValidNext | _T_4; // @[TensorLoadNarrowVME.scala 523:34]
  wire [3:0] _rdDataDestColNext_T_1 = rdDataCol + 4'h1; // @[TensorLoadNarrowVME.scala 530:38]
  wire [3:0] _rdDataDestColNext_T_3 = rdDataDestColNext + 4'h1; // @[TensorLoadNarrowVME.scala 534:46]
  wire [3:0] rdDataDestCol = _T_5 ? rdDataCol : rdDataDestColNext; // @[TensorLoadNarrowVME.scala 525:59 528:21 533:21]
  wire [15:0] _rdDataDestIdxNext_T_1 = rdDataDestIdxNext + 16'h1; // @[TensorLoadNarrowVME.scala 537:48]
  wire [15:0] _GEN_2 = rdDataDestCol == 4'hf ? _rdDataDestIdxNext_T_1 : rdDataDestIdxNext; // @[TensorLoadNarrowVME.scala 536:54 537:27 506:30]
  wire [16:0] _GEN_5 = _T_5 ? rdDataIdx : {{1'd0}, rdDataDestIdxNext}; // @[TensorLoadNarrowVME.scala 525:59 529:21 535:21]
  wire [16:0] _GEN_7 = _T_5 ? rdDataIdx : {{1'd0}, _GEN_2}; // @[TensorLoadNarrowVME.scala 525:59 531:25]
  wire [16:0] _GEN_12 = _T ? _GEN_7 : {{1'd0}, rdDataDestIdxNext}; // @[TensorLoadNarrowVME.scala 521:25 506:30]
  wire [15:0] rdDataDestIdx = _GEN_5[15:0]; // @[TensorLoadNarrowVME.scala 497:27]
  assign io_vmeData_ready = 1'h1; // @[TensorLoadNarrowVME.scala 498:20]
  assign io_idx = rdDataDestIdx[6:0]; // @[TensorLoadNarrowVME.scala 542:10]
  assign io_col = _T_5 ? rdDataCol : rdDataDestColNext; // @[TensorLoadNarrowVME.scala 525:59 528:21 533:21]
  always @(posedge clock) begin
    if (_T) begin // @[TensorLoadNarrowVME.scala 521:25]
      if (_T_5) begin // @[TensorLoadNarrowVME.scala 525:59]
        vmeTagDecodeLast <= io_vmeData_bits_tag; // @[TensorLoadNarrowVME.scala 527:24]
      end
    end
    if (_T) begin // @[TensorLoadNarrowVME.scala 521:25]
      if (_T_5) begin // @[TensorLoadNarrowVME.scala 525:59]
        rdDataDestColNext <= _rdDataDestColNext_T_1; // @[TensorLoadNarrowVME.scala 530:25]
      end else begin
        rdDataDestColNext <= _rdDataDestColNext_T_3; // @[TensorLoadNarrowVME.scala 534:25]
      end
    end
    rdDataDestIdxNext <= _GEN_12[15:0];
    if (reset) begin // @[TensorLoadNarrowVME.scala 509:42]
      vmeTagDecodeLastValidNext <= 1'h0; // @[TensorLoadNarrowVME.scala 509:42]
    end else if (io_start) begin // @[TensorLoadNarrowVME.scala 512:18]
      vmeTagDecodeLastValidNext <= 1'h0; // @[TensorLoadNarrowVME.scala 513:27]
    end else begin
      vmeTagDecodeLastValidNext <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  vmeTagDecodeLast = _RAND_0[20:0];
  _RAND_1 = {1{`RANDOM}};
  rdDataDestColNext = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  rdDataDestIdxNext = _RAND_2[15:0];
  _RAND_3 = {1{`RANDOM}};
  vmeTagDecodeLastValidNext = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TensorLoadNarrowVME_2(
  input          clock,
  input          reset,
  input          io_start,
  output         io_done,
  input  [127:0] io_inst,
  input  [31:0]  io_baddr,
  input          io_vme_rd_cmd_ready,
  output         io_vme_rd_cmd_valid,
  output [31:0]  io_vme_rd_cmd_bits_addr,
  output [3:0]   io_vme_rd_cmd_bits_len,
  output [20:0]  io_vme_rd_cmd_bits_tag,
  output         io_vme_rd_data_ready,
  input          io_vme_rd_data_valid,
  input  [63:0]  io_vme_rd_data_bits_data,
  input  [20:0]  io_vme_rd_data_bits_tag,
  input          io_tensor_rd_0_idx_valid,
  input  [6:0]   io_tensor_rd_0_idx_bits,
  output         io_tensor_rd_0_data_valid,
  output [31:0]  io_tensor_rd_0_data_bits_0_0,
  output [31:0]  io_tensor_rd_0_data_bits_0_1,
  output [31:0]  io_tensor_rd_0_data_bits_0_2,
  output [31:0]  io_tensor_rd_0_data_bits_0_3,
  output [31:0]  io_tensor_rd_0_data_bits_0_4,
  output [31:0]  io_tensor_rd_0_data_bits_0_5,
  output [31:0]  io_tensor_rd_0_data_bits_0_6,
  output [31:0]  io_tensor_rd_0_data_bits_0_7,
  output [31:0]  io_tensor_rd_0_data_bits_0_8,
  output [31:0]  io_tensor_rd_0_data_bits_0_9,
  output [31:0]  io_tensor_rd_0_data_bits_0_10,
  output [31:0]  io_tensor_rd_0_data_bits_0_11,
  output [31:0]  io_tensor_rd_0_data_bits_0_12,
  output [31:0]  io_tensor_rd_0_data_bits_0_13,
  output [31:0]  io_tensor_rd_0_data_bits_0_14,
  output [31:0]  io_tensor_rd_0_data_bits_0_15,
  output [31:0]  io_tensor_rd_0_data_bits_0_16,
  output [31:0]  io_tensor_rd_0_data_bits_0_17,
  output [31:0]  io_tensor_rd_0_data_bits_0_18,
  output [31:0]  io_tensor_rd_0_data_bits_0_19,
  output [31:0]  io_tensor_rd_0_data_bits_0_20,
  output [31:0]  io_tensor_rd_0_data_bits_0_21,
  output [31:0]  io_tensor_rd_0_data_bits_0_22,
  output [31:0]  io_tensor_rd_0_data_bits_0_23,
  output [31:0]  io_tensor_rd_0_data_bits_0_24,
  output [31:0]  io_tensor_rd_0_data_bits_0_25,
  output [31:0]  io_tensor_rd_0_data_bits_0_26,
  output [31:0]  io_tensor_rd_0_data_bits_0_27,
  output [31:0]  io_tensor_rd_0_data_bits_0_28,
  output [31:0]  io_tensor_rd_0_data_bits_0_29,
  output [31:0]  io_tensor_rd_0_data_bits_0_30,
  output [31:0]  io_tensor_rd_0_data_bits_0_31,
  input          io_tensor_wr_0_valid,
  input  [6:0]   io_tensor_wr_0_bits_idx,
  input  [31:0]  io_tensor_wr_0_bits_data_0_0,
  input  [31:0]  io_tensor_wr_0_bits_data_0_1,
  input  [31:0]  io_tensor_wr_0_bits_data_0_2,
  input  [31:0]  io_tensor_wr_0_bits_data_0_3,
  input  [31:0]  io_tensor_wr_0_bits_data_0_4,
  input  [31:0]  io_tensor_wr_0_bits_data_0_5,
  input  [31:0]  io_tensor_wr_0_bits_data_0_6,
  input  [31:0]  io_tensor_wr_0_bits_data_0_7,
  input  [31:0]  io_tensor_wr_0_bits_data_0_8,
  input  [31:0]  io_tensor_wr_0_bits_data_0_9,
  input  [31:0]  io_tensor_wr_0_bits_data_0_10,
  input  [31:0]  io_tensor_wr_0_bits_data_0_11,
  input  [31:0]  io_tensor_wr_0_bits_data_0_12,
  input  [31:0]  io_tensor_wr_0_bits_data_0_13,
  input  [31:0]  io_tensor_wr_0_bits_data_0_14,
  input  [31:0]  io_tensor_wr_0_bits_data_0_15,
  input  [31:0]  io_tensor_wr_0_bits_data_0_16,
  input  [31:0]  io_tensor_wr_0_bits_data_0_17,
  input  [31:0]  io_tensor_wr_0_bits_data_0_18,
  input  [31:0]  io_tensor_wr_0_bits_data_0_19,
  input  [31:0]  io_tensor_wr_0_bits_data_0_20,
  input  [31:0]  io_tensor_wr_0_bits_data_0_21,
  input  [31:0]  io_tensor_wr_0_bits_data_0_22,
  input  [31:0]  io_tensor_wr_0_bits_data_0_23,
  input  [31:0]  io_tensor_wr_0_bits_data_0_24,
  input  [31:0]  io_tensor_wr_0_bits_data_0_25,
  input  [31:0]  io_tensor_wr_0_bits_data_0_26,
  input  [31:0]  io_tensor_wr_0_bits_data_0_27,
  input  [31:0]  io_tensor_wr_0_bits_data_0_28,
  input  [31:0]  io_tensor_wr_0_bits_data_0_29,
  input  [31:0]  io_tensor_wr_0_bits_data_0_30,
  input  [31:0]  io_tensor_wr_0_bits_data_0_31
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_27;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_33;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_39;
  reg [63:0] _RAND_42;
  reg [63:0] _RAND_45;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [63:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [127:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
`endif // RANDOMIZE_REG_INIT
  wire  vmeCmd_clock; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_reset; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_start; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_isBusy; // @[TensorLoadNarrowVME.scala 75:23]
  wire [127:0] vmeCmd_io_inst; // @[TensorLoadNarrowVME.scala 75:23]
  wire [31:0] vmeCmd_io_baddr; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_vmeCmd_ready; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_vmeCmd_valid; // @[TensorLoadNarrowVME.scala 75:23]
  wire [31:0] vmeCmd_io_vmeCmd_bits_addr; // @[TensorLoadNarrowVME.scala 75:23]
  wire [3:0] vmeCmd_io_vmeCmd_bits_len; // @[TensorLoadNarrowVME.scala 75:23]
  wire [20:0] vmeCmd_io_vmeCmd_bits_tag; // @[TensorLoadNarrowVME.scala 75:23]
  wire [4:0] vmeCmd_io_readLen; // @[TensorLoadNarrowVME.scala 75:23]
  wire  vmeCmd_io_done; // @[TensorLoadNarrowVME.scala 75:23]
  wire  readData_clock; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_reset; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_io_start; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_io_vmeData_ready; // @[TensorLoadNarrowVME.scala 105:24]
  wire  readData_io_vmeData_valid; // @[TensorLoadNarrowVME.scala 105:24]
  wire [20:0] readData_io_vmeData_bits_tag; // @[TensorLoadNarrowVME.scala 105:24]
  wire [6:0] readData_io_idx; // @[TensorLoadNarrowVME.scala 105:24]
  wire [3:0] readData_io_col; // @[TensorLoadNarrowVME.scala 105:24]
  wire  fillPadding_clock; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_reset; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_io_canWriteMem; // @[TensorLoadNarrowVME.scala 119:27]
  wire [127:0] fillPadding_io_inst; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_io_tensorIdx_valid; // @[TensorLoadNarrowVME.scala 119:27]
  wire [6:0] fillPadding_io_tensorIdx_bits; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_io_start; // @[TensorLoadNarrowVME.scala 119:27]
  wire  fillPadding_io_done; // @[TensorLoadNarrowVME.scala 119:27]
  reg [63:0] tensorFile_0 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_0_MPORT_16_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_0_MPORT_16_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_0_MPORT_16_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_0_MPORT_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_0_MPORT_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_0_MPORT_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_0_MPORT_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_0_MPORT_16_en_pipe_0;
  reg [6:0] tensorFile_0_MPORT_16_addr_pipe_0;
  reg [63:0] tensorFile_1 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_1_MPORT_17_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_1_MPORT_17_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_1_MPORT_17_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_1_MPORT_1_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_1_MPORT_1_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_1_MPORT_1_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_1_MPORT_1_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_1_MPORT_17_en_pipe_0;
  reg [6:0] tensorFile_1_MPORT_17_addr_pipe_0;
  reg [63:0] tensorFile_2 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_2_MPORT_18_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_2_MPORT_18_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_2_MPORT_18_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_2_MPORT_2_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_2_MPORT_2_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_2_MPORT_2_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_2_MPORT_2_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_2_MPORT_18_en_pipe_0;
  reg [6:0] tensorFile_2_MPORT_18_addr_pipe_0;
  reg [63:0] tensorFile_3 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_3_MPORT_19_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_3_MPORT_19_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_3_MPORT_19_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_3_MPORT_3_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_3_MPORT_3_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_3_MPORT_3_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_3_MPORT_3_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_3_MPORT_19_en_pipe_0;
  reg [6:0] tensorFile_3_MPORT_19_addr_pipe_0;
  reg [63:0] tensorFile_4 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_4_MPORT_20_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_4_MPORT_20_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_4_MPORT_20_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_4_MPORT_4_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_4_MPORT_4_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_4_MPORT_4_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_4_MPORT_4_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_4_MPORT_20_en_pipe_0;
  reg [6:0] tensorFile_4_MPORT_20_addr_pipe_0;
  reg [63:0] tensorFile_5 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_5_MPORT_21_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_5_MPORT_21_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_5_MPORT_21_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_5_MPORT_5_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_5_MPORT_5_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_5_MPORT_5_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_5_MPORT_5_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_5_MPORT_21_en_pipe_0;
  reg [6:0] tensorFile_5_MPORT_21_addr_pipe_0;
  reg [63:0] tensorFile_6 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_6_MPORT_22_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_6_MPORT_22_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_6_MPORT_22_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_6_MPORT_6_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_6_MPORT_6_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_6_MPORT_6_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_6_MPORT_6_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_6_MPORT_22_en_pipe_0;
  reg [6:0] tensorFile_6_MPORT_22_addr_pipe_0;
  reg [63:0] tensorFile_7 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_7_MPORT_23_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_7_MPORT_23_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_7_MPORT_23_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_7_MPORT_7_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_7_MPORT_7_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_7_MPORT_7_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_7_MPORT_7_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_7_MPORT_23_en_pipe_0;
  reg [6:0] tensorFile_7_MPORT_23_addr_pipe_0;
  reg [63:0] tensorFile_8 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_8_MPORT_24_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_8_MPORT_24_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_8_MPORT_24_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_8_MPORT_8_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_8_MPORT_8_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_8_MPORT_8_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_8_MPORT_8_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_8_MPORT_24_en_pipe_0;
  reg [6:0] tensorFile_8_MPORT_24_addr_pipe_0;
  reg [63:0] tensorFile_9 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_9_MPORT_25_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_9_MPORT_25_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_9_MPORT_25_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_9_MPORT_9_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_9_MPORT_9_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_9_MPORT_9_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_9_MPORT_9_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_9_MPORT_25_en_pipe_0;
  reg [6:0] tensorFile_9_MPORT_25_addr_pipe_0;
  reg [63:0] tensorFile_10 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_10_MPORT_26_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_10_MPORT_26_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_10_MPORT_26_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_10_MPORT_10_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_10_MPORT_10_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_10_MPORT_10_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_10_MPORT_10_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_10_MPORT_26_en_pipe_0;
  reg [6:0] tensorFile_10_MPORT_26_addr_pipe_0;
  reg [63:0] tensorFile_11 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_11_MPORT_27_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_11_MPORT_27_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_11_MPORT_27_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_11_MPORT_11_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_11_MPORT_11_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_11_MPORT_11_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_11_MPORT_11_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_11_MPORT_27_en_pipe_0;
  reg [6:0] tensorFile_11_MPORT_27_addr_pipe_0;
  reg [63:0] tensorFile_12 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_12_MPORT_28_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_12_MPORT_28_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_12_MPORT_28_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_12_MPORT_12_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_12_MPORT_12_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_12_MPORT_12_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_12_MPORT_12_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_12_MPORT_28_en_pipe_0;
  reg [6:0] tensorFile_12_MPORT_28_addr_pipe_0;
  reg [63:0] tensorFile_13 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_13_MPORT_29_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_13_MPORT_29_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_13_MPORT_29_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_13_MPORT_13_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_13_MPORT_13_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_13_MPORT_13_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_13_MPORT_13_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_13_MPORT_29_en_pipe_0;
  reg [6:0] tensorFile_13_MPORT_29_addr_pipe_0;
  reg [63:0] tensorFile_14 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_14_MPORT_30_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_14_MPORT_30_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_14_MPORT_30_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_14_MPORT_14_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_14_MPORT_14_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_14_MPORT_14_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_14_MPORT_14_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_14_MPORT_30_en_pipe_0;
  reg [6:0] tensorFile_14_MPORT_30_addr_pipe_0;
  reg [63:0] tensorFile_15 [0:127]; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_15_MPORT_31_en; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_15_MPORT_31_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_15_MPORT_31_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [63:0] tensorFile_15_MPORT_15_data; // @[TensorLoadNarrowVME.scala 152:16]
  wire [6:0] tensorFile_15_MPORT_15_addr; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_15_MPORT_15_mask; // @[TensorLoadNarrowVME.scala 152:16]
  wire  tensorFile_15_MPORT_15_en; // @[TensorLoadNarrowVME.scala 152:16]
  reg  tensorFile_15_MPORT_31_en_pipe_0;
  reg [6:0] tensorFile_15_MPORT_31_addr_pipe_0;
  reg  state; // @[TensorLoadNarrowVME.scala 54:22]
  reg [10:0] blocksInFlight; // @[TensorLoadNarrowVME.scala 87:27]
  wire  loadDone = blocksInFlight == 11'h0 & vmeCmd_io_done & state; // @[TensorLoadNarrowVME.scala 292:57]
  wire  localDone = loadDone & fillPadding_io_done; // @[TensorLoadNarrowVME.scala 293:25]
  wire  _GEN_0 = localDone ? 1'h0 : state; // @[TensorLoadNarrowVME.scala 61:25 62:11 54:22]
  wire  _GEN_1 = io_start | _GEN_0; // @[TensorLoadNarrowVME.scala 59:18 60:11]
  reg [63:0] vmeDataBitsPipe_data; // @[TensorLoadNarrowVME.scala 67:32]
  reg [20:0] vmeDataBitsPipe_tag; // @[TensorLoadNarrowVME.scala 67:32]
  reg  vmeDataValidPipe; // @[TensorLoadNarrowVME.scala 68:33]
  reg  vmeDataReadyPipe; // @[TensorLoadNarrowVME.scala 69:33]
  wire  vmeDataFirePipe = vmeDataValidPipe & vmeDataReadyPipe; // @[TensorLoadNarrowVME.scala 70:42]
  wire  _T = io_vme_rd_cmd_ready & io_vme_rd_cmd_valid; // @[Decoupled.scala 50:35]
  wire  _T_1 = state & _T; // @[TensorLoadNarrowVME.scala 90:21]
  wire  _T_3 = state & _T & ~vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 90:43]
  wire [10:0] _GEN_106 = {{6'd0}, vmeCmd_io_readLen}; // @[TensorLoadNarrowVME.scala 91:38]
  wire [10:0] _blocksInFlight_T_1 = blocksInFlight + _GEN_106; // @[TensorLoadNarrowVME.scala 91:38]
  wire  _T_6 = _T_1 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 92:43]
  wire [10:0] _blocksInFlight_T_5 = _blocksInFlight_T_1 - 11'h1; // @[TensorLoadNarrowVME.scala 93:48]
  wire  _T_10 = state & ~_T & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 94:44]
  wire  _T_13 = ~reset; // @[TensorLoadNarrowVME.scala 95:11]
  wire [10:0] _blocksInFlight_T_7 = blocksInFlight - 11'h1; // @[TensorLoadNarrowVME.scala 96:38]
  reg [127:0] fillPadding_io_inst_REG; // @[TensorLoadNarrowVME.scala 121:33]
  reg  fillPadding_io_start_REG; // @[TensorLoadNarrowVME.scala 122:34]
  wire [6:0] waddrTensInstrTmp = fillPadding_io_tensorIdx_valid ? fillPadding_io_tensorIdx_bits : readData_io_idx; // @[TensorLoadNarrowVME.scala 166:30]
  wire [55:0] waddrDirect_lo = {io_tensor_wr_0_bits_idx,io_tensor_wr_0_bits_idx,io_tensor_wr_0_bits_idx,
    io_tensor_wr_0_bits_idx,io_tensor_wr_0_bits_idx,io_tensor_wr_0_bits_idx,io_tensor_wr_0_bits_idx,
    io_tensor_wr_0_bits_idx}; // @[TensorLoadNarrowVME.scala 178:85]
  wire [111:0] _waddrDirect_T = {io_tensor_wr_0_bits_idx,io_tensor_wr_0_bits_idx,io_tensor_wr_0_bits_idx,
    io_tensor_wr_0_bits_idx,io_tensor_wr_0_bits_idx,io_tensor_wr_0_bits_idx,io_tensor_wr_0_bits_idx,
    io_tensor_wr_0_bits_idx,waddrDirect_lo}; // @[TensorLoadNarrowVME.scala 178:85]
  wire [6:0] waddrDirect_0 = _waddrDirect_T[6:0]; // @[TensorLoadNarrowVME.scala 178:85]
  wire [6:0] waddrDirect_1 = _waddrDirect_T[13:7]; // @[TensorLoadNarrowVME.scala 178:85]
  wire [6:0] waddrDirect_2 = _waddrDirect_T[20:14]; // @[TensorLoadNarrowVME.scala 178:85]
  wire [6:0] waddrDirect_3 = _waddrDirect_T[27:21]; // @[TensorLoadNarrowVME.scala 178:85]
  wire [6:0] waddrDirect_4 = _waddrDirect_T[34:28]; // @[TensorLoadNarrowVME.scala 178:85]
  wire [6:0] waddrDirect_5 = _waddrDirect_T[41:35]; // @[TensorLoadNarrowVME.scala 178:85]
  wire [6:0] waddrDirect_6 = _waddrDirect_T[48:42]; // @[TensorLoadNarrowVME.scala 178:85]
  wire [6:0] waddrDirect_7 = _waddrDirect_T[55:49]; // @[TensorLoadNarrowVME.scala 178:85]
  wire [6:0] waddrDirect_8 = _waddrDirect_T[62:56]; // @[TensorLoadNarrowVME.scala 178:85]
  wire [6:0] waddrDirect_9 = _waddrDirect_T[69:63]; // @[TensorLoadNarrowVME.scala 178:85]
  wire [6:0] waddrDirect_10 = _waddrDirect_T[76:70]; // @[TensorLoadNarrowVME.scala 178:85]
  wire [6:0] waddrDirect_11 = _waddrDirect_T[83:77]; // @[TensorLoadNarrowVME.scala 178:85]
  wire [6:0] waddrDirect_12 = _waddrDirect_T[90:84]; // @[TensorLoadNarrowVME.scala 178:85]
  wire [6:0] waddrDirect_13 = _waddrDirect_T[97:91]; // @[TensorLoadNarrowVME.scala 178:85]
  wire [6:0] waddrDirect_14 = _waddrDirect_T[104:98]; // @[TensorLoadNarrowVME.scala 178:85]
  wire [6:0] waddrDirect_15 = _waddrDirect_T[111:105]; // @[TensorLoadNarrowVME.scala 178:85]
  wire  _waddr_0_T = ~state; // @[TensorLoadNarrowVME.scala 186:27]
  wire  wenTensInstr_0 = fillPadding_io_tensorIdx_valid | readData_io_col == 4'h0 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_1 = fillPadding_io_tensorIdx_valid | readData_io_col == 4'h1 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_2 = fillPadding_io_tensorIdx_valid | readData_io_col == 4'h2 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_3 = fillPadding_io_tensorIdx_valid | readData_io_col == 4'h3 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_4 = fillPadding_io_tensorIdx_valid | readData_io_col == 4'h4 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_5 = fillPadding_io_tensorIdx_valid | readData_io_col == 4'h5 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_6 = fillPadding_io_tensorIdx_valid | readData_io_col == 4'h6 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_7 = fillPadding_io_tensorIdx_valid | readData_io_col == 4'h7 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_8 = fillPadding_io_tensorIdx_valid | readData_io_col == 4'h8 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_9 = fillPadding_io_tensorIdx_valid | readData_io_col == 4'h9 & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_10 = fillPadding_io_tensorIdx_valid | readData_io_col == 4'ha & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_11 = fillPadding_io_tensorIdx_valid | readData_io_col == 4'hb & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_12 = fillPadding_io_tensorIdx_valid | readData_io_col == 4'hc & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_13 = fillPadding_io_tensorIdx_valid | readData_io_col == 4'hd & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_14 = fillPadding_io_tensorIdx_valid | readData_io_col == 4'he & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire  wenTensInstr_15 = fillPadding_io_tensorIdx_valid | readData_io_col == 4'hf & vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 197:8]
  wire [63:0] wdataTensInstr_0 = fillPadding_io_tensorIdx_valid ? 64'h0 : vmeDataBitsPipe_data; // @[TensorLoadNarrowVME.scala 234:29]
  wire [255:0] wdataDirect_lo_lo = {io_tensor_wr_0_bits_data_0_7,io_tensor_wr_0_bits_data_0_6,
    io_tensor_wr_0_bits_data_0_5,io_tensor_wr_0_bits_data_0_4,io_tensor_wr_0_bits_data_0_3,io_tensor_wr_0_bits_data_0_2,
    io_tensor_wr_0_bits_data_0_1,io_tensor_wr_0_bits_data_0_0}; // @[TensorLoadNarrowVME.scala 247:18]
  wire [511:0] wdataDirect_lo = {io_tensor_wr_0_bits_data_0_15,io_tensor_wr_0_bits_data_0_14,
    io_tensor_wr_0_bits_data_0_13,io_tensor_wr_0_bits_data_0_12,io_tensor_wr_0_bits_data_0_11,
    io_tensor_wr_0_bits_data_0_10,io_tensor_wr_0_bits_data_0_9,io_tensor_wr_0_bits_data_0_8,wdataDirect_lo_lo}; // @[TensorLoadNarrowVME.scala 247:18]
  wire [255:0] wdataDirect_hi_lo = {io_tensor_wr_0_bits_data_0_23,io_tensor_wr_0_bits_data_0_22,
    io_tensor_wr_0_bits_data_0_21,io_tensor_wr_0_bits_data_0_20,io_tensor_wr_0_bits_data_0_19,
    io_tensor_wr_0_bits_data_0_18,io_tensor_wr_0_bits_data_0_17,io_tensor_wr_0_bits_data_0_16}; // @[TensorLoadNarrowVME.scala 247:18]
  wire [1023:0] _wdataDirect_T = {io_tensor_wr_0_bits_data_0_31,io_tensor_wr_0_bits_data_0_30,
    io_tensor_wr_0_bits_data_0_29,io_tensor_wr_0_bits_data_0_28,io_tensor_wr_0_bits_data_0_27,
    io_tensor_wr_0_bits_data_0_26,io_tensor_wr_0_bits_data_0_25,io_tensor_wr_0_bits_data_0_24,wdataDirect_hi_lo,
    wdataDirect_lo}; // @[TensorLoadNarrowVME.scala 247:18]
  wire [63:0] wdataDirect_0 = _wdataDirect_T[63:0]; // @[TensorLoadNarrowVME.scala 247:18]
  reg  rvalid; // @[Reg.scala 28:20]
  wire [63:0] _WIRE_16_1 = tensorFile_1_MPORT_17_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_16_0 = tensorFile_0_MPORT_16_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_16_3 = tensorFile_3_MPORT_19_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_16_2 = tensorFile_2_MPORT_18_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_16_5 = tensorFile_5_MPORT_21_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_16_4 = tensorFile_4_MPORT_20_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_16_7 = tensorFile_7_MPORT_23_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_16_6 = tensorFile_6_MPORT_22_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [511:0] lo = {_WIRE_16_7,_WIRE_16_6,_WIRE_16_5,_WIRE_16_4,_WIRE_16_3,_WIRE_16_2,_WIRE_16_1,_WIRE_16_0}; // @[TensorLoadNarrowVME.scala 288:18]
  wire [63:0] _WIRE_16_9 = tensorFile_9_MPORT_25_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_16_8 = tensorFile_8_MPORT_24_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_16_11 = tensorFile_11_MPORT_27_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_16_10 = tensorFile_10_MPORT_26_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_16_13 = tensorFile_13_MPORT_29_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_16_12 = tensorFile_12_MPORT_28_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_16_15 = tensorFile_15_MPORT_31_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [63:0] _WIRE_16_14 = tensorFile_14_MPORT_30_data; // @[TensorLoadNarrowVME.scala 284:{14,14}]
  wire [1023:0] _T_52 = {_WIRE_16_15,_WIRE_16_14,_WIRE_16_13,_WIRE_16_12,_WIRE_16_11,_WIRE_16_10,_WIRE_16_9,_WIRE_16_8,
    lo}; // @[TensorLoadNarrowVME.scala 288:18]
  GenVMECmd_2 vmeCmd ( // @[TensorLoadNarrowVME.scala 75:23]
    .clock(vmeCmd_clock),
    .reset(vmeCmd_reset),
    .io_start(vmeCmd_io_start),
    .io_isBusy(vmeCmd_io_isBusy),
    .io_inst(vmeCmd_io_inst),
    .io_baddr(vmeCmd_io_baddr),
    .io_vmeCmd_ready(vmeCmd_io_vmeCmd_ready),
    .io_vmeCmd_valid(vmeCmd_io_vmeCmd_valid),
    .io_vmeCmd_bits_addr(vmeCmd_io_vmeCmd_bits_addr),
    .io_vmeCmd_bits_len(vmeCmd_io_vmeCmd_bits_len),
    .io_vmeCmd_bits_tag(vmeCmd_io_vmeCmd_bits_tag),
    .io_readLen(vmeCmd_io_readLen),
    .io_done(vmeCmd_io_done)
  );
  ReadVMEData_2 readData ( // @[TensorLoadNarrowVME.scala 105:24]
    .clock(readData_clock),
    .reset(readData_reset),
    .io_start(readData_io_start),
    .io_vmeData_ready(readData_io_vmeData_ready),
    .io_vmeData_valid(readData_io_vmeData_valid),
    .io_vmeData_bits_tag(readData_io_vmeData_bits_tag),
    .io_idx(readData_io_idx),
    .io_col(readData_io_col)
  );
  ZeroPadding fillPadding ( // @[TensorLoadNarrowVME.scala 119:27]
    .clock(fillPadding_clock),
    .reset(fillPadding_reset),
    .io_canWriteMem(fillPadding_io_canWriteMem),
    .io_inst(fillPadding_io_inst),
    .io_tensorIdx_valid(fillPadding_io_tensorIdx_valid),
    .io_tensorIdx_bits(fillPadding_io_tensorIdx_bits),
    .io_start(fillPadding_io_start),
    .io_done(fillPadding_io_done)
  );
  assign tensorFile_0_MPORT_16_en = tensorFile_0_MPORT_16_en_pipe_0;
  assign tensorFile_0_MPORT_16_addr = tensorFile_0_MPORT_16_addr_pipe_0;
  assign tensorFile_0_MPORT_16_data = tensorFile_0[tensorFile_0_MPORT_16_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_0_MPORT_data = _waddr_0_T ? wdataDirect_0 : wdataTensInstr_0;
  assign tensorFile_0_MPORT_addr = _waddr_0_T ? waddrDirect_0 : waddrTensInstrTmp;
  assign tensorFile_0_MPORT_mask = 1'h1;
  assign tensorFile_0_MPORT_en = _waddr_0_T ? io_tensor_wr_0_valid : wenTensInstr_0;
  assign tensorFile_1_MPORT_17_en = tensorFile_1_MPORT_17_en_pipe_0;
  assign tensorFile_1_MPORT_17_addr = tensorFile_1_MPORT_17_addr_pipe_0;
  assign tensorFile_1_MPORT_17_data = tensorFile_1[tensorFile_1_MPORT_17_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_1_MPORT_1_data = _waddr_0_T ? _wdataDirect_T[127:64] : wdataTensInstr_0;
  assign tensorFile_1_MPORT_1_addr = _waddr_0_T ? waddrDirect_1 : waddrTensInstrTmp;
  assign tensorFile_1_MPORT_1_mask = 1'h1;
  assign tensorFile_1_MPORT_1_en = _waddr_0_T ? io_tensor_wr_0_valid : wenTensInstr_1;
  assign tensorFile_2_MPORT_18_en = tensorFile_2_MPORT_18_en_pipe_0;
  assign tensorFile_2_MPORT_18_addr = tensorFile_2_MPORT_18_addr_pipe_0;
  assign tensorFile_2_MPORT_18_data = tensorFile_2[tensorFile_2_MPORT_18_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_2_MPORT_2_data = _waddr_0_T ? _wdataDirect_T[191:128] : wdataTensInstr_0;
  assign tensorFile_2_MPORT_2_addr = _waddr_0_T ? waddrDirect_2 : waddrTensInstrTmp;
  assign tensorFile_2_MPORT_2_mask = 1'h1;
  assign tensorFile_2_MPORT_2_en = _waddr_0_T ? io_tensor_wr_0_valid : wenTensInstr_2;
  assign tensorFile_3_MPORT_19_en = tensorFile_3_MPORT_19_en_pipe_0;
  assign tensorFile_3_MPORT_19_addr = tensorFile_3_MPORT_19_addr_pipe_0;
  assign tensorFile_3_MPORT_19_data = tensorFile_3[tensorFile_3_MPORT_19_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_3_MPORT_3_data = _waddr_0_T ? _wdataDirect_T[255:192] : wdataTensInstr_0;
  assign tensorFile_3_MPORT_3_addr = _waddr_0_T ? waddrDirect_3 : waddrTensInstrTmp;
  assign tensorFile_3_MPORT_3_mask = 1'h1;
  assign tensorFile_3_MPORT_3_en = _waddr_0_T ? io_tensor_wr_0_valid : wenTensInstr_3;
  assign tensorFile_4_MPORT_20_en = tensorFile_4_MPORT_20_en_pipe_0;
  assign tensorFile_4_MPORT_20_addr = tensorFile_4_MPORT_20_addr_pipe_0;
  assign tensorFile_4_MPORT_20_data = tensorFile_4[tensorFile_4_MPORT_20_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_4_MPORT_4_data = _waddr_0_T ? _wdataDirect_T[319:256] : wdataTensInstr_0;
  assign tensorFile_4_MPORT_4_addr = _waddr_0_T ? waddrDirect_4 : waddrTensInstrTmp;
  assign tensorFile_4_MPORT_4_mask = 1'h1;
  assign tensorFile_4_MPORT_4_en = _waddr_0_T ? io_tensor_wr_0_valid : wenTensInstr_4;
  assign tensorFile_5_MPORT_21_en = tensorFile_5_MPORT_21_en_pipe_0;
  assign tensorFile_5_MPORT_21_addr = tensorFile_5_MPORT_21_addr_pipe_0;
  assign tensorFile_5_MPORT_21_data = tensorFile_5[tensorFile_5_MPORT_21_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_5_MPORT_5_data = _waddr_0_T ? _wdataDirect_T[383:320] : wdataTensInstr_0;
  assign tensorFile_5_MPORT_5_addr = _waddr_0_T ? waddrDirect_5 : waddrTensInstrTmp;
  assign tensorFile_5_MPORT_5_mask = 1'h1;
  assign tensorFile_5_MPORT_5_en = _waddr_0_T ? io_tensor_wr_0_valid : wenTensInstr_5;
  assign tensorFile_6_MPORT_22_en = tensorFile_6_MPORT_22_en_pipe_0;
  assign tensorFile_6_MPORT_22_addr = tensorFile_6_MPORT_22_addr_pipe_0;
  assign tensorFile_6_MPORT_22_data = tensorFile_6[tensorFile_6_MPORT_22_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_6_MPORT_6_data = _waddr_0_T ? _wdataDirect_T[447:384] : wdataTensInstr_0;
  assign tensorFile_6_MPORT_6_addr = _waddr_0_T ? waddrDirect_6 : waddrTensInstrTmp;
  assign tensorFile_6_MPORT_6_mask = 1'h1;
  assign tensorFile_6_MPORT_6_en = _waddr_0_T ? io_tensor_wr_0_valid : wenTensInstr_6;
  assign tensorFile_7_MPORT_23_en = tensorFile_7_MPORT_23_en_pipe_0;
  assign tensorFile_7_MPORT_23_addr = tensorFile_7_MPORT_23_addr_pipe_0;
  assign tensorFile_7_MPORT_23_data = tensorFile_7[tensorFile_7_MPORT_23_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_7_MPORT_7_data = _waddr_0_T ? _wdataDirect_T[511:448] : wdataTensInstr_0;
  assign tensorFile_7_MPORT_7_addr = _waddr_0_T ? waddrDirect_7 : waddrTensInstrTmp;
  assign tensorFile_7_MPORT_7_mask = 1'h1;
  assign tensorFile_7_MPORT_7_en = _waddr_0_T ? io_tensor_wr_0_valid : wenTensInstr_7;
  assign tensorFile_8_MPORT_24_en = tensorFile_8_MPORT_24_en_pipe_0;
  assign tensorFile_8_MPORT_24_addr = tensorFile_8_MPORT_24_addr_pipe_0;
  assign tensorFile_8_MPORT_24_data = tensorFile_8[tensorFile_8_MPORT_24_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_8_MPORT_8_data = _waddr_0_T ? _wdataDirect_T[575:512] : wdataTensInstr_0;
  assign tensorFile_8_MPORT_8_addr = _waddr_0_T ? waddrDirect_8 : waddrTensInstrTmp;
  assign tensorFile_8_MPORT_8_mask = 1'h1;
  assign tensorFile_8_MPORT_8_en = _waddr_0_T ? io_tensor_wr_0_valid : wenTensInstr_8;
  assign tensorFile_9_MPORT_25_en = tensorFile_9_MPORT_25_en_pipe_0;
  assign tensorFile_9_MPORT_25_addr = tensorFile_9_MPORT_25_addr_pipe_0;
  assign tensorFile_9_MPORT_25_data = tensorFile_9[tensorFile_9_MPORT_25_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_9_MPORT_9_data = _waddr_0_T ? _wdataDirect_T[639:576] : wdataTensInstr_0;
  assign tensorFile_9_MPORT_9_addr = _waddr_0_T ? waddrDirect_9 : waddrTensInstrTmp;
  assign tensorFile_9_MPORT_9_mask = 1'h1;
  assign tensorFile_9_MPORT_9_en = _waddr_0_T ? io_tensor_wr_0_valid : wenTensInstr_9;
  assign tensorFile_10_MPORT_26_en = tensorFile_10_MPORT_26_en_pipe_0;
  assign tensorFile_10_MPORT_26_addr = tensorFile_10_MPORT_26_addr_pipe_0;
  assign tensorFile_10_MPORT_26_data = tensorFile_10[tensorFile_10_MPORT_26_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_10_MPORT_10_data = _waddr_0_T ? _wdataDirect_T[703:640] : wdataTensInstr_0;
  assign tensorFile_10_MPORT_10_addr = _waddr_0_T ? waddrDirect_10 : waddrTensInstrTmp;
  assign tensorFile_10_MPORT_10_mask = 1'h1;
  assign tensorFile_10_MPORT_10_en = _waddr_0_T ? io_tensor_wr_0_valid : wenTensInstr_10;
  assign tensorFile_11_MPORT_27_en = tensorFile_11_MPORT_27_en_pipe_0;
  assign tensorFile_11_MPORT_27_addr = tensorFile_11_MPORT_27_addr_pipe_0;
  assign tensorFile_11_MPORT_27_data = tensorFile_11[tensorFile_11_MPORT_27_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_11_MPORT_11_data = _waddr_0_T ? _wdataDirect_T[767:704] : wdataTensInstr_0;
  assign tensorFile_11_MPORT_11_addr = _waddr_0_T ? waddrDirect_11 : waddrTensInstrTmp;
  assign tensorFile_11_MPORT_11_mask = 1'h1;
  assign tensorFile_11_MPORT_11_en = _waddr_0_T ? io_tensor_wr_0_valid : wenTensInstr_11;
  assign tensorFile_12_MPORT_28_en = tensorFile_12_MPORT_28_en_pipe_0;
  assign tensorFile_12_MPORT_28_addr = tensorFile_12_MPORT_28_addr_pipe_0;
  assign tensorFile_12_MPORT_28_data = tensorFile_12[tensorFile_12_MPORT_28_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_12_MPORT_12_data = _waddr_0_T ? _wdataDirect_T[831:768] : wdataTensInstr_0;
  assign tensorFile_12_MPORT_12_addr = _waddr_0_T ? waddrDirect_12 : waddrTensInstrTmp;
  assign tensorFile_12_MPORT_12_mask = 1'h1;
  assign tensorFile_12_MPORT_12_en = _waddr_0_T ? io_tensor_wr_0_valid : wenTensInstr_12;
  assign tensorFile_13_MPORT_29_en = tensorFile_13_MPORT_29_en_pipe_0;
  assign tensorFile_13_MPORT_29_addr = tensorFile_13_MPORT_29_addr_pipe_0;
  assign tensorFile_13_MPORT_29_data = tensorFile_13[tensorFile_13_MPORT_29_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_13_MPORT_13_data = _waddr_0_T ? _wdataDirect_T[895:832] : wdataTensInstr_0;
  assign tensorFile_13_MPORT_13_addr = _waddr_0_T ? waddrDirect_13 : waddrTensInstrTmp;
  assign tensorFile_13_MPORT_13_mask = 1'h1;
  assign tensorFile_13_MPORT_13_en = _waddr_0_T ? io_tensor_wr_0_valid : wenTensInstr_13;
  assign tensorFile_14_MPORT_30_en = tensorFile_14_MPORT_30_en_pipe_0;
  assign tensorFile_14_MPORT_30_addr = tensorFile_14_MPORT_30_addr_pipe_0;
  assign tensorFile_14_MPORT_30_data = tensorFile_14[tensorFile_14_MPORT_30_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_14_MPORT_14_data = _waddr_0_T ? _wdataDirect_T[959:896] : wdataTensInstr_0;
  assign tensorFile_14_MPORT_14_addr = _waddr_0_T ? waddrDirect_14 : waddrTensInstrTmp;
  assign tensorFile_14_MPORT_14_mask = 1'h1;
  assign tensorFile_14_MPORT_14_en = _waddr_0_T ? io_tensor_wr_0_valid : wenTensInstr_14;
  assign tensorFile_15_MPORT_31_en = tensorFile_15_MPORT_31_en_pipe_0;
  assign tensorFile_15_MPORT_31_addr = tensorFile_15_MPORT_31_addr_pipe_0;
  assign tensorFile_15_MPORT_31_data = tensorFile_15[tensorFile_15_MPORT_31_addr]; // @[TensorLoadNarrowVME.scala 152:16]
  assign tensorFile_15_MPORT_15_data = _waddr_0_T ? _wdataDirect_T[1023:960] : wdataTensInstr_0;
  assign tensorFile_15_MPORT_15_addr = _waddr_0_T ? waddrDirect_15 : waddrTensInstrTmp;
  assign tensorFile_15_MPORT_15_mask = 1'h1;
  assign tensorFile_15_MPORT_15_en = _waddr_0_T ? io_tensor_wr_0_valid : wenTensInstr_15;
  assign io_done = loadDone & fillPadding_io_done; // @[TensorLoadNarrowVME.scala 293:25]
  assign io_vme_rd_cmd_valid = vmeCmd_io_vmeCmd_valid; // @[TensorLoadNarrowVME.scala 80:20]
  assign io_vme_rd_cmd_bits_addr = vmeCmd_io_vmeCmd_bits_addr; // @[TensorLoadNarrowVME.scala 80:20]
  assign io_vme_rd_cmd_bits_len = vmeCmd_io_vmeCmd_bits_len; // @[TensorLoadNarrowVME.scala 80:20]
  assign io_vme_rd_cmd_bits_tag = vmeCmd_io_vmeCmd_bits_tag; // @[TensorLoadNarrowVME.scala 80:20]
  assign io_vme_rd_data_ready = 1'h1; // @[TensorLoadNarrowVME.scala 111:24]
  assign io_tensor_rd_0_data_valid = rvalid; // @[TensorLoadNarrowVME.scala 278:36]
  assign io_tensor_rd_0_data_bits_0_0 = _T_52[31:0]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_1 = _T_52[63:32]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_2 = _T_52[95:64]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_3 = _T_52[127:96]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_4 = _T_52[159:128]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_5 = _T_52[191:160]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_6 = _T_52[223:192]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_7 = _T_52[255:224]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_8 = _T_52[287:256]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_9 = _T_52[319:288]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_10 = _T_52[351:320]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_11 = _T_52[383:352]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_12 = _T_52[415:384]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_13 = _T_52[447:416]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_14 = _T_52[479:448]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_15 = _T_52[511:480]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_16 = _T_52[543:512]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_17 = _T_52[575:544]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_18 = _T_52[607:576]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_19 = _T_52[639:608]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_20 = _T_52[671:640]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_21 = _T_52[703:672]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_22 = _T_52[735:704]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_23 = _T_52[767:736]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_24 = _T_52[799:768]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_25 = _T_52[831:800]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_26 = _T_52[863:832]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_27 = _T_52[895:864]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_28 = _T_52[927:896]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_29 = _T_52[959:928]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_30 = _T_52[991:960]; // @[TensorLoadNarrowVME.scala 288:18]
  assign io_tensor_rd_0_data_bits_0_31 = _T_52[1023:992]; // @[TensorLoadNarrowVME.scala 288:18]
  assign vmeCmd_clock = clock;
  assign vmeCmd_reset = reset;
  assign vmeCmd_io_start = io_start; // @[TensorLoadNarrowVME.scala 76:19]
  assign vmeCmd_io_isBusy = state; // @[TensorLoadNarrowVME.scala 56:22]
  assign vmeCmd_io_inst = io_inst; // @[TensorLoadNarrowVME.scala 78:18]
  assign vmeCmd_io_baddr = io_baddr; // @[TensorLoadNarrowVME.scala 79:19]
  assign vmeCmd_io_vmeCmd_ready = io_vme_rd_cmd_ready; // @[TensorLoadNarrowVME.scala 80:20]
  assign readData_clock = clock;
  assign readData_reset = reset;
  assign readData_io_start = io_start; // @[TensorLoadNarrowVME.scala 106:21]
  assign readData_io_vmeData_valid = vmeDataValidPipe; // @[TensorLoadNarrowVME.scala 107:29]
  assign readData_io_vmeData_bits_tag = vmeDataBitsPipe_tag; // @[TensorLoadNarrowVME.scala 108:28]
  assign fillPadding_clock = clock;
  assign fillPadding_reset = reset;
  assign fillPadding_io_canWriteMem = ~vmeDataFirePipe; // @[TensorLoadNarrowVME.scala 120:33]
  assign fillPadding_io_inst = fillPadding_io_inst_REG; // @[TensorLoadNarrowVME.scala 121:23]
  assign fillPadding_io_start = fillPadding_io_start_REG; // @[TensorLoadNarrowVME.scala 122:24]
  always @(posedge clock) begin
    if (tensorFile_0_MPORT_en & tensorFile_0_MPORT_mask) begin
      tensorFile_0[tensorFile_0_MPORT_addr] <= tensorFile_0_MPORT_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_0_MPORT_16_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_0_MPORT_16_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_1_MPORT_1_en & tensorFile_1_MPORT_1_mask) begin
      tensorFile_1[tensorFile_1_MPORT_1_addr] <= tensorFile_1_MPORT_1_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_1_MPORT_17_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_1_MPORT_17_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_2_MPORT_2_en & tensorFile_2_MPORT_2_mask) begin
      tensorFile_2[tensorFile_2_MPORT_2_addr] <= tensorFile_2_MPORT_2_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_2_MPORT_18_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_2_MPORT_18_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_3_MPORT_3_en & tensorFile_3_MPORT_3_mask) begin
      tensorFile_3[tensorFile_3_MPORT_3_addr] <= tensorFile_3_MPORT_3_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_3_MPORT_19_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_3_MPORT_19_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_4_MPORT_4_en & tensorFile_4_MPORT_4_mask) begin
      tensorFile_4[tensorFile_4_MPORT_4_addr] <= tensorFile_4_MPORT_4_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_4_MPORT_20_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_4_MPORT_20_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_5_MPORT_5_en & tensorFile_5_MPORT_5_mask) begin
      tensorFile_5[tensorFile_5_MPORT_5_addr] <= tensorFile_5_MPORT_5_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_5_MPORT_21_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_5_MPORT_21_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_6_MPORT_6_en & tensorFile_6_MPORT_6_mask) begin
      tensorFile_6[tensorFile_6_MPORT_6_addr] <= tensorFile_6_MPORT_6_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_6_MPORT_22_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_6_MPORT_22_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_7_MPORT_7_en & tensorFile_7_MPORT_7_mask) begin
      tensorFile_7[tensorFile_7_MPORT_7_addr] <= tensorFile_7_MPORT_7_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_7_MPORT_23_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_7_MPORT_23_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_8_MPORT_8_en & tensorFile_8_MPORT_8_mask) begin
      tensorFile_8[tensorFile_8_MPORT_8_addr] <= tensorFile_8_MPORT_8_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_8_MPORT_24_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_8_MPORT_24_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_9_MPORT_9_en & tensorFile_9_MPORT_9_mask) begin
      tensorFile_9[tensorFile_9_MPORT_9_addr] <= tensorFile_9_MPORT_9_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_9_MPORT_25_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_9_MPORT_25_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_10_MPORT_10_en & tensorFile_10_MPORT_10_mask) begin
      tensorFile_10[tensorFile_10_MPORT_10_addr] <= tensorFile_10_MPORT_10_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_10_MPORT_26_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_10_MPORT_26_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_11_MPORT_11_en & tensorFile_11_MPORT_11_mask) begin
      tensorFile_11[tensorFile_11_MPORT_11_addr] <= tensorFile_11_MPORT_11_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_11_MPORT_27_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_11_MPORT_27_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_12_MPORT_12_en & tensorFile_12_MPORT_12_mask) begin
      tensorFile_12[tensorFile_12_MPORT_12_addr] <= tensorFile_12_MPORT_12_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_12_MPORT_28_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_12_MPORT_28_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_13_MPORT_13_en & tensorFile_13_MPORT_13_mask) begin
      tensorFile_13[tensorFile_13_MPORT_13_addr] <= tensorFile_13_MPORT_13_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_13_MPORT_29_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_13_MPORT_29_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_14_MPORT_14_en & tensorFile_14_MPORT_14_mask) begin
      tensorFile_14[tensorFile_14_MPORT_14_addr] <= tensorFile_14_MPORT_14_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_14_MPORT_30_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_14_MPORT_30_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (tensorFile_15_MPORT_15_en & tensorFile_15_MPORT_15_mask) begin
      tensorFile_15[tensorFile_15_MPORT_15_addr] <= tensorFile_15_MPORT_15_data; // @[TensorLoadNarrowVME.scala 152:16]
    end
    tensorFile_15_MPORT_31_en_pipe_0 <= io_tensor_rd_0_idx_valid;
    if (io_tensor_rd_0_idx_valid) begin
      tensorFile_15_MPORT_31_addr_pipe_0 <= io_tensor_rd_0_idx_bits;
    end
    if (reset) begin // @[TensorLoadNarrowVME.scala 54:22]
      state <= 1'h0; // @[TensorLoadNarrowVME.scala 54:22]
    end else begin
      state <= _GEN_1;
    end
    if (io_start) begin // @[TensorLoadNarrowVME.scala 88:18]
      blocksInFlight <= 11'h0; // @[TensorLoadNarrowVME.scala 89:20]
    end else if (state & _T & ~vmeDataFirePipe) begin // @[TensorLoadNarrowVME.scala 90:64]
      blocksInFlight <= _blocksInFlight_T_1; // @[TensorLoadNarrowVME.scala 91:20]
    end else if (_T_1 & vmeDataFirePipe) begin // @[TensorLoadNarrowVME.scala 92:63]
      blocksInFlight <= _blocksInFlight_T_5; // @[TensorLoadNarrowVME.scala 93:20]
    end else if (state & ~_T & vmeDataFirePipe) begin // @[TensorLoadNarrowVME.scala 94:64]
      blocksInFlight <= _blocksInFlight_T_7; // @[TensorLoadNarrowVME.scala 96:20]
    end
    vmeDataBitsPipe_data <= io_vme_rd_data_bits_data; // @[TensorLoadNarrowVME.scala 67:32]
    vmeDataBitsPipe_tag <= io_vme_rd_data_bits_tag; // @[TensorLoadNarrowVME.scala 67:32]
    if (reset) begin // @[TensorLoadNarrowVME.scala 68:33]
      vmeDataValidPipe <= 1'h0; // @[TensorLoadNarrowVME.scala 68:33]
    end else begin
      vmeDataValidPipe <= io_vme_rd_data_valid; // @[TensorLoadNarrowVME.scala 68:33]
    end
    if (reset) begin // @[TensorLoadNarrowVME.scala 69:33]
      vmeDataReadyPipe <= 1'h0; // @[TensorLoadNarrowVME.scala 69:33]
    end else begin
      vmeDataReadyPipe <= io_vme_rd_data_ready; // @[TensorLoadNarrowVME.scala 69:33]
    end
    fillPadding_io_inst_REG <= io_inst; // @[TensorLoadNarrowVME.scala 121:33]
    if (reset) begin // @[TensorLoadNarrowVME.scala 122:34]
      fillPadding_io_start_REG <= 1'h0; // @[TensorLoadNarrowVME.scala 122:34]
    end else begin
      fillPadding_io_start_REG <= io_start; // @[TensorLoadNarrowVME.scala 122:34]
    end
    if (reset) begin // @[Reg.scala 28:20]
      rvalid <= 1'h0; // @[Reg.scala 28:20]
    end else begin
      rvalid <= io_tensor_rd_0_idx_valid;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~io_start & ~_T_3 & ~_T_6 & _T_10 & ~reset & ~(blocksInFlight > 11'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TensorLoadNarrowVME.scala:95 assert(blocksInFlight > 0.U)\n"); // @[TensorLoadNarrowVME.scala 95:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_0[initvar] = _RAND_0[63:0];
  _RAND_3 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_1[initvar] = _RAND_3[63:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_2[initvar] = _RAND_6[63:0];
  _RAND_9 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_3[initvar] = _RAND_9[63:0];
  _RAND_12 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_4[initvar] = _RAND_12[63:0];
  _RAND_15 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_5[initvar] = _RAND_15[63:0];
  _RAND_18 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_6[initvar] = _RAND_18[63:0];
  _RAND_21 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_7[initvar] = _RAND_21[63:0];
  _RAND_24 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_8[initvar] = _RAND_24[63:0];
  _RAND_27 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_9[initvar] = _RAND_27[63:0];
  _RAND_30 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_10[initvar] = _RAND_30[63:0];
  _RAND_33 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_11[initvar] = _RAND_33[63:0];
  _RAND_36 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_12[initvar] = _RAND_36[63:0];
  _RAND_39 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_13[initvar] = _RAND_39[63:0];
  _RAND_42 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_14[initvar] = _RAND_42[63:0];
  _RAND_45 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_15[initvar] = _RAND_45[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tensorFile_0_MPORT_16_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  tensorFile_0_MPORT_16_addr_pipe_0 = _RAND_2[6:0];
  _RAND_4 = {1{`RANDOM}};
  tensorFile_1_MPORT_17_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  tensorFile_1_MPORT_17_addr_pipe_0 = _RAND_5[6:0];
  _RAND_7 = {1{`RANDOM}};
  tensorFile_2_MPORT_18_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  tensorFile_2_MPORT_18_addr_pipe_0 = _RAND_8[6:0];
  _RAND_10 = {1{`RANDOM}};
  tensorFile_3_MPORT_19_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  tensorFile_3_MPORT_19_addr_pipe_0 = _RAND_11[6:0];
  _RAND_13 = {1{`RANDOM}};
  tensorFile_4_MPORT_20_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  tensorFile_4_MPORT_20_addr_pipe_0 = _RAND_14[6:0];
  _RAND_16 = {1{`RANDOM}};
  tensorFile_5_MPORT_21_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  tensorFile_5_MPORT_21_addr_pipe_0 = _RAND_17[6:0];
  _RAND_19 = {1{`RANDOM}};
  tensorFile_6_MPORT_22_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  tensorFile_6_MPORT_22_addr_pipe_0 = _RAND_20[6:0];
  _RAND_22 = {1{`RANDOM}};
  tensorFile_7_MPORT_23_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  tensorFile_7_MPORT_23_addr_pipe_0 = _RAND_23[6:0];
  _RAND_25 = {1{`RANDOM}};
  tensorFile_8_MPORT_24_en_pipe_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  tensorFile_8_MPORT_24_addr_pipe_0 = _RAND_26[6:0];
  _RAND_28 = {1{`RANDOM}};
  tensorFile_9_MPORT_25_en_pipe_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  tensorFile_9_MPORT_25_addr_pipe_0 = _RAND_29[6:0];
  _RAND_31 = {1{`RANDOM}};
  tensorFile_10_MPORT_26_en_pipe_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  tensorFile_10_MPORT_26_addr_pipe_0 = _RAND_32[6:0];
  _RAND_34 = {1{`RANDOM}};
  tensorFile_11_MPORT_27_en_pipe_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  tensorFile_11_MPORT_27_addr_pipe_0 = _RAND_35[6:0];
  _RAND_37 = {1{`RANDOM}};
  tensorFile_12_MPORT_28_en_pipe_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  tensorFile_12_MPORT_28_addr_pipe_0 = _RAND_38[6:0];
  _RAND_40 = {1{`RANDOM}};
  tensorFile_13_MPORT_29_en_pipe_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  tensorFile_13_MPORT_29_addr_pipe_0 = _RAND_41[6:0];
  _RAND_43 = {1{`RANDOM}};
  tensorFile_14_MPORT_30_en_pipe_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  tensorFile_14_MPORT_30_addr_pipe_0 = _RAND_44[6:0];
  _RAND_46 = {1{`RANDOM}};
  tensorFile_15_MPORT_31_en_pipe_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  tensorFile_15_MPORT_31_addr_pipe_0 = _RAND_47[6:0];
  _RAND_48 = {1{`RANDOM}};
  state = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  blocksInFlight = _RAND_49[10:0];
  _RAND_50 = {2{`RANDOM}};
  vmeDataBitsPipe_data = _RAND_50[63:0];
  _RAND_51 = {1{`RANDOM}};
  vmeDataBitsPipe_tag = _RAND_51[20:0];
  _RAND_52 = {1{`RANDOM}};
  vmeDataValidPipe = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  vmeDataReadyPipe = _RAND_53[0:0];
  _RAND_54 = {4{`RANDOM}};
  fillPadding_io_inst_REG = _RAND_54[127:0];
  _RAND_55 = {1{`RANDOM}};
  fillPadding_io_start_REG = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  rvalid = _RAND_56[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~io_start & ~_T_3 & ~_T_6 & _T_10 & ~reset) begin
      assert(blocksInFlight > 11'h0); // @[TensorLoadNarrowVME.scala 95:11]
    end
    //
    if (_T_13) begin
      assert(1'h1); // @[TensorLoadNarrowVME.scala 109:9]
    end
  end
endmodule
module TensorLoadAcc(
  input          clock,
  input          reset,
  input          io_start,
  output         io_done,
  input  [127:0] io_inst,
  input  [31:0]  io_baddr,
  input          io_vme_rd_cmd_ready,
  output         io_vme_rd_cmd_valid,
  output [31:0]  io_vme_rd_cmd_bits_addr,
  output [3:0]   io_vme_rd_cmd_bits_len,
  output [20:0]  io_vme_rd_cmd_bits_tag,
  input          io_vme_rd_data_valid,
  input  [63:0]  io_vme_rd_data_bits_data,
  input  [20:0]  io_vme_rd_data_bits_tag,
  input          io_tensor_rd_0_idx_valid,
  input  [6:0]   io_tensor_rd_0_idx_bits,
  output         io_tensor_rd_0_data_valid,
  output [31:0]  io_tensor_rd_0_data_bits_0_0,
  output [31:0]  io_tensor_rd_0_data_bits_0_1,
  output [31:0]  io_tensor_rd_0_data_bits_0_2,
  output [31:0]  io_tensor_rd_0_data_bits_0_3,
  output [31:0]  io_tensor_rd_0_data_bits_0_4,
  output [31:0]  io_tensor_rd_0_data_bits_0_5,
  output [31:0]  io_tensor_rd_0_data_bits_0_6,
  output [31:0]  io_tensor_rd_0_data_bits_0_7,
  output [31:0]  io_tensor_rd_0_data_bits_0_8,
  output [31:0]  io_tensor_rd_0_data_bits_0_9,
  output [31:0]  io_tensor_rd_0_data_bits_0_10,
  output [31:0]  io_tensor_rd_0_data_bits_0_11,
  output [31:0]  io_tensor_rd_0_data_bits_0_12,
  output [31:0]  io_tensor_rd_0_data_bits_0_13,
  output [31:0]  io_tensor_rd_0_data_bits_0_14,
  output [31:0]  io_tensor_rd_0_data_bits_0_15,
  output [31:0]  io_tensor_rd_0_data_bits_0_16,
  output [31:0]  io_tensor_rd_0_data_bits_0_17,
  output [31:0]  io_tensor_rd_0_data_bits_0_18,
  output [31:0]  io_tensor_rd_0_data_bits_0_19,
  output [31:0]  io_tensor_rd_0_data_bits_0_20,
  output [31:0]  io_tensor_rd_0_data_bits_0_21,
  output [31:0]  io_tensor_rd_0_data_bits_0_22,
  output [31:0]  io_tensor_rd_0_data_bits_0_23,
  output [31:0]  io_tensor_rd_0_data_bits_0_24,
  output [31:0]  io_tensor_rd_0_data_bits_0_25,
  output [31:0]  io_tensor_rd_0_data_bits_0_26,
  output [31:0]  io_tensor_rd_0_data_bits_0_27,
  output [31:0]  io_tensor_rd_0_data_bits_0_28,
  output [31:0]  io_tensor_rd_0_data_bits_0_29,
  output [31:0]  io_tensor_rd_0_data_bits_0_30,
  output [31:0]  io_tensor_rd_0_data_bits_0_31,
  input          io_tensor_wr_0_valid,
  input  [6:0]   io_tensor_wr_0_bits_idx,
  input  [31:0]  io_tensor_wr_0_bits_data_0_0,
  input  [31:0]  io_tensor_wr_0_bits_data_0_1,
  input  [31:0]  io_tensor_wr_0_bits_data_0_2,
  input  [31:0]  io_tensor_wr_0_bits_data_0_3,
  input  [31:0]  io_tensor_wr_0_bits_data_0_4,
  input  [31:0]  io_tensor_wr_0_bits_data_0_5,
  input  [31:0]  io_tensor_wr_0_bits_data_0_6,
  input  [31:0]  io_tensor_wr_0_bits_data_0_7,
  input  [31:0]  io_tensor_wr_0_bits_data_0_8,
  input  [31:0]  io_tensor_wr_0_bits_data_0_9,
  input  [31:0]  io_tensor_wr_0_bits_data_0_10,
  input  [31:0]  io_tensor_wr_0_bits_data_0_11,
  input  [31:0]  io_tensor_wr_0_bits_data_0_12,
  input  [31:0]  io_tensor_wr_0_bits_data_0_13,
  input  [31:0]  io_tensor_wr_0_bits_data_0_14,
  input  [31:0]  io_tensor_wr_0_bits_data_0_15,
  input  [31:0]  io_tensor_wr_0_bits_data_0_16,
  input  [31:0]  io_tensor_wr_0_bits_data_0_17,
  input  [31:0]  io_tensor_wr_0_bits_data_0_18,
  input  [31:0]  io_tensor_wr_0_bits_data_0_19,
  input  [31:0]  io_tensor_wr_0_bits_data_0_20,
  input  [31:0]  io_tensor_wr_0_bits_data_0_21,
  input  [31:0]  io_tensor_wr_0_bits_data_0_22,
  input  [31:0]  io_tensor_wr_0_bits_data_0_23,
  input  [31:0]  io_tensor_wr_0_bits_data_0_24,
  input  [31:0]  io_tensor_wr_0_bits_data_0_25,
  input  [31:0]  io_tensor_wr_0_bits_data_0_26,
  input  [31:0]  io_tensor_wr_0_bits_data_0_27,
  input  [31:0]  io_tensor_wr_0_bits_data_0_28,
  input  [31:0]  io_tensor_wr_0_bits_data_0_29,
  input  [31:0]  io_tensor_wr_0_bits_data_0_30,
  input  [31:0]  io_tensor_wr_0_bits_data_0_31
);
  wire  tensorLoad_clock; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_reset; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_start; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_done; // @[TensorLoad.scala 71:28]
  wire [127:0] tensorLoad_io_inst; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_baddr; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_vme_rd_cmd_ready; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_vme_rd_cmd_valid; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_vme_rd_cmd_bits_addr; // @[TensorLoad.scala 71:28]
  wire [3:0] tensorLoad_io_vme_rd_cmd_bits_len; // @[TensorLoad.scala 71:28]
  wire [20:0] tensorLoad_io_vme_rd_cmd_bits_tag; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_vme_rd_data_ready; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_vme_rd_data_valid; // @[TensorLoad.scala 71:28]
  wire [63:0] tensorLoad_io_vme_rd_data_bits_data; // @[TensorLoad.scala 71:28]
  wire [20:0] tensorLoad_io_vme_rd_data_bits_tag; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_tensor_rd_0_idx_valid; // @[TensorLoad.scala 71:28]
  wire [6:0] tensorLoad_io_tensor_rd_0_idx_bits; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_tensor_rd_0_data_valid; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_0; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_1; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_2; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_3; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_4; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_5; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_6; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_7; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_8; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_9; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_10; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_11; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_12; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_13; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_14; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_15; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_16; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_17; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_18; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_19; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_20; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_21; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_22; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_23; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_24; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_25; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_26; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_27; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_28; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_29; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_30; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_rd_0_data_bits_0_31; // @[TensorLoad.scala 71:28]
  wire  tensorLoad_io_tensor_wr_0_valid; // @[TensorLoad.scala 71:28]
  wire [6:0] tensorLoad_io_tensor_wr_0_bits_idx; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_0; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_1; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_2; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_3; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_4; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_5; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_6; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_7; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_8; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_9; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_10; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_11; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_12; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_13; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_14; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_15; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_16; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_17; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_18; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_19; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_20; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_21; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_22; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_23; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_24; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_25; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_26; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_27; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_28; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_29; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_30; // @[TensorLoad.scala 71:28]
  wire [31:0] tensorLoad_io_tensor_wr_0_bits_data_0_31; // @[TensorLoad.scala 71:28]
  TensorLoadNarrowVME_2 tensorLoad ( // @[TensorLoad.scala 71:28]
    .clock(tensorLoad_clock),
    .reset(tensorLoad_reset),
    .io_start(tensorLoad_io_start),
    .io_done(tensorLoad_io_done),
    .io_inst(tensorLoad_io_inst),
    .io_baddr(tensorLoad_io_baddr),
    .io_vme_rd_cmd_ready(tensorLoad_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(tensorLoad_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(tensorLoad_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(tensorLoad_io_vme_rd_cmd_bits_len),
    .io_vme_rd_cmd_bits_tag(tensorLoad_io_vme_rd_cmd_bits_tag),
    .io_vme_rd_data_ready(tensorLoad_io_vme_rd_data_ready),
    .io_vme_rd_data_valid(tensorLoad_io_vme_rd_data_valid),
    .io_vme_rd_data_bits_data(tensorLoad_io_vme_rd_data_bits_data),
    .io_vme_rd_data_bits_tag(tensorLoad_io_vme_rd_data_bits_tag),
    .io_tensor_rd_0_idx_valid(tensorLoad_io_tensor_rd_0_idx_valid),
    .io_tensor_rd_0_idx_bits(tensorLoad_io_tensor_rd_0_idx_bits),
    .io_tensor_rd_0_data_valid(tensorLoad_io_tensor_rd_0_data_valid),
    .io_tensor_rd_0_data_bits_0_0(tensorLoad_io_tensor_rd_0_data_bits_0_0),
    .io_tensor_rd_0_data_bits_0_1(tensorLoad_io_tensor_rd_0_data_bits_0_1),
    .io_tensor_rd_0_data_bits_0_2(tensorLoad_io_tensor_rd_0_data_bits_0_2),
    .io_tensor_rd_0_data_bits_0_3(tensorLoad_io_tensor_rd_0_data_bits_0_3),
    .io_tensor_rd_0_data_bits_0_4(tensorLoad_io_tensor_rd_0_data_bits_0_4),
    .io_tensor_rd_0_data_bits_0_5(tensorLoad_io_tensor_rd_0_data_bits_0_5),
    .io_tensor_rd_0_data_bits_0_6(tensorLoad_io_tensor_rd_0_data_bits_0_6),
    .io_tensor_rd_0_data_bits_0_7(tensorLoad_io_tensor_rd_0_data_bits_0_7),
    .io_tensor_rd_0_data_bits_0_8(tensorLoad_io_tensor_rd_0_data_bits_0_8),
    .io_tensor_rd_0_data_bits_0_9(tensorLoad_io_tensor_rd_0_data_bits_0_9),
    .io_tensor_rd_0_data_bits_0_10(tensorLoad_io_tensor_rd_0_data_bits_0_10),
    .io_tensor_rd_0_data_bits_0_11(tensorLoad_io_tensor_rd_0_data_bits_0_11),
    .io_tensor_rd_0_data_bits_0_12(tensorLoad_io_tensor_rd_0_data_bits_0_12),
    .io_tensor_rd_0_data_bits_0_13(tensorLoad_io_tensor_rd_0_data_bits_0_13),
    .io_tensor_rd_0_data_bits_0_14(tensorLoad_io_tensor_rd_0_data_bits_0_14),
    .io_tensor_rd_0_data_bits_0_15(tensorLoad_io_tensor_rd_0_data_bits_0_15),
    .io_tensor_rd_0_data_bits_0_16(tensorLoad_io_tensor_rd_0_data_bits_0_16),
    .io_tensor_rd_0_data_bits_0_17(tensorLoad_io_tensor_rd_0_data_bits_0_17),
    .io_tensor_rd_0_data_bits_0_18(tensorLoad_io_tensor_rd_0_data_bits_0_18),
    .io_tensor_rd_0_data_bits_0_19(tensorLoad_io_tensor_rd_0_data_bits_0_19),
    .io_tensor_rd_0_data_bits_0_20(tensorLoad_io_tensor_rd_0_data_bits_0_20),
    .io_tensor_rd_0_data_bits_0_21(tensorLoad_io_tensor_rd_0_data_bits_0_21),
    .io_tensor_rd_0_data_bits_0_22(tensorLoad_io_tensor_rd_0_data_bits_0_22),
    .io_tensor_rd_0_data_bits_0_23(tensorLoad_io_tensor_rd_0_data_bits_0_23),
    .io_tensor_rd_0_data_bits_0_24(tensorLoad_io_tensor_rd_0_data_bits_0_24),
    .io_tensor_rd_0_data_bits_0_25(tensorLoad_io_tensor_rd_0_data_bits_0_25),
    .io_tensor_rd_0_data_bits_0_26(tensorLoad_io_tensor_rd_0_data_bits_0_26),
    .io_tensor_rd_0_data_bits_0_27(tensorLoad_io_tensor_rd_0_data_bits_0_27),
    .io_tensor_rd_0_data_bits_0_28(tensorLoad_io_tensor_rd_0_data_bits_0_28),
    .io_tensor_rd_0_data_bits_0_29(tensorLoad_io_tensor_rd_0_data_bits_0_29),
    .io_tensor_rd_0_data_bits_0_30(tensorLoad_io_tensor_rd_0_data_bits_0_30),
    .io_tensor_rd_0_data_bits_0_31(tensorLoad_io_tensor_rd_0_data_bits_0_31),
    .io_tensor_wr_0_valid(tensorLoad_io_tensor_wr_0_valid),
    .io_tensor_wr_0_bits_idx(tensorLoad_io_tensor_wr_0_bits_idx),
    .io_tensor_wr_0_bits_data_0_0(tensorLoad_io_tensor_wr_0_bits_data_0_0),
    .io_tensor_wr_0_bits_data_0_1(tensorLoad_io_tensor_wr_0_bits_data_0_1),
    .io_tensor_wr_0_bits_data_0_2(tensorLoad_io_tensor_wr_0_bits_data_0_2),
    .io_tensor_wr_0_bits_data_0_3(tensorLoad_io_tensor_wr_0_bits_data_0_3),
    .io_tensor_wr_0_bits_data_0_4(tensorLoad_io_tensor_wr_0_bits_data_0_4),
    .io_tensor_wr_0_bits_data_0_5(tensorLoad_io_tensor_wr_0_bits_data_0_5),
    .io_tensor_wr_0_bits_data_0_6(tensorLoad_io_tensor_wr_0_bits_data_0_6),
    .io_tensor_wr_0_bits_data_0_7(tensorLoad_io_tensor_wr_0_bits_data_0_7),
    .io_tensor_wr_0_bits_data_0_8(tensorLoad_io_tensor_wr_0_bits_data_0_8),
    .io_tensor_wr_0_bits_data_0_9(tensorLoad_io_tensor_wr_0_bits_data_0_9),
    .io_tensor_wr_0_bits_data_0_10(tensorLoad_io_tensor_wr_0_bits_data_0_10),
    .io_tensor_wr_0_bits_data_0_11(tensorLoad_io_tensor_wr_0_bits_data_0_11),
    .io_tensor_wr_0_bits_data_0_12(tensorLoad_io_tensor_wr_0_bits_data_0_12),
    .io_tensor_wr_0_bits_data_0_13(tensorLoad_io_tensor_wr_0_bits_data_0_13),
    .io_tensor_wr_0_bits_data_0_14(tensorLoad_io_tensor_wr_0_bits_data_0_14),
    .io_tensor_wr_0_bits_data_0_15(tensorLoad_io_tensor_wr_0_bits_data_0_15),
    .io_tensor_wr_0_bits_data_0_16(tensorLoad_io_tensor_wr_0_bits_data_0_16),
    .io_tensor_wr_0_bits_data_0_17(tensorLoad_io_tensor_wr_0_bits_data_0_17),
    .io_tensor_wr_0_bits_data_0_18(tensorLoad_io_tensor_wr_0_bits_data_0_18),
    .io_tensor_wr_0_bits_data_0_19(tensorLoad_io_tensor_wr_0_bits_data_0_19),
    .io_tensor_wr_0_bits_data_0_20(tensorLoad_io_tensor_wr_0_bits_data_0_20),
    .io_tensor_wr_0_bits_data_0_21(tensorLoad_io_tensor_wr_0_bits_data_0_21),
    .io_tensor_wr_0_bits_data_0_22(tensorLoad_io_tensor_wr_0_bits_data_0_22),
    .io_tensor_wr_0_bits_data_0_23(tensorLoad_io_tensor_wr_0_bits_data_0_23),
    .io_tensor_wr_0_bits_data_0_24(tensorLoad_io_tensor_wr_0_bits_data_0_24),
    .io_tensor_wr_0_bits_data_0_25(tensorLoad_io_tensor_wr_0_bits_data_0_25),
    .io_tensor_wr_0_bits_data_0_26(tensorLoad_io_tensor_wr_0_bits_data_0_26),
    .io_tensor_wr_0_bits_data_0_27(tensorLoad_io_tensor_wr_0_bits_data_0_27),
    .io_tensor_wr_0_bits_data_0_28(tensorLoad_io_tensor_wr_0_bits_data_0_28),
    .io_tensor_wr_0_bits_data_0_29(tensorLoad_io_tensor_wr_0_bits_data_0_29),
    .io_tensor_wr_0_bits_data_0_30(tensorLoad_io_tensor_wr_0_bits_data_0_30),
    .io_tensor_wr_0_bits_data_0_31(tensorLoad_io_tensor_wr_0_bits_data_0_31)
  );
  assign io_done = tensorLoad_io_done; // @[TensorLoad.scala 72:8]
  assign io_vme_rd_cmd_valid = tensorLoad_io_vme_rd_cmd_valid; // @[TensorLoad.scala 72:8]
  assign io_vme_rd_cmd_bits_addr = tensorLoad_io_vme_rd_cmd_bits_addr; // @[TensorLoad.scala 72:8]
  assign io_vme_rd_cmd_bits_len = tensorLoad_io_vme_rd_cmd_bits_len; // @[TensorLoad.scala 72:8]
  assign io_vme_rd_cmd_bits_tag = tensorLoad_io_vme_rd_cmd_bits_tag; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_valid = tensorLoad_io_tensor_rd_0_data_valid; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_0 = tensorLoad_io_tensor_rd_0_data_bits_0_0; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_1 = tensorLoad_io_tensor_rd_0_data_bits_0_1; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_2 = tensorLoad_io_tensor_rd_0_data_bits_0_2; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_3 = tensorLoad_io_tensor_rd_0_data_bits_0_3; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_4 = tensorLoad_io_tensor_rd_0_data_bits_0_4; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_5 = tensorLoad_io_tensor_rd_0_data_bits_0_5; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_6 = tensorLoad_io_tensor_rd_0_data_bits_0_6; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_7 = tensorLoad_io_tensor_rd_0_data_bits_0_7; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_8 = tensorLoad_io_tensor_rd_0_data_bits_0_8; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_9 = tensorLoad_io_tensor_rd_0_data_bits_0_9; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_10 = tensorLoad_io_tensor_rd_0_data_bits_0_10; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_11 = tensorLoad_io_tensor_rd_0_data_bits_0_11; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_12 = tensorLoad_io_tensor_rd_0_data_bits_0_12; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_13 = tensorLoad_io_tensor_rd_0_data_bits_0_13; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_14 = tensorLoad_io_tensor_rd_0_data_bits_0_14; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_15 = tensorLoad_io_tensor_rd_0_data_bits_0_15; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_16 = tensorLoad_io_tensor_rd_0_data_bits_0_16; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_17 = tensorLoad_io_tensor_rd_0_data_bits_0_17; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_18 = tensorLoad_io_tensor_rd_0_data_bits_0_18; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_19 = tensorLoad_io_tensor_rd_0_data_bits_0_19; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_20 = tensorLoad_io_tensor_rd_0_data_bits_0_20; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_21 = tensorLoad_io_tensor_rd_0_data_bits_0_21; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_22 = tensorLoad_io_tensor_rd_0_data_bits_0_22; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_23 = tensorLoad_io_tensor_rd_0_data_bits_0_23; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_24 = tensorLoad_io_tensor_rd_0_data_bits_0_24; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_25 = tensorLoad_io_tensor_rd_0_data_bits_0_25; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_26 = tensorLoad_io_tensor_rd_0_data_bits_0_26; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_27 = tensorLoad_io_tensor_rd_0_data_bits_0_27; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_28 = tensorLoad_io_tensor_rd_0_data_bits_0_28; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_29 = tensorLoad_io_tensor_rd_0_data_bits_0_29; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_30 = tensorLoad_io_tensor_rd_0_data_bits_0_30; // @[TensorLoad.scala 72:8]
  assign io_tensor_rd_0_data_bits_0_31 = tensorLoad_io_tensor_rd_0_data_bits_0_31; // @[TensorLoad.scala 72:8]
  assign tensorLoad_clock = clock;
  assign tensorLoad_reset = reset;
  assign tensorLoad_io_start = io_start; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_inst = io_inst; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_baddr = io_baddr; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_vme_rd_cmd_ready = io_vme_rd_cmd_ready; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_vme_rd_data_valid = io_vme_rd_data_valid; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_vme_rd_data_bits_data = io_vme_rd_data_bits_data; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_vme_rd_data_bits_tag = io_vme_rd_data_bits_tag; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_rd_0_idx_valid = io_tensor_rd_0_idx_valid; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_rd_0_idx_bits = io_tensor_rd_0_idx_bits; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_valid = io_tensor_wr_0_valid; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_idx = io_tensor_wr_0_bits_idx; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_0 = io_tensor_wr_0_bits_data_0_0; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_1 = io_tensor_wr_0_bits_data_0_1; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_2 = io_tensor_wr_0_bits_data_0_2; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_3 = io_tensor_wr_0_bits_data_0_3; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_4 = io_tensor_wr_0_bits_data_0_4; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_5 = io_tensor_wr_0_bits_data_0_5; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_6 = io_tensor_wr_0_bits_data_0_6; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_7 = io_tensor_wr_0_bits_data_0_7; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_8 = io_tensor_wr_0_bits_data_0_8; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_9 = io_tensor_wr_0_bits_data_0_9; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_10 = io_tensor_wr_0_bits_data_0_10; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_11 = io_tensor_wr_0_bits_data_0_11; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_12 = io_tensor_wr_0_bits_data_0_12; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_13 = io_tensor_wr_0_bits_data_0_13; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_14 = io_tensor_wr_0_bits_data_0_14; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_15 = io_tensor_wr_0_bits_data_0_15; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_16 = io_tensor_wr_0_bits_data_0_16; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_17 = io_tensor_wr_0_bits_data_0_17; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_18 = io_tensor_wr_0_bits_data_0_18; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_19 = io_tensor_wr_0_bits_data_0_19; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_20 = io_tensor_wr_0_bits_data_0_20; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_21 = io_tensor_wr_0_bits_data_0_21; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_22 = io_tensor_wr_0_bits_data_0_22; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_23 = io_tensor_wr_0_bits_data_0_23; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_24 = io_tensor_wr_0_bits_data_0_24; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_25 = io_tensor_wr_0_bits_data_0_25; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_26 = io_tensor_wr_0_bits_data_0_26; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_27 = io_tensor_wr_0_bits_data_0_27; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_28 = io_tensor_wr_0_bits_data_0_28; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_29 = io_tensor_wr_0_bits_data_0_29; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_30 = io_tensor_wr_0_bits_data_0_30; // @[TensorLoad.scala 72:8]
  assign tensorLoad_io_tensor_wr_0_bits_data_0_31 = io_tensor_wr_0_bits_data_0_31; // @[TensorLoad.scala 72:8]
endmodule
module TensorGemmIndexGenerator(
  input         clock,
  input         reset,
  input         io_start,
  output        io_last,
  input  [9:0]  io_dec_wgt_1,
  input  [9:0]  io_dec_wgt_0,
  input  [10:0] io_dec_inp_1,
  input  [10:0] io_dec_inp_0,
  input  [10:0] io_dec_acc_1,
  input  [10:0] io_dec_acc_0,
  input  [13:0] io_dec_lp_1,
  input  [13:0] io_dec_lp_0,
  input  [13:0] io_dec_uop_end,
  input  [12:0] io_dec_uop_begin,
  output [6:0]  io_acc_i,
  output [6:0]  io_inp_i,
  output [5:0]  io_wgt_i,
  output [6:0]  io_uop_idx,
  output        io_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg  running; // @[TensorGemm.scala 238:24]
  wire  _T = ~running; // @[TensorGemm.scala 239:8]
  wire  _GEN_0 = io_last ? 1'h0 : running; // @[TensorGemm.scala 241:23 242:13 238:24]
  wire  _GEN_1 = ~running & io_start | _GEN_0; // @[TensorGemm.scala 239:30 240:13]
  reg [13:0] cnt_i; // @[TensorGemm.scala 245:18]
  reg [6:0] acc_i; // @[TensorGemm.scala 246:18]
  reg [6:0] inp_i; // @[TensorGemm.scala 247:18]
  reg [5:0] wgt_i; // @[TensorGemm.scala 248:18]
  reg [13:0] cnt_o; // @[TensorGemm.scala 250:18]
  reg [6:0] acc_o; // @[TensorGemm.scala 251:18]
  reg [6:0] inp_o; // @[TensorGemm.scala 252:18]
  reg [5:0] wgt_o; // @[TensorGemm.scala 253:18]
  reg [13:0] uop_idx; // @[TensorGemm.scala 255:20]
  wire [13:0] _T_4 = io_dec_uop_end - 14'h1; // @[TensorGemm.scala 268:38]
  wire [13:0] _uop_idx_T_1 = uop_idx + 14'h1; // @[TensorGemm.scala 269:26]
  wire [13:0] _T_7 = io_dec_lp_1 - 14'h1; // @[TensorGemm.scala 272:35]
  wire [13:0] _cnt_i_T_1 = cnt_i + 14'h1; // @[TensorGemm.scala 273:24]
  wire [10:0] _GEN_40 = {{4'd0}, acc_i}; // @[TensorGemm.scala 274:24]
  wire [10:0] _acc_i_T_1 = _GEN_40 + io_dec_acc_1; // @[TensorGemm.scala 274:24]
  wire [10:0] _GEN_41 = {{4'd0}, inp_i}; // @[TensorGemm.scala 275:24]
  wire [10:0] _inp_i_T_1 = _GEN_41 + io_dec_inp_1; // @[TensorGemm.scala 275:24]
  wire [9:0] _GEN_42 = {{4'd0}, wgt_i}; // @[TensorGemm.scala 276:24]
  wire [9:0] _wgt_i_T_1 = _GEN_42 + io_dec_wgt_1; // @[TensorGemm.scala 276:24]
  wire [13:0] _T_10 = io_dec_lp_0 - 14'h1; // @[TensorGemm.scala 278:37]
  wire [10:0] _GEN_43 = {{4'd0}, acc_o}; // @[TensorGemm.scala 279:31]
  wire [10:0] acc_tmp = _GEN_43 + io_dec_acc_0; // @[TensorGemm.scala 279:31]
  wire [10:0] _GEN_44 = {{4'd0}, inp_o}; // @[TensorGemm.scala 280:31]
  wire [10:0] inp_tmp = _GEN_44 + io_dec_inp_0; // @[TensorGemm.scala 280:31]
  wire [9:0] _GEN_45 = {{4'd0}, wgt_o}; // @[TensorGemm.scala 281:31]
  wire [9:0] wgt_tmp = _GEN_45 + io_dec_wgt_0; // @[TensorGemm.scala 281:31]
  wire [13:0] _cnt_o_T_1 = cnt_o + 14'h1; // @[TensorGemm.scala 282:26]
  wire [10:0] _GEN_3 = cnt_o != _T_10 ? acc_tmp : {{4'd0}, acc_o}; // @[TensorGemm.scala 278:44 283:17 251:18]
  wire [10:0] _GEN_4 = cnt_o != _T_10 ? inp_tmp : {{4'd0}, inp_o}; // @[TensorGemm.scala 278:44 284:17 252:18]
  wire [9:0] _GEN_5 = cnt_o != _T_10 ? wgt_tmp : {{4'd0}, wgt_o}; // @[TensorGemm.scala 278:44 285:17 253:18]
  wire [10:0] _GEN_7 = cnt_o != _T_10 ? acc_tmp : {{4'd0}, acc_i}; // @[TensorGemm.scala 278:44 287:17 246:18]
  wire [10:0] _GEN_8 = cnt_o != _T_10 ? inp_tmp : {{4'd0}, inp_i}; // @[TensorGemm.scala 278:44 288:17 247:18]
  wire [9:0] _GEN_9 = cnt_o != _T_10 ? wgt_tmp : {{4'd0}, wgt_i}; // @[TensorGemm.scala 278:44 289:17 248:18]
  wire  _GEN_10 = cnt_o != _T_10 ? 1'h0 : 1'h1; // @[TensorGemm.scala 236:11 278:44 291:19]
  wire [10:0] _GEN_12 = cnt_i != _T_7 ? _acc_i_T_1 : _GEN_7; // @[TensorGemm.scala 272:42 274:15]
  wire [10:0] _GEN_13 = cnt_i != _T_7 ? _inp_i_T_1 : _GEN_8; // @[TensorGemm.scala 272:42 275:15]
  wire [9:0] _GEN_14 = cnt_i != _T_7 ? _wgt_i_T_1 : _GEN_9; // @[TensorGemm.scala 272:42 276:15]
  wire [10:0] _GEN_16 = cnt_i != _T_7 ? {{4'd0}, acc_o} : _GEN_3; // @[TensorGemm.scala 251:18 272:42]
  wire [10:0] _GEN_17 = cnt_i != _T_7 ? {{4'd0}, inp_o} : _GEN_4; // @[TensorGemm.scala 252:18 272:42]
  wire [9:0] _GEN_18 = cnt_i != _T_7 ? {{4'd0}, wgt_o} : _GEN_5; // @[TensorGemm.scala 253:18 272:42]
  wire  _GEN_19 = cnt_i != _T_7 ? 1'h0 : _GEN_10; // @[TensorGemm.scala 236:11 272:42]
  wire [10:0] _GEN_22 = uop_idx != _T_4 ? {{4'd0}, acc_i} : _GEN_12; // @[TensorGemm.scala 246:18 268:45]
  wire [10:0] _GEN_23 = uop_idx != _T_4 ? {{4'd0}, inp_i} : _GEN_13; // @[TensorGemm.scala 247:18 268:45]
  wire [9:0] _GEN_24 = uop_idx != _T_4 ? {{4'd0}, wgt_i} : _GEN_14; // @[TensorGemm.scala 248:18 268:45]
  wire [10:0] _GEN_26 = uop_idx != _T_4 ? {{4'd0}, acc_o} : _GEN_16; // @[TensorGemm.scala 251:18 268:45]
  wire [10:0] _GEN_27 = uop_idx != _T_4 ? {{4'd0}, inp_o} : _GEN_17; // @[TensorGemm.scala 252:18 268:45]
  wire [9:0] _GEN_28 = uop_idx != _T_4 ? {{4'd0}, wgt_o} : _GEN_18; // @[TensorGemm.scala 253:18 268:45]
  wire  _GEN_29 = uop_idx != _T_4 ? 1'h0 : _GEN_19; // @[TensorGemm.scala 236:11 268:45]
  wire [10:0] _GEN_31 = _T ? 11'h0 : _GEN_22; // @[TensorGemm.scala 263:18 264:25]
  wire [10:0] _GEN_32 = _T ? 11'h0 : _GEN_23; // @[TensorGemm.scala 263:18 264:39]
  wire [9:0] _GEN_33 = _T ? 10'h0 : _GEN_24; // @[TensorGemm.scala 263:18 264:53]
  wire [10:0] _GEN_35 = _T ? 11'h0 : _GEN_26; // @[TensorGemm.scala 263:18 265:25]
  wire [10:0] _GEN_36 = _T ? 11'h0 : _GEN_27; // @[TensorGemm.scala 263:18 265:39]
  wire [9:0] _GEN_37 = _T ? 10'h0 : _GEN_28; // @[TensorGemm.scala 263:18 265:53]
  assign io_last = _T ? 1'h0 : _GEN_29; // @[TensorGemm.scala 236:11 263:18]
  assign io_acc_i = acc_i; // @[TensorGemm.scala 258:12]
  assign io_inp_i = inp_i; // @[TensorGemm.scala 259:12]
  assign io_wgt_i = wgt_i; // @[TensorGemm.scala 260:12]
  assign io_uop_idx = uop_idx[6:0]; // @[TensorGemm.scala 261:14]
  assign io_valid = running; // @[TensorGemm.scala 257:12]
  always @(posedge clock) begin
    if (reset) begin // @[TensorGemm.scala 238:24]
      running <= 1'h0; // @[TensorGemm.scala 238:24]
    end else begin
      running <= _GEN_1;
    end
    if (_T) begin // @[TensorGemm.scala 263:18]
      cnt_i <= 14'h0; // @[TensorGemm.scala 264:11]
    end else if (!(uop_idx != _T_4)) begin // @[TensorGemm.scala 268:45]
      if (cnt_i != _T_7) begin // @[TensorGemm.scala 272:42]
        cnt_i <= _cnt_i_T_1; // @[TensorGemm.scala 273:15]
      end else if (cnt_o != _T_10) begin // @[TensorGemm.scala 278:44]
        cnt_i <= 14'h0; // @[TensorGemm.scala 286:17]
      end
    end
    acc_i <= _GEN_31[6:0];
    inp_i <= _GEN_32[6:0];
    wgt_i <= _GEN_33[5:0];
    if (_T) begin // @[TensorGemm.scala 263:18]
      cnt_o <= 14'h0; // @[TensorGemm.scala 265:11]
    end else if (!(uop_idx != _T_4)) begin // @[TensorGemm.scala 268:45]
      if (!(cnt_i != _T_7)) begin // @[TensorGemm.scala 272:42]
        if (cnt_o != _T_10) begin // @[TensorGemm.scala 278:44]
          cnt_o <= _cnt_o_T_1; // @[TensorGemm.scala 282:17]
        end
      end
    end
    acc_o <= _GEN_35[6:0];
    inp_o <= _GEN_36[6:0];
    wgt_o <= _GEN_37[5:0];
    if (_T) begin // @[TensorGemm.scala 263:18]
      uop_idx <= {{1'd0}, io_dec_uop_begin}; // @[TensorGemm.scala 266:13]
    end else if (uop_idx != _T_4) begin // @[TensorGemm.scala 268:45]
      uop_idx <= _uop_idx_T_1; // @[TensorGemm.scala 269:15]
    end else begin
      uop_idx <= {{1'd0}, io_dec_uop_begin}; // @[TensorGemm.scala 271:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  running = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  cnt_i = _RAND_1[13:0];
  _RAND_2 = {1{`RANDOM}};
  acc_i = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  inp_i = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  wgt_i = _RAND_4[5:0];
  _RAND_5 = {1{`RANDOM}};
  cnt_o = _RAND_5[13:0];
  _RAND_6 = {1{`RANDOM}};
  acc_o = _RAND_6[6:0];
  _RAND_7 = {1{`RANDOM}};
  inp_o = _RAND_7[6:0];
  _RAND_8 = {1{`RANDOM}};
  wgt_o = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  uop_idx = _RAND_9[13:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Pipe(
  input   clock,
  input   reset,
  input   io_enq_valid,
  input   io_enq_bits,
  output  io_deq_valid,
  output  io_deq_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  io_deq_v; // @[Valid.scala 127:22]
  reg  io_deq_b; // @[Reg.scala 16:16]
  reg  io_deq_outPipe_valid; // @[Valid.scala 127:22]
  reg  io_deq_outPipe_bits; // @[Reg.scala 16:16]
  reg  io_deq_outPipe_valid_1; // @[Valid.scala 127:22]
  reg  io_deq_outPipe_bits_1; // @[Reg.scala 16:16]
  assign io_deq_valid = io_deq_outPipe_valid_1; // @[Valid.scala 122:21 123:17]
  assign io_deq_bits = io_deq_outPipe_bits_1; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      io_deq_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_deq_v <= io_enq_valid; // @[Valid.scala 127:22]
    end
    if (io_enq_valid) begin // @[Reg.scala 17:18]
      io_deq_b <= io_enq_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_deq_outPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_deq_outPipe_valid <= io_deq_v; // @[Valid.scala 127:22]
    end
    if (io_deq_v) begin // @[Reg.scala 17:18]
      io_deq_outPipe_bits <= io_deq_b; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_deq_outPipe_valid_1 <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_deq_outPipe_valid_1 <= io_deq_outPipe_valid; // @[Valid.scala 127:22]
    end
    if (io_deq_outPipe_valid) begin // @[Reg.scala 17:18]
      io_deq_outPipe_bits_1 <= io_deq_outPipe_bits; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_deq_v = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  io_deq_b = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  io_deq_outPipe_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  io_deq_outPipe_bits = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  io_deq_outPipe_valid_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  io_deq_outPipe_bits_1 = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Pipe_1(
  input        clock,
  input        reset,
  input        io_enq_valid,
  input  [6:0] io_enq_bits,
  output       io_deq_valid,
  output [6:0] io_deq_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  io_deq_v; // @[Valid.scala 127:22]
  reg [6:0] io_deq_b; // @[Reg.scala 16:16]
  assign io_deq_valid = io_deq_v; // @[Valid.scala 122:21 123:17]
  assign io_deq_bits = io_deq_b; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      io_deq_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_deq_v <= io_enq_valid; // @[Valid.scala 127:22]
    end
    if (io_enq_valid) begin // @[Reg.scala 17:18]
      io_deq_b <= io_enq_bits; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_deq_v = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  io_deq_b = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Pipe_2(
  input        clock,
  input        reset,
  input        io_enq_valid,
  input  [6:0] io_enq_bits,
  output       io_deq_valid,
  output [6:0] io_deq_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg  io_deq_v; // @[Valid.scala 127:22]
  reg [6:0] io_deq_b; // @[Reg.scala 16:16]
  reg  io_deq_outPipe_valid; // @[Valid.scala 127:22]
  reg [6:0] io_deq_outPipe_bits; // @[Reg.scala 16:16]
  assign io_deq_valid = io_deq_outPipe_valid; // @[Valid.scala 122:21 123:17]
  assign io_deq_bits = io_deq_outPipe_bits; // @[Valid.scala 122:21 124:16]
  always @(posedge clock) begin
    if (reset) begin // @[Valid.scala 127:22]
      io_deq_v <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_deq_v <= io_enq_valid; // @[Valid.scala 127:22]
    end
    if (io_enq_valid) begin // @[Reg.scala 17:18]
      io_deq_b <= io_enq_bits; // @[Reg.scala 17:22]
    end
    if (reset) begin // @[Valid.scala 127:22]
      io_deq_outPipe_valid <= 1'h0; // @[Valid.scala 127:22]
    end else begin
      io_deq_outPipe_valid <= io_deq_v; // @[Valid.scala 127:22]
    end
    if (io_deq_v) begin // @[Reg.scala 17:18]
      io_deq_outPipe_bits <= io_deq_b; // @[Reg.scala 17:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  io_deq_v = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  io_deq_b = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  io_deq_outPipe_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  io_deq_outPipe_bits = _RAND_3[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module MAC(
  input         clock,
  input  [7:0]  io_a,
  input  [7:0]  io_b,
  output [16:0] io_y
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] rA; // @[TensorGemm.scala 38:31]
  reg [7:0] rB; // @[TensorGemm.scala 39:31]
  wire [15:0] mult = $signed(rA) * $signed(rB); // @[TensorGemm.scala 42:14]
  assign io_y = {{1{mult[15]}},mult}; // @[TensorGemm.scala 43:30]
  always @(posedge clock) begin
    rA <= io_a; // @[TensorGemm.scala 38:31]
    rB <= io_b; // @[TensorGemm.scala 39:31]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rA = _RAND_0[7:0];
  _RAND_1 = {1{`RANDOM}};
  rB = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Adder(
  input  [16:0] io_a,
  input  [16:0] io_b,
  output [17:0] io_y
);
  assign io_y = $signed(io_a) + $signed(io_b); // @[TensorGemm.scala 81:13]
endmodule
module Adder_8(
  input  [17:0] io_a,
  input  [17:0] io_b,
  output [18:0] io_y
);
  assign io_y = $signed(io_a) + $signed(io_b); // @[TensorGemm.scala 81:13]
endmodule
module PipeAdder(
  input         clock,
  input  [18:0] io_a,
  input  [18:0] io_b,
  output [19:0] io_y
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [18:0] rA; // @[TensorGemm.scala 63:19]
  reg [18:0] rB; // @[TensorGemm.scala 64:19]
  assign io_y = $signed(rA) + $signed(rB); // @[TensorGemm.scala 65:13]
  always @(posedge clock) begin
    rA <= io_a; // @[TensorGemm.scala 63:19]
    rB <= io_b; // @[TensorGemm.scala 64:19]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rA = _RAND_0[18:0];
  _RAND_1 = {1{`RANDOM}};
  rB = _RAND_1[18:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Adder_12(
  input  [19:0] io_a,
  input  [19:0] io_b,
  output [20:0] io_y
);
  assign io_y = $signed(io_a) + $signed(io_b); // @[TensorGemm.scala 81:13]
endmodule
module DotProduct(
  input         clock,
  input  [7:0]  io_a_0,
  input  [7:0]  io_a_1,
  input  [7:0]  io_a_2,
  input  [7:0]  io_a_3,
  input  [7:0]  io_a_4,
  input  [7:0]  io_a_5,
  input  [7:0]  io_a_6,
  input  [7:0]  io_a_7,
  input  [7:0]  io_a_8,
  input  [7:0]  io_a_9,
  input  [7:0]  io_a_10,
  input  [7:0]  io_a_11,
  input  [7:0]  io_a_12,
  input  [7:0]  io_a_13,
  input  [7:0]  io_a_14,
  input  [7:0]  io_a_15,
  input  [7:0]  io_b_0,
  input  [7:0]  io_b_1,
  input  [7:0]  io_b_2,
  input  [7:0]  io_b_3,
  input  [7:0]  io_b_4,
  input  [7:0]  io_b_5,
  input  [7:0]  io_b_6,
  input  [7:0]  io_b_7,
  input  [7:0]  io_b_8,
  input  [7:0]  io_b_9,
  input  [7:0]  io_b_10,
  input  [7:0]  io_b_11,
  input  [7:0]  io_b_12,
  input  [7:0]  io_b_13,
  input  [7:0]  io_b_14,
  input  [7:0]  io_b_15,
  output [20:0] io_y
);
  wire  m_0_clock; // @[TensorGemm.scala 100:32]
  wire [7:0] m_0_io_a; // @[TensorGemm.scala 100:32]
  wire [7:0] m_0_io_b; // @[TensorGemm.scala 100:32]
  wire [16:0] m_0_io_y; // @[TensorGemm.scala 100:32]
  wire  m_1_clock; // @[TensorGemm.scala 100:32]
  wire [7:0] m_1_io_a; // @[TensorGemm.scala 100:32]
  wire [7:0] m_1_io_b; // @[TensorGemm.scala 100:32]
  wire [16:0] m_1_io_y; // @[TensorGemm.scala 100:32]
  wire  m_2_clock; // @[TensorGemm.scala 100:32]
  wire [7:0] m_2_io_a; // @[TensorGemm.scala 100:32]
  wire [7:0] m_2_io_b; // @[TensorGemm.scala 100:32]
  wire [16:0] m_2_io_y; // @[TensorGemm.scala 100:32]
  wire  m_3_clock; // @[TensorGemm.scala 100:32]
  wire [7:0] m_3_io_a; // @[TensorGemm.scala 100:32]
  wire [7:0] m_3_io_b; // @[TensorGemm.scala 100:32]
  wire [16:0] m_3_io_y; // @[TensorGemm.scala 100:32]
  wire  m_4_clock; // @[TensorGemm.scala 100:32]
  wire [7:0] m_4_io_a; // @[TensorGemm.scala 100:32]
  wire [7:0] m_4_io_b; // @[TensorGemm.scala 100:32]
  wire [16:0] m_4_io_y; // @[TensorGemm.scala 100:32]
  wire  m_5_clock; // @[TensorGemm.scala 100:32]
  wire [7:0] m_5_io_a; // @[TensorGemm.scala 100:32]
  wire [7:0] m_5_io_b; // @[TensorGemm.scala 100:32]
  wire [16:0] m_5_io_y; // @[TensorGemm.scala 100:32]
  wire  m_6_clock; // @[TensorGemm.scala 100:32]
  wire [7:0] m_6_io_a; // @[TensorGemm.scala 100:32]
  wire [7:0] m_6_io_b; // @[TensorGemm.scala 100:32]
  wire [16:0] m_6_io_y; // @[TensorGemm.scala 100:32]
  wire  m_7_clock; // @[TensorGemm.scala 100:32]
  wire [7:0] m_7_io_a; // @[TensorGemm.scala 100:32]
  wire [7:0] m_7_io_b; // @[TensorGemm.scala 100:32]
  wire [16:0] m_7_io_y; // @[TensorGemm.scala 100:32]
  wire  m_8_clock; // @[TensorGemm.scala 100:32]
  wire [7:0] m_8_io_a; // @[TensorGemm.scala 100:32]
  wire [7:0] m_8_io_b; // @[TensorGemm.scala 100:32]
  wire [16:0] m_8_io_y; // @[TensorGemm.scala 100:32]
  wire  m_9_clock; // @[TensorGemm.scala 100:32]
  wire [7:0] m_9_io_a; // @[TensorGemm.scala 100:32]
  wire [7:0] m_9_io_b; // @[TensorGemm.scala 100:32]
  wire [16:0] m_9_io_y; // @[TensorGemm.scala 100:32]
  wire  m_10_clock; // @[TensorGemm.scala 100:32]
  wire [7:0] m_10_io_a; // @[TensorGemm.scala 100:32]
  wire [7:0] m_10_io_b; // @[TensorGemm.scala 100:32]
  wire [16:0] m_10_io_y; // @[TensorGemm.scala 100:32]
  wire  m_11_clock; // @[TensorGemm.scala 100:32]
  wire [7:0] m_11_io_a; // @[TensorGemm.scala 100:32]
  wire [7:0] m_11_io_b; // @[TensorGemm.scala 100:32]
  wire [16:0] m_11_io_y; // @[TensorGemm.scala 100:32]
  wire  m_12_clock; // @[TensorGemm.scala 100:32]
  wire [7:0] m_12_io_a; // @[TensorGemm.scala 100:32]
  wire [7:0] m_12_io_b; // @[TensorGemm.scala 100:32]
  wire [16:0] m_12_io_y; // @[TensorGemm.scala 100:32]
  wire  m_13_clock; // @[TensorGemm.scala 100:32]
  wire [7:0] m_13_io_a; // @[TensorGemm.scala 100:32]
  wire [7:0] m_13_io_b; // @[TensorGemm.scala 100:32]
  wire [16:0] m_13_io_y; // @[TensorGemm.scala 100:32]
  wire  m_14_clock; // @[TensorGemm.scala 100:32]
  wire [7:0] m_14_io_a; // @[TensorGemm.scala 100:32]
  wire [7:0] m_14_io_b; // @[TensorGemm.scala 100:32]
  wire [16:0] m_14_io_y; // @[TensorGemm.scala 100:32]
  wire  m_15_clock; // @[TensorGemm.scala 100:32]
  wire [7:0] m_15_io_a; // @[TensorGemm.scala 100:32]
  wire [7:0] m_15_io_b; // @[TensorGemm.scala 100:32]
  wire [16:0] m_15_io_y; // @[TensorGemm.scala 100:32]
  wire [16:0] a_0_0_io_a; // @[TensorGemm.scala 108:17]
  wire [16:0] a_0_0_io_b; // @[TensorGemm.scala 108:17]
  wire [17:0] a_0_0_io_y; // @[TensorGemm.scala 108:17]
  wire [16:0] a_0_1_io_a; // @[TensorGemm.scala 108:17]
  wire [16:0] a_0_1_io_b; // @[TensorGemm.scala 108:17]
  wire [17:0] a_0_1_io_y; // @[TensorGemm.scala 108:17]
  wire [16:0] a_0_2_io_a; // @[TensorGemm.scala 108:17]
  wire [16:0] a_0_2_io_b; // @[TensorGemm.scala 108:17]
  wire [17:0] a_0_2_io_y; // @[TensorGemm.scala 108:17]
  wire [16:0] a_0_3_io_a; // @[TensorGemm.scala 108:17]
  wire [16:0] a_0_3_io_b; // @[TensorGemm.scala 108:17]
  wire [17:0] a_0_3_io_y; // @[TensorGemm.scala 108:17]
  wire [16:0] a_0_4_io_a; // @[TensorGemm.scala 108:17]
  wire [16:0] a_0_4_io_b; // @[TensorGemm.scala 108:17]
  wire [17:0] a_0_4_io_y; // @[TensorGemm.scala 108:17]
  wire [16:0] a_0_5_io_a; // @[TensorGemm.scala 108:17]
  wire [16:0] a_0_5_io_b; // @[TensorGemm.scala 108:17]
  wire [17:0] a_0_5_io_y; // @[TensorGemm.scala 108:17]
  wire [16:0] a_0_6_io_a; // @[TensorGemm.scala 108:17]
  wire [16:0] a_0_6_io_b; // @[TensorGemm.scala 108:17]
  wire [17:0] a_0_6_io_y; // @[TensorGemm.scala 108:17]
  wire [16:0] a_0_7_io_a; // @[TensorGemm.scala 108:17]
  wire [16:0] a_0_7_io_b; // @[TensorGemm.scala 108:17]
  wire [17:0] a_0_7_io_y; // @[TensorGemm.scala 108:17]
  wire [17:0] a_1_0_io_a; // @[TensorGemm.scala 108:17]
  wire [17:0] a_1_0_io_b; // @[TensorGemm.scala 108:17]
  wire [18:0] a_1_0_io_y; // @[TensorGemm.scala 108:17]
  wire [17:0] a_1_1_io_a; // @[TensorGemm.scala 108:17]
  wire [17:0] a_1_1_io_b; // @[TensorGemm.scala 108:17]
  wire [18:0] a_1_1_io_y; // @[TensorGemm.scala 108:17]
  wire [17:0] a_1_2_io_a; // @[TensorGemm.scala 108:17]
  wire [17:0] a_1_2_io_b; // @[TensorGemm.scala 108:17]
  wire [18:0] a_1_2_io_y; // @[TensorGemm.scala 108:17]
  wire [17:0] a_1_3_io_a; // @[TensorGemm.scala 108:17]
  wire [17:0] a_1_3_io_b; // @[TensorGemm.scala 108:17]
  wire [18:0] a_1_3_io_y; // @[TensorGemm.scala 108:17]
  wire  a_2_0_clock; // @[TensorGemm.scala 105:17]
  wire [18:0] a_2_0_io_a; // @[TensorGemm.scala 105:17]
  wire [18:0] a_2_0_io_b; // @[TensorGemm.scala 105:17]
  wire [19:0] a_2_0_io_y; // @[TensorGemm.scala 105:17]
  wire  a_2_1_clock; // @[TensorGemm.scala 105:17]
  wire [18:0] a_2_1_io_a; // @[TensorGemm.scala 105:17]
  wire [18:0] a_2_1_io_b; // @[TensorGemm.scala 105:17]
  wire [19:0] a_2_1_io_y; // @[TensorGemm.scala 105:17]
  wire [19:0] a_3_0_io_a; // @[TensorGemm.scala 108:17]
  wire [19:0] a_3_0_io_b; // @[TensorGemm.scala 108:17]
  wire [20:0] a_3_0_io_y; // @[TensorGemm.scala 108:17]
  MAC m_0 ( // @[TensorGemm.scala 100:32]
    .clock(m_0_clock),
    .io_a(m_0_io_a),
    .io_b(m_0_io_b),
    .io_y(m_0_io_y)
  );
  MAC m_1 ( // @[TensorGemm.scala 100:32]
    .clock(m_1_clock),
    .io_a(m_1_io_a),
    .io_b(m_1_io_b),
    .io_y(m_1_io_y)
  );
  MAC m_2 ( // @[TensorGemm.scala 100:32]
    .clock(m_2_clock),
    .io_a(m_2_io_a),
    .io_b(m_2_io_b),
    .io_y(m_2_io_y)
  );
  MAC m_3 ( // @[TensorGemm.scala 100:32]
    .clock(m_3_clock),
    .io_a(m_3_io_a),
    .io_b(m_3_io_b),
    .io_y(m_3_io_y)
  );
  MAC m_4 ( // @[TensorGemm.scala 100:32]
    .clock(m_4_clock),
    .io_a(m_4_io_a),
    .io_b(m_4_io_b),
    .io_y(m_4_io_y)
  );
  MAC m_5 ( // @[TensorGemm.scala 100:32]
    .clock(m_5_clock),
    .io_a(m_5_io_a),
    .io_b(m_5_io_b),
    .io_y(m_5_io_y)
  );
  MAC m_6 ( // @[TensorGemm.scala 100:32]
    .clock(m_6_clock),
    .io_a(m_6_io_a),
    .io_b(m_6_io_b),
    .io_y(m_6_io_y)
  );
  MAC m_7 ( // @[TensorGemm.scala 100:32]
    .clock(m_7_clock),
    .io_a(m_7_io_a),
    .io_b(m_7_io_b),
    .io_y(m_7_io_y)
  );
  MAC m_8 ( // @[TensorGemm.scala 100:32]
    .clock(m_8_clock),
    .io_a(m_8_io_a),
    .io_b(m_8_io_b),
    .io_y(m_8_io_y)
  );
  MAC m_9 ( // @[TensorGemm.scala 100:32]
    .clock(m_9_clock),
    .io_a(m_9_io_a),
    .io_b(m_9_io_b),
    .io_y(m_9_io_y)
  );
  MAC m_10 ( // @[TensorGemm.scala 100:32]
    .clock(m_10_clock),
    .io_a(m_10_io_a),
    .io_b(m_10_io_b),
    .io_y(m_10_io_y)
  );
  MAC m_11 ( // @[TensorGemm.scala 100:32]
    .clock(m_11_clock),
    .io_a(m_11_io_a),
    .io_b(m_11_io_b),
    .io_y(m_11_io_y)
  );
  MAC m_12 ( // @[TensorGemm.scala 100:32]
    .clock(m_12_clock),
    .io_a(m_12_io_a),
    .io_b(m_12_io_b),
    .io_y(m_12_io_y)
  );
  MAC m_13 ( // @[TensorGemm.scala 100:32]
    .clock(m_13_clock),
    .io_a(m_13_io_a),
    .io_b(m_13_io_b),
    .io_y(m_13_io_y)
  );
  MAC m_14 ( // @[TensorGemm.scala 100:32]
    .clock(m_14_clock),
    .io_a(m_14_io_a),
    .io_b(m_14_io_b),
    .io_y(m_14_io_y)
  );
  MAC m_15 ( // @[TensorGemm.scala 100:32]
    .clock(m_15_clock),
    .io_a(m_15_io_a),
    .io_b(m_15_io_b),
    .io_y(m_15_io_y)
  );
  Adder a_0_0 ( // @[TensorGemm.scala 108:17]
    .io_a(a_0_0_io_a),
    .io_b(a_0_0_io_b),
    .io_y(a_0_0_io_y)
  );
  Adder a_0_1 ( // @[TensorGemm.scala 108:17]
    .io_a(a_0_1_io_a),
    .io_b(a_0_1_io_b),
    .io_y(a_0_1_io_y)
  );
  Adder a_0_2 ( // @[TensorGemm.scala 108:17]
    .io_a(a_0_2_io_a),
    .io_b(a_0_2_io_b),
    .io_y(a_0_2_io_y)
  );
  Adder a_0_3 ( // @[TensorGemm.scala 108:17]
    .io_a(a_0_3_io_a),
    .io_b(a_0_3_io_b),
    .io_y(a_0_3_io_y)
  );
  Adder a_0_4 ( // @[TensorGemm.scala 108:17]
    .io_a(a_0_4_io_a),
    .io_b(a_0_4_io_b),
    .io_y(a_0_4_io_y)
  );
  Adder a_0_5 ( // @[TensorGemm.scala 108:17]
    .io_a(a_0_5_io_a),
    .io_b(a_0_5_io_b),
    .io_y(a_0_5_io_y)
  );
  Adder a_0_6 ( // @[TensorGemm.scala 108:17]
    .io_a(a_0_6_io_a),
    .io_b(a_0_6_io_b),
    .io_y(a_0_6_io_y)
  );
  Adder a_0_7 ( // @[TensorGemm.scala 108:17]
    .io_a(a_0_7_io_a),
    .io_b(a_0_7_io_b),
    .io_y(a_0_7_io_y)
  );
  Adder_8 a_1_0 ( // @[TensorGemm.scala 108:17]
    .io_a(a_1_0_io_a),
    .io_b(a_1_0_io_b),
    .io_y(a_1_0_io_y)
  );
  Adder_8 a_1_1 ( // @[TensorGemm.scala 108:17]
    .io_a(a_1_1_io_a),
    .io_b(a_1_1_io_b),
    .io_y(a_1_1_io_y)
  );
  Adder_8 a_1_2 ( // @[TensorGemm.scala 108:17]
    .io_a(a_1_2_io_a),
    .io_b(a_1_2_io_b),
    .io_y(a_1_2_io_y)
  );
  Adder_8 a_1_3 ( // @[TensorGemm.scala 108:17]
    .io_a(a_1_3_io_a),
    .io_b(a_1_3_io_b),
    .io_y(a_1_3_io_y)
  );
  PipeAdder a_2_0 ( // @[TensorGemm.scala 105:17]
    .clock(a_2_0_clock),
    .io_a(a_2_0_io_a),
    .io_b(a_2_0_io_b),
    .io_y(a_2_0_io_y)
  );
  PipeAdder a_2_1 ( // @[TensorGemm.scala 105:17]
    .clock(a_2_1_clock),
    .io_a(a_2_1_io_a),
    .io_b(a_2_1_io_b),
    .io_y(a_2_1_io_y)
  );
  Adder_12 a_3_0 ( // @[TensorGemm.scala 108:17]
    .io_a(a_3_0_io_a),
    .io_b(a_3_0_io_b),
    .io_y(a_3_0_io_y)
  );
  assign io_y = a_3_0_io_y; // @[TensorGemm.scala 134:8]
  assign m_0_clock = clock;
  assign m_0_io_a = io_a_0; // @[TensorGemm.scala 114:15]
  assign m_0_io_b = io_b_0; // @[TensorGemm.scala 115:15]
  assign m_1_clock = clock;
  assign m_1_io_a = io_a_1; // @[TensorGemm.scala 114:15]
  assign m_1_io_b = io_b_1; // @[TensorGemm.scala 115:15]
  assign m_2_clock = clock;
  assign m_2_io_a = io_a_2; // @[TensorGemm.scala 114:15]
  assign m_2_io_b = io_b_2; // @[TensorGemm.scala 115:15]
  assign m_3_clock = clock;
  assign m_3_io_a = io_a_3; // @[TensorGemm.scala 114:15]
  assign m_3_io_b = io_b_3; // @[TensorGemm.scala 115:15]
  assign m_4_clock = clock;
  assign m_4_io_a = io_a_4; // @[TensorGemm.scala 114:15]
  assign m_4_io_b = io_b_4; // @[TensorGemm.scala 115:15]
  assign m_5_clock = clock;
  assign m_5_io_a = io_a_5; // @[TensorGemm.scala 114:15]
  assign m_5_io_b = io_b_5; // @[TensorGemm.scala 115:15]
  assign m_6_clock = clock;
  assign m_6_io_a = io_a_6; // @[TensorGemm.scala 114:15]
  assign m_6_io_b = io_b_6; // @[TensorGemm.scala 115:15]
  assign m_7_clock = clock;
  assign m_7_io_a = io_a_7; // @[TensorGemm.scala 114:15]
  assign m_7_io_b = io_b_7; // @[TensorGemm.scala 115:15]
  assign m_8_clock = clock;
  assign m_8_io_a = io_a_8; // @[TensorGemm.scala 114:15]
  assign m_8_io_b = io_b_8; // @[TensorGemm.scala 115:15]
  assign m_9_clock = clock;
  assign m_9_io_a = io_a_9; // @[TensorGemm.scala 114:15]
  assign m_9_io_b = io_b_9; // @[TensorGemm.scala 115:15]
  assign m_10_clock = clock;
  assign m_10_io_a = io_a_10; // @[TensorGemm.scala 114:15]
  assign m_10_io_b = io_b_10; // @[TensorGemm.scala 115:15]
  assign m_11_clock = clock;
  assign m_11_io_a = io_a_11; // @[TensorGemm.scala 114:15]
  assign m_11_io_b = io_b_11; // @[TensorGemm.scala 115:15]
  assign m_12_clock = clock;
  assign m_12_io_a = io_a_12; // @[TensorGemm.scala 114:15]
  assign m_12_io_b = io_b_12; // @[TensorGemm.scala 115:15]
  assign m_13_clock = clock;
  assign m_13_io_a = io_a_13; // @[TensorGemm.scala 114:15]
  assign m_13_io_b = io_b_13; // @[TensorGemm.scala 115:15]
  assign m_14_clock = clock;
  assign m_14_io_a = io_a_14; // @[TensorGemm.scala 114:15]
  assign m_14_io_b = io_b_14; // @[TensorGemm.scala 115:15]
  assign m_15_clock = clock;
  assign m_15_io_a = io_a_15; // @[TensorGemm.scala 114:15]
  assign m_15_io_b = io_b_15; // @[TensorGemm.scala 115:15]
  assign a_0_0_io_a = m_0_io_y; // @[TensorGemm.scala 124:22]
  assign a_0_0_io_b = m_1_io_y; // @[TensorGemm.scala 125:22]
  assign a_0_1_io_a = m_2_io_y; // @[TensorGemm.scala 124:22]
  assign a_0_1_io_b = m_3_io_y; // @[TensorGemm.scala 125:22]
  assign a_0_2_io_a = m_4_io_y; // @[TensorGemm.scala 124:22]
  assign a_0_2_io_b = m_5_io_y; // @[TensorGemm.scala 125:22]
  assign a_0_3_io_a = m_6_io_y; // @[TensorGemm.scala 124:22]
  assign a_0_3_io_b = m_7_io_y; // @[TensorGemm.scala 125:22]
  assign a_0_4_io_a = m_8_io_y; // @[TensorGemm.scala 124:22]
  assign a_0_4_io_b = m_9_io_y; // @[TensorGemm.scala 125:22]
  assign a_0_5_io_a = m_10_io_y; // @[TensorGemm.scala 124:22]
  assign a_0_5_io_b = m_11_io_y; // @[TensorGemm.scala 125:22]
  assign a_0_6_io_a = m_12_io_y; // @[TensorGemm.scala 124:22]
  assign a_0_6_io_b = m_13_io_y; // @[TensorGemm.scala 125:22]
  assign a_0_7_io_a = m_14_io_y; // @[TensorGemm.scala 124:22]
  assign a_0_7_io_b = m_15_io_y; // @[TensorGemm.scala 125:22]
  assign a_1_0_io_a = a_0_0_io_y; // @[TensorGemm.scala 127:22]
  assign a_1_0_io_b = a_0_1_io_y; // @[TensorGemm.scala 128:22]
  assign a_1_1_io_a = a_0_2_io_y; // @[TensorGemm.scala 127:22]
  assign a_1_1_io_b = a_0_3_io_y; // @[TensorGemm.scala 128:22]
  assign a_1_2_io_a = a_0_4_io_y; // @[TensorGemm.scala 127:22]
  assign a_1_2_io_b = a_0_5_io_y; // @[TensorGemm.scala 128:22]
  assign a_1_3_io_a = a_0_6_io_y; // @[TensorGemm.scala 127:22]
  assign a_1_3_io_b = a_0_7_io_y; // @[TensorGemm.scala 128:22]
  assign a_2_0_clock = clock;
  assign a_2_0_io_a = a_1_0_io_y; // @[TensorGemm.scala 127:22]
  assign a_2_0_io_b = a_1_1_io_y; // @[TensorGemm.scala 128:22]
  assign a_2_1_clock = clock;
  assign a_2_1_io_a = a_1_2_io_y; // @[TensorGemm.scala 127:22]
  assign a_2_1_io_b = a_1_3_io_y; // @[TensorGemm.scala 128:22]
  assign a_3_0_io_a = a_2_0_io_y; // @[TensorGemm.scala 127:22]
  assign a_3_0_io_b = a_2_1_io_y; // @[TensorGemm.scala 128:22]
endmodule
module MatrixVectorMultiplicationBypass(
  input         clock,
  input         io_valid_reset,
  input  [7:0]  io_inp_data_bits_0_0,
  input  [7:0]  io_inp_data_bits_0_1,
  input  [7:0]  io_inp_data_bits_0_2,
  input  [7:0]  io_inp_data_bits_0_3,
  input  [7:0]  io_inp_data_bits_0_4,
  input  [7:0]  io_inp_data_bits_0_5,
  input  [7:0]  io_inp_data_bits_0_6,
  input  [7:0]  io_inp_data_bits_0_7,
  input  [7:0]  io_inp_data_bits_0_8,
  input  [7:0]  io_inp_data_bits_0_9,
  input  [7:0]  io_inp_data_bits_0_10,
  input  [7:0]  io_inp_data_bits_0_11,
  input  [7:0]  io_inp_data_bits_0_12,
  input  [7:0]  io_inp_data_bits_0_13,
  input  [7:0]  io_inp_data_bits_0_14,
  input  [7:0]  io_inp_data_bits_0_15,
  input  [7:0]  io_wgt_data_bits_0_0,
  input  [7:0]  io_wgt_data_bits_0_1,
  input  [7:0]  io_wgt_data_bits_0_2,
  input  [7:0]  io_wgt_data_bits_0_3,
  input  [7:0]  io_wgt_data_bits_0_4,
  input  [7:0]  io_wgt_data_bits_0_5,
  input  [7:0]  io_wgt_data_bits_0_6,
  input  [7:0]  io_wgt_data_bits_0_7,
  input  [7:0]  io_wgt_data_bits_0_8,
  input  [7:0]  io_wgt_data_bits_0_9,
  input  [7:0]  io_wgt_data_bits_0_10,
  input  [7:0]  io_wgt_data_bits_0_11,
  input  [7:0]  io_wgt_data_bits_0_12,
  input  [7:0]  io_wgt_data_bits_0_13,
  input  [7:0]  io_wgt_data_bits_0_14,
  input  [7:0]  io_wgt_data_bits_0_15,
  input  [7:0]  io_wgt_data_bits_1_0,
  input  [7:0]  io_wgt_data_bits_1_1,
  input  [7:0]  io_wgt_data_bits_1_2,
  input  [7:0]  io_wgt_data_bits_1_3,
  input  [7:0]  io_wgt_data_bits_1_4,
  input  [7:0]  io_wgt_data_bits_1_5,
  input  [7:0]  io_wgt_data_bits_1_6,
  input  [7:0]  io_wgt_data_bits_1_7,
  input  [7:0]  io_wgt_data_bits_1_8,
  input  [7:0]  io_wgt_data_bits_1_9,
  input  [7:0]  io_wgt_data_bits_1_10,
  input  [7:0]  io_wgt_data_bits_1_11,
  input  [7:0]  io_wgt_data_bits_1_12,
  input  [7:0]  io_wgt_data_bits_1_13,
  input  [7:0]  io_wgt_data_bits_1_14,
  input  [7:0]  io_wgt_data_bits_1_15,
  input  [7:0]  io_wgt_data_bits_2_0,
  input  [7:0]  io_wgt_data_bits_2_1,
  input  [7:0]  io_wgt_data_bits_2_2,
  input  [7:0]  io_wgt_data_bits_2_3,
  input  [7:0]  io_wgt_data_bits_2_4,
  input  [7:0]  io_wgt_data_bits_2_5,
  input  [7:0]  io_wgt_data_bits_2_6,
  input  [7:0]  io_wgt_data_bits_2_7,
  input  [7:0]  io_wgt_data_bits_2_8,
  input  [7:0]  io_wgt_data_bits_2_9,
  input  [7:0]  io_wgt_data_bits_2_10,
  input  [7:0]  io_wgt_data_bits_2_11,
  input  [7:0]  io_wgt_data_bits_2_12,
  input  [7:0]  io_wgt_data_bits_2_13,
  input  [7:0]  io_wgt_data_bits_2_14,
  input  [7:0]  io_wgt_data_bits_2_15,
  input  [7:0]  io_wgt_data_bits_3_0,
  input  [7:0]  io_wgt_data_bits_3_1,
  input  [7:0]  io_wgt_data_bits_3_2,
  input  [7:0]  io_wgt_data_bits_3_3,
  input  [7:0]  io_wgt_data_bits_3_4,
  input  [7:0]  io_wgt_data_bits_3_5,
  input  [7:0]  io_wgt_data_bits_3_6,
  input  [7:0]  io_wgt_data_bits_3_7,
  input  [7:0]  io_wgt_data_bits_3_8,
  input  [7:0]  io_wgt_data_bits_3_9,
  input  [7:0]  io_wgt_data_bits_3_10,
  input  [7:0]  io_wgt_data_bits_3_11,
  input  [7:0]  io_wgt_data_bits_3_12,
  input  [7:0]  io_wgt_data_bits_3_13,
  input  [7:0]  io_wgt_data_bits_3_14,
  input  [7:0]  io_wgt_data_bits_3_15,
  input  [7:0]  io_wgt_data_bits_4_0,
  input  [7:0]  io_wgt_data_bits_4_1,
  input  [7:0]  io_wgt_data_bits_4_2,
  input  [7:0]  io_wgt_data_bits_4_3,
  input  [7:0]  io_wgt_data_bits_4_4,
  input  [7:0]  io_wgt_data_bits_4_5,
  input  [7:0]  io_wgt_data_bits_4_6,
  input  [7:0]  io_wgt_data_bits_4_7,
  input  [7:0]  io_wgt_data_bits_4_8,
  input  [7:0]  io_wgt_data_bits_4_9,
  input  [7:0]  io_wgt_data_bits_4_10,
  input  [7:0]  io_wgt_data_bits_4_11,
  input  [7:0]  io_wgt_data_bits_4_12,
  input  [7:0]  io_wgt_data_bits_4_13,
  input  [7:0]  io_wgt_data_bits_4_14,
  input  [7:0]  io_wgt_data_bits_4_15,
  input  [7:0]  io_wgt_data_bits_5_0,
  input  [7:0]  io_wgt_data_bits_5_1,
  input  [7:0]  io_wgt_data_bits_5_2,
  input  [7:0]  io_wgt_data_bits_5_3,
  input  [7:0]  io_wgt_data_bits_5_4,
  input  [7:0]  io_wgt_data_bits_5_5,
  input  [7:0]  io_wgt_data_bits_5_6,
  input  [7:0]  io_wgt_data_bits_5_7,
  input  [7:0]  io_wgt_data_bits_5_8,
  input  [7:0]  io_wgt_data_bits_5_9,
  input  [7:0]  io_wgt_data_bits_5_10,
  input  [7:0]  io_wgt_data_bits_5_11,
  input  [7:0]  io_wgt_data_bits_5_12,
  input  [7:0]  io_wgt_data_bits_5_13,
  input  [7:0]  io_wgt_data_bits_5_14,
  input  [7:0]  io_wgt_data_bits_5_15,
  input  [7:0]  io_wgt_data_bits_6_0,
  input  [7:0]  io_wgt_data_bits_6_1,
  input  [7:0]  io_wgt_data_bits_6_2,
  input  [7:0]  io_wgt_data_bits_6_3,
  input  [7:0]  io_wgt_data_bits_6_4,
  input  [7:0]  io_wgt_data_bits_6_5,
  input  [7:0]  io_wgt_data_bits_6_6,
  input  [7:0]  io_wgt_data_bits_6_7,
  input  [7:0]  io_wgt_data_bits_6_8,
  input  [7:0]  io_wgt_data_bits_6_9,
  input  [7:0]  io_wgt_data_bits_6_10,
  input  [7:0]  io_wgt_data_bits_6_11,
  input  [7:0]  io_wgt_data_bits_6_12,
  input  [7:0]  io_wgt_data_bits_6_13,
  input  [7:0]  io_wgt_data_bits_6_14,
  input  [7:0]  io_wgt_data_bits_6_15,
  input  [7:0]  io_wgt_data_bits_7_0,
  input  [7:0]  io_wgt_data_bits_7_1,
  input  [7:0]  io_wgt_data_bits_7_2,
  input  [7:0]  io_wgt_data_bits_7_3,
  input  [7:0]  io_wgt_data_bits_7_4,
  input  [7:0]  io_wgt_data_bits_7_5,
  input  [7:0]  io_wgt_data_bits_7_6,
  input  [7:0]  io_wgt_data_bits_7_7,
  input  [7:0]  io_wgt_data_bits_7_8,
  input  [7:0]  io_wgt_data_bits_7_9,
  input  [7:0]  io_wgt_data_bits_7_10,
  input  [7:0]  io_wgt_data_bits_7_11,
  input  [7:0]  io_wgt_data_bits_7_12,
  input  [7:0]  io_wgt_data_bits_7_13,
  input  [7:0]  io_wgt_data_bits_7_14,
  input  [7:0]  io_wgt_data_bits_7_15,
  input  [7:0]  io_wgt_data_bits_8_0,
  input  [7:0]  io_wgt_data_bits_8_1,
  input  [7:0]  io_wgt_data_bits_8_2,
  input  [7:0]  io_wgt_data_bits_8_3,
  input  [7:0]  io_wgt_data_bits_8_4,
  input  [7:0]  io_wgt_data_bits_8_5,
  input  [7:0]  io_wgt_data_bits_8_6,
  input  [7:0]  io_wgt_data_bits_8_7,
  input  [7:0]  io_wgt_data_bits_8_8,
  input  [7:0]  io_wgt_data_bits_8_9,
  input  [7:0]  io_wgt_data_bits_8_10,
  input  [7:0]  io_wgt_data_bits_8_11,
  input  [7:0]  io_wgt_data_bits_8_12,
  input  [7:0]  io_wgt_data_bits_8_13,
  input  [7:0]  io_wgt_data_bits_8_14,
  input  [7:0]  io_wgt_data_bits_8_15,
  input  [7:0]  io_wgt_data_bits_9_0,
  input  [7:0]  io_wgt_data_bits_9_1,
  input  [7:0]  io_wgt_data_bits_9_2,
  input  [7:0]  io_wgt_data_bits_9_3,
  input  [7:0]  io_wgt_data_bits_9_4,
  input  [7:0]  io_wgt_data_bits_9_5,
  input  [7:0]  io_wgt_data_bits_9_6,
  input  [7:0]  io_wgt_data_bits_9_7,
  input  [7:0]  io_wgt_data_bits_9_8,
  input  [7:0]  io_wgt_data_bits_9_9,
  input  [7:0]  io_wgt_data_bits_9_10,
  input  [7:0]  io_wgt_data_bits_9_11,
  input  [7:0]  io_wgt_data_bits_9_12,
  input  [7:0]  io_wgt_data_bits_9_13,
  input  [7:0]  io_wgt_data_bits_9_14,
  input  [7:0]  io_wgt_data_bits_9_15,
  input  [7:0]  io_wgt_data_bits_10_0,
  input  [7:0]  io_wgt_data_bits_10_1,
  input  [7:0]  io_wgt_data_bits_10_2,
  input  [7:0]  io_wgt_data_bits_10_3,
  input  [7:0]  io_wgt_data_bits_10_4,
  input  [7:0]  io_wgt_data_bits_10_5,
  input  [7:0]  io_wgt_data_bits_10_6,
  input  [7:0]  io_wgt_data_bits_10_7,
  input  [7:0]  io_wgt_data_bits_10_8,
  input  [7:0]  io_wgt_data_bits_10_9,
  input  [7:0]  io_wgt_data_bits_10_10,
  input  [7:0]  io_wgt_data_bits_10_11,
  input  [7:0]  io_wgt_data_bits_10_12,
  input  [7:0]  io_wgt_data_bits_10_13,
  input  [7:0]  io_wgt_data_bits_10_14,
  input  [7:0]  io_wgt_data_bits_10_15,
  input  [7:0]  io_wgt_data_bits_11_0,
  input  [7:0]  io_wgt_data_bits_11_1,
  input  [7:0]  io_wgt_data_bits_11_2,
  input  [7:0]  io_wgt_data_bits_11_3,
  input  [7:0]  io_wgt_data_bits_11_4,
  input  [7:0]  io_wgt_data_bits_11_5,
  input  [7:0]  io_wgt_data_bits_11_6,
  input  [7:0]  io_wgt_data_bits_11_7,
  input  [7:0]  io_wgt_data_bits_11_8,
  input  [7:0]  io_wgt_data_bits_11_9,
  input  [7:0]  io_wgt_data_bits_11_10,
  input  [7:0]  io_wgt_data_bits_11_11,
  input  [7:0]  io_wgt_data_bits_11_12,
  input  [7:0]  io_wgt_data_bits_11_13,
  input  [7:0]  io_wgt_data_bits_11_14,
  input  [7:0]  io_wgt_data_bits_11_15,
  input  [7:0]  io_wgt_data_bits_12_0,
  input  [7:0]  io_wgt_data_bits_12_1,
  input  [7:0]  io_wgt_data_bits_12_2,
  input  [7:0]  io_wgt_data_bits_12_3,
  input  [7:0]  io_wgt_data_bits_12_4,
  input  [7:0]  io_wgt_data_bits_12_5,
  input  [7:0]  io_wgt_data_bits_12_6,
  input  [7:0]  io_wgt_data_bits_12_7,
  input  [7:0]  io_wgt_data_bits_12_8,
  input  [7:0]  io_wgt_data_bits_12_9,
  input  [7:0]  io_wgt_data_bits_12_10,
  input  [7:0]  io_wgt_data_bits_12_11,
  input  [7:0]  io_wgt_data_bits_12_12,
  input  [7:0]  io_wgt_data_bits_12_13,
  input  [7:0]  io_wgt_data_bits_12_14,
  input  [7:0]  io_wgt_data_bits_12_15,
  input  [7:0]  io_wgt_data_bits_13_0,
  input  [7:0]  io_wgt_data_bits_13_1,
  input  [7:0]  io_wgt_data_bits_13_2,
  input  [7:0]  io_wgt_data_bits_13_3,
  input  [7:0]  io_wgt_data_bits_13_4,
  input  [7:0]  io_wgt_data_bits_13_5,
  input  [7:0]  io_wgt_data_bits_13_6,
  input  [7:0]  io_wgt_data_bits_13_7,
  input  [7:0]  io_wgt_data_bits_13_8,
  input  [7:0]  io_wgt_data_bits_13_9,
  input  [7:0]  io_wgt_data_bits_13_10,
  input  [7:0]  io_wgt_data_bits_13_11,
  input  [7:0]  io_wgt_data_bits_13_12,
  input  [7:0]  io_wgt_data_bits_13_13,
  input  [7:0]  io_wgt_data_bits_13_14,
  input  [7:0]  io_wgt_data_bits_13_15,
  input  [7:0]  io_wgt_data_bits_14_0,
  input  [7:0]  io_wgt_data_bits_14_1,
  input  [7:0]  io_wgt_data_bits_14_2,
  input  [7:0]  io_wgt_data_bits_14_3,
  input  [7:0]  io_wgt_data_bits_14_4,
  input  [7:0]  io_wgt_data_bits_14_5,
  input  [7:0]  io_wgt_data_bits_14_6,
  input  [7:0]  io_wgt_data_bits_14_7,
  input  [7:0]  io_wgt_data_bits_14_8,
  input  [7:0]  io_wgt_data_bits_14_9,
  input  [7:0]  io_wgt_data_bits_14_10,
  input  [7:0]  io_wgt_data_bits_14_11,
  input  [7:0]  io_wgt_data_bits_14_12,
  input  [7:0]  io_wgt_data_bits_14_13,
  input  [7:0]  io_wgt_data_bits_14_14,
  input  [7:0]  io_wgt_data_bits_14_15,
  input  [7:0]  io_wgt_data_bits_15_0,
  input  [7:0]  io_wgt_data_bits_15_1,
  input  [7:0]  io_wgt_data_bits_15_2,
  input  [7:0]  io_wgt_data_bits_15_3,
  input  [7:0]  io_wgt_data_bits_15_4,
  input  [7:0]  io_wgt_data_bits_15_5,
  input  [7:0]  io_wgt_data_bits_15_6,
  input  [7:0]  io_wgt_data_bits_15_7,
  input  [7:0]  io_wgt_data_bits_15_8,
  input  [7:0]  io_wgt_data_bits_15_9,
  input  [7:0]  io_wgt_data_bits_15_10,
  input  [7:0]  io_wgt_data_bits_15_11,
  input  [7:0]  io_wgt_data_bits_15_12,
  input  [7:0]  io_wgt_data_bits_15_13,
  input  [7:0]  io_wgt_data_bits_15_14,
  input  [7:0]  io_wgt_data_bits_15_15,
  input  [7:0]  io_wgt_data_bits_16_0,
  input  [7:0]  io_wgt_data_bits_16_1,
  input  [7:0]  io_wgt_data_bits_16_2,
  input  [7:0]  io_wgt_data_bits_16_3,
  input  [7:0]  io_wgt_data_bits_16_4,
  input  [7:0]  io_wgt_data_bits_16_5,
  input  [7:0]  io_wgt_data_bits_16_6,
  input  [7:0]  io_wgt_data_bits_16_7,
  input  [7:0]  io_wgt_data_bits_16_8,
  input  [7:0]  io_wgt_data_bits_16_9,
  input  [7:0]  io_wgt_data_bits_16_10,
  input  [7:0]  io_wgt_data_bits_16_11,
  input  [7:0]  io_wgt_data_bits_16_12,
  input  [7:0]  io_wgt_data_bits_16_13,
  input  [7:0]  io_wgt_data_bits_16_14,
  input  [7:0]  io_wgt_data_bits_16_15,
  input  [7:0]  io_wgt_data_bits_17_0,
  input  [7:0]  io_wgt_data_bits_17_1,
  input  [7:0]  io_wgt_data_bits_17_2,
  input  [7:0]  io_wgt_data_bits_17_3,
  input  [7:0]  io_wgt_data_bits_17_4,
  input  [7:0]  io_wgt_data_bits_17_5,
  input  [7:0]  io_wgt_data_bits_17_6,
  input  [7:0]  io_wgt_data_bits_17_7,
  input  [7:0]  io_wgt_data_bits_17_8,
  input  [7:0]  io_wgt_data_bits_17_9,
  input  [7:0]  io_wgt_data_bits_17_10,
  input  [7:0]  io_wgt_data_bits_17_11,
  input  [7:0]  io_wgt_data_bits_17_12,
  input  [7:0]  io_wgt_data_bits_17_13,
  input  [7:0]  io_wgt_data_bits_17_14,
  input  [7:0]  io_wgt_data_bits_17_15,
  input  [7:0]  io_wgt_data_bits_18_0,
  input  [7:0]  io_wgt_data_bits_18_1,
  input  [7:0]  io_wgt_data_bits_18_2,
  input  [7:0]  io_wgt_data_bits_18_3,
  input  [7:0]  io_wgt_data_bits_18_4,
  input  [7:0]  io_wgt_data_bits_18_5,
  input  [7:0]  io_wgt_data_bits_18_6,
  input  [7:0]  io_wgt_data_bits_18_7,
  input  [7:0]  io_wgt_data_bits_18_8,
  input  [7:0]  io_wgt_data_bits_18_9,
  input  [7:0]  io_wgt_data_bits_18_10,
  input  [7:0]  io_wgt_data_bits_18_11,
  input  [7:0]  io_wgt_data_bits_18_12,
  input  [7:0]  io_wgt_data_bits_18_13,
  input  [7:0]  io_wgt_data_bits_18_14,
  input  [7:0]  io_wgt_data_bits_18_15,
  input  [7:0]  io_wgt_data_bits_19_0,
  input  [7:0]  io_wgt_data_bits_19_1,
  input  [7:0]  io_wgt_data_bits_19_2,
  input  [7:0]  io_wgt_data_bits_19_3,
  input  [7:0]  io_wgt_data_bits_19_4,
  input  [7:0]  io_wgt_data_bits_19_5,
  input  [7:0]  io_wgt_data_bits_19_6,
  input  [7:0]  io_wgt_data_bits_19_7,
  input  [7:0]  io_wgt_data_bits_19_8,
  input  [7:0]  io_wgt_data_bits_19_9,
  input  [7:0]  io_wgt_data_bits_19_10,
  input  [7:0]  io_wgt_data_bits_19_11,
  input  [7:0]  io_wgt_data_bits_19_12,
  input  [7:0]  io_wgt_data_bits_19_13,
  input  [7:0]  io_wgt_data_bits_19_14,
  input  [7:0]  io_wgt_data_bits_19_15,
  input  [7:0]  io_wgt_data_bits_20_0,
  input  [7:0]  io_wgt_data_bits_20_1,
  input  [7:0]  io_wgt_data_bits_20_2,
  input  [7:0]  io_wgt_data_bits_20_3,
  input  [7:0]  io_wgt_data_bits_20_4,
  input  [7:0]  io_wgt_data_bits_20_5,
  input  [7:0]  io_wgt_data_bits_20_6,
  input  [7:0]  io_wgt_data_bits_20_7,
  input  [7:0]  io_wgt_data_bits_20_8,
  input  [7:0]  io_wgt_data_bits_20_9,
  input  [7:0]  io_wgt_data_bits_20_10,
  input  [7:0]  io_wgt_data_bits_20_11,
  input  [7:0]  io_wgt_data_bits_20_12,
  input  [7:0]  io_wgt_data_bits_20_13,
  input  [7:0]  io_wgt_data_bits_20_14,
  input  [7:0]  io_wgt_data_bits_20_15,
  input  [7:0]  io_wgt_data_bits_21_0,
  input  [7:0]  io_wgt_data_bits_21_1,
  input  [7:0]  io_wgt_data_bits_21_2,
  input  [7:0]  io_wgt_data_bits_21_3,
  input  [7:0]  io_wgt_data_bits_21_4,
  input  [7:0]  io_wgt_data_bits_21_5,
  input  [7:0]  io_wgt_data_bits_21_6,
  input  [7:0]  io_wgt_data_bits_21_7,
  input  [7:0]  io_wgt_data_bits_21_8,
  input  [7:0]  io_wgt_data_bits_21_9,
  input  [7:0]  io_wgt_data_bits_21_10,
  input  [7:0]  io_wgt_data_bits_21_11,
  input  [7:0]  io_wgt_data_bits_21_12,
  input  [7:0]  io_wgt_data_bits_21_13,
  input  [7:0]  io_wgt_data_bits_21_14,
  input  [7:0]  io_wgt_data_bits_21_15,
  input  [7:0]  io_wgt_data_bits_22_0,
  input  [7:0]  io_wgt_data_bits_22_1,
  input  [7:0]  io_wgt_data_bits_22_2,
  input  [7:0]  io_wgt_data_bits_22_3,
  input  [7:0]  io_wgt_data_bits_22_4,
  input  [7:0]  io_wgt_data_bits_22_5,
  input  [7:0]  io_wgt_data_bits_22_6,
  input  [7:0]  io_wgt_data_bits_22_7,
  input  [7:0]  io_wgt_data_bits_22_8,
  input  [7:0]  io_wgt_data_bits_22_9,
  input  [7:0]  io_wgt_data_bits_22_10,
  input  [7:0]  io_wgt_data_bits_22_11,
  input  [7:0]  io_wgt_data_bits_22_12,
  input  [7:0]  io_wgt_data_bits_22_13,
  input  [7:0]  io_wgt_data_bits_22_14,
  input  [7:0]  io_wgt_data_bits_22_15,
  input  [7:0]  io_wgt_data_bits_23_0,
  input  [7:0]  io_wgt_data_bits_23_1,
  input  [7:0]  io_wgt_data_bits_23_2,
  input  [7:0]  io_wgt_data_bits_23_3,
  input  [7:0]  io_wgt_data_bits_23_4,
  input  [7:0]  io_wgt_data_bits_23_5,
  input  [7:0]  io_wgt_data_bits_23_6,
  input  [7:0]  io_wgt_data_bits_23_7,
  input  [7:0]  io_wgt_data_bits_23_8,
  input  [7:0]  io_wgt_data_bits_23_9,
  input  [7:0]  io_wgt_data_bits_23_10,
  input  [7:0]  io_wgt_data_bits_23_11,
  input  [7:0]  io_wgt_data_bits_23_12,
  input  [7:0]  io_wgt_data_bits_23_13,
  input  [7:0]  io_wgt_data_bits_23_14,
  input  [7:0]  io_wgt_data_bits_23_15,
  input  [7:0]  io_wgt_data_bits_24_0,
  input  [7:0]  io_wgt_data_bits_24_1,
  input  [7:0]  io_wgt_data_bits_24_2,
  input  [7:0]  io_wgt_data_bits_24_3,
  input  [7:0]  io_wgt_data_bits_24_4,
  input  [7:0]  io_wgt_data_bits_24_5,
  input  [7:0]  io_wgt_data_bits_24_6,
  input  [7:0]  io_wgt_data_bits_24_7,
  input  [7:0]  io_wgt_data_bits_24_8,
  input  [7:0]  io_wgt_data_bits_24_9,
  input  [7:0]  io_wgt_data_bits_24_10,
  input  [7:0]  io_wgt_data_bits_24_11,
  input  [7:0]  io_wgt_data_bits_24_12,
  input  [7:0]  io_wgt_data_bits_24_13,
  input  [7:0]  io_wgt_data_bits_24_14,
  input  [7:0]  io_wgt_data_bits_24_15,
  input  [7:0]  io_wgt_data_bits_25_0,
  input  [7:0]  io_wgt_data_bits_25_1,
  input  [7:0]  io_wgt_data_bits_25_2,
  input  [7:0]  io_wgt_data_bits_25_3,
  input  [7:0]  io_wgt_data_bits_25_4,
  input  [7:0]  io_wgt_data_bits_25_5,
  input  [7:0]  io_wgt_data_bits_25_6,
  input  [7:0]  io_wgt_data_bits_25_7,
  input  [7:0]  io_wgt_data_bits_25_8,
  input  [7:0]  io_wgt_data_bits_25_9,
  input  [7:0]  io_wgt_data_bits_25_10,
  input  [7:0]  io_wgt_data_bits_25_11,
  input  [7:0]  io_wgt_data_bits_25_12,
  input  [7:0]  io_wgt_data_bits_25_13,
  input  [7:0]  io_wgt_data_bits_25_14,
  input  [7:0]  io_wgt_data_bits_25_15,
  input  [7:0]  io_wgt_data_bits_26_0,
  input  [7:0]  io_wgt_data_bits_26_1,
  input  [7:0]  io_wgt_data_bits_26_2,
  input  [7:0]  io_wgt_data_bits_26_3,
  input  [7:0]  io_wgt_data_bits_26_4,
  input  [7:0]  io_wgt_data_bits_26_5,
  input  [7:0]  io_wgt_data_bits_26_6,
  input  [7:0]  io_wgt_data_bits_26_7,
  input  [7:0]  io_wgt_data_bits_26_8,
  input  [7:0]  io_wgt_data_bits_26_9,
  input  [7:0]  io_wgt_data_bits_26_10,
  input  [7:0]  io_wgt_data_bits_26_11,
  input  [7:0]  io_wgt_data_bits_26_12,
  input  [7:0]  io_wgt_data_bits_26_13,
  input  [7:0]  io_wgt_data_bits_26_14,
  input  [7:0]  io_wgt_data_bits_26_15,
  input  [7:0]  io_wgt_data_bits_27_0,
  input  [7:0]  io_wgt_data_bits_27_1,
  input  [7:0]  io_wgt_data_bits_27_2,
  input  [7:0]  io_wgt_data_bits_27_3,
  input  [7:0]  io_wgt_data_bits_27_4,
  input  [7:0]  io_wgt_data_bits_27_5,
  input  [7:0]  io_wgt_data_bits_27_6,
  input  [7:0]  io_wgt_data_bits_27_7,
  input  [7:0]  io_wgt_data_bits_27_8,
  input  [7:0]  io_wgt_data_bits_27_9,
  input  [7:0]  io_wgt_data_bits_27_10,
  input  [7:0]  io_wgt_data_bits_27_11,
  input  [7:0]  io_wgt_data_bits_27_12,
  input  [7:0]  io_wgt_data_bits_27_13,
  input  [7:0]  io_wgt_data_bits_27_14,
  input  [7:0]  io_wgt_data_bits_27_15,
  input  [7:0]  io_wgt_data_bits_28_0,
  input  [7:0]  io_wgt_data_bits_28_1,
  input  [7:0]  io_wgt_data_bits_28_2,
  input  [7:0]  io_wgt_data_bits_28_3,
  input  [7:0]  io_wgt_data_bits_28_4,
  input  [7:0]  io_wgt_data_bits_28_5,
  input  [7:0]  io_wgt_data_bits_28_6,
  input  [7:0]  io_wgt_data_bits_28_7,
  input  [7:0]  io_wgt_data_bits_28_8,
  input  [7:0]  io_wgt_data_bits_28_9,
  input  [7:0]  io_wgt_data_bits_28_10,
  input  [7:0]  io_wgt_data_bits_28_11,
  input  [7:0]  io_wgt_data_bits_28_12,
  input  [7:0]  io_wgt_data_bits_28_13,
  input  [7:0]  io_wgt_data_bits_28_14,
  input  [7:0]  io_wgt_data_bits_28_15,
  input  [7:0]  io_wgt_data_bits_29_0,
  input  [7:0]  io_wgt_data_bits_29_1,
  input  [7:0]  io_wgt_data_bits_29_2,
  input  [7:0]  io_wgt_data_bits_29_3,
  input  [7:0]  io_wgt_data_bits_29_4,
  input  [7:0]  io_wgt_data_bits_29_5,
  input  [7:0]  io_wgt_data_bits_29_6,
  input  [7:0]  io_wgt_data_bits_29_7,
  input  [7:0]  io_wgt_data_bits_29_8,
  input  [7:0]  io_wgt_data_bits_29_9,
  input  [7:0]  io_wgt_data_bits_29_10,
  input  [7:0]  io_wgt_data_bits_29_11,
  input  [7:0]  io_wgt_data_bits_29_12,
  input  [7:0]  io_wgt_data_bits_29_13,
  input  [7:0]  io_wgt_data_bits_29_14,
  input  [7:0]  io_wgt_data_bits_29_15,
  input  [7:0]  io_wgt_data_bits_30_0,
  input  [7:0]  io_wgt_data_bits_30_1,
  input  [7:0]  io_wgt_data_bits_30_2,
  input  [7:0]  io_wgt_data_bits_30_3,
  input  [7:0]  io_wgt_data_bits_30_4,
  input  [7:0]  io_wgt_data_bits_30_5,
  input  [7:0]  io_wgt_data_bits_30_6,
  input  [7:0]  io_wgt_data_bits_30_7,
  input  [7:0]  io_wgt_data_bits_30_8,
  input  [7:0]  io_wgt_data_bits_30_9,
  input  [7:0]  io_wgt_data_bits_30_10,
  input  [7:0]  io_wgt_data_bits_30_11,
  input  [7:0]  io_wgt_data_bits_30_12,
  input  [7:0]  io_wgt_data_bits_30_13,
  input  [7:0]  io_wgt_data_bits_30_14,
  input  [7:0]  io_wgt_data_bits_30_15,
  input  [7:0]  io_wgt_data_bits_31_0,
  input  [7:0]  io_wgt_data_bits_31_1,
  input  [7:0]  io_wgt_data_bits_31_2,
  input  [7:0]  io_wgt_data_bits_31_3,
  input  [7:0]  io_wgt_data_bits_31_4,
  input  [7:0]  io_wgt_data_bits_31_5,
  input  [7:0]  io_wgt_data_bits_31_6,
  input  [7:0]  io_wgt_data_bits_31_7,
  input  [7:0]  io_wgt_data_bits_31_8,
  input  [7:0]  io_wgt_data_bits_31_9,
  input  [7:0]  io_wgt_data_bits_31_10,
  input  [7:0]  io_wgt_data_bits_31_11,
  input  [7:0]  io_wgt_data_bits_31_12,
  input  [7:0]  io_wgt_data_bits_31_13,
  input  [7:0]  io_wgt_data_bits_31_14,
  input  [7:0]  io_wgt_data_bits_31_15,
  input         io_acc_i_data_valid,
  input  [31:0] io_acc_i_data_bits_0_0,
  input  [31:0] io_acc_i_data_bits_0_1,
  input  [31:0] io_acc_i_data_bits_0_2,
  input  [31:0] io_acc_i_data_bits_0_3,
  input  [31:0] io_acc_i_data_bits_0_4,
  input  [31:0] io_acc_i_data_bits_0_5,
  input  [31:0] io_acc_i_data_bits_0_6,
  input  [31:0] io_acc_i_data_bits_0_7,
  input  [31:0] io_acc_i_data_bits_0_8,
  input  [31:0] io_acc_i_data_bits_0_9,
  input  [31:0] io_acc_i_data_bits_0_10,
  input  [31:0] io_acc_i_data_bits_0_11,
  input  [31:0] io_acc_i_data_bits_0_12,
  input  [31:0] io_acc_i_data_bits_0_13,
  input  [31:0] io_acc_i_data_bits_0_14,
  input  [31:0] io_acc_i_data_bits_0_15,
  input  [31:0] io_acc_i_data_bits_0_16,
  input  [31:0] io_acc_i_data_bits_0_17,
  input  [31:0] io_acc_i_data_bits_0_18,
  input  [31:0] io_acc_i_data_bits_0_19,
  input  [31:0] io_acc_i_data_bits_0_20,
  input  [31:0] io_acc_i_data_bits_0_21,
  input  [31:0] io_acc_i_data_bits_0_22,
  input  [31:0] io_acc_i_data_bits_0_23,
  input  [31:0] io_acc_i_data_bits_0_24,
  input  [31:0] io_acc_i_data_bits_0_25,
  input  [31:0] io_acc_i_data_bits_0_26,
  input  [31:0] io_acc_i_data_bits_0_27,
  input  [31:0] io_acc_i_data_bits_0_28,
  input  [31:0] io_acc_i_data_bits_0_29,
  input  [31:0] io_acc_i_data_bits_0_30,
  input  [31:0] io_acc_i_data_bits_0_31,
  output        io_acc_o_data_valid,
  output [31:0] io_acc_o_data_bits_0_0,
  output [31:0] io_acc_o_data_bits_0_1,
  output [31:0] io_acc_o_data_bits_0_2,
  output [31:0] io_acc_o_data_bits_0_3,
  output [31:0] io_acc_o_data_bits_0_4,
  output [31:0] io_acc_o_data_bits_0_5,
  output [31:0] io_acc_o_data_bits_0_6,
  output [31:0] io_acc_o_data_bits_0_7,
  output [31:0] io_acc_o_data_bits_0_8,
  output [31:0] io_acc_o_data_bits_0_9,
  output [31:0] io_acc_o_data_bits_0_10,
  output [31:0] io_acc_o_data_bits_0_11,
  output [31:0] io_acc_o_data_bits_0_12,
  output [31:0] io_acc_o_data_bits_0_13,
  output [31:0] io_acc_o_data_bits_0_14,
  output [31:0] io_acc_o_data_bits_0_15,
  output [31:0] io_acc_o_data_bits_0_16,
  output [31:0] io_acc_o_data_bits_0_17,
  output [31:0] io_acc_o_data_bits_0_18,
  output [31:0] io_acc_o_data_bits_0_19,
  output [31:0] io_acc_o_data_bits_0_20,
  output [31:0] io_acc_o_data_bits_0_21,
  output [31:0] io_acc_o_data_bits_0_22,
  output [31:0] io_acc_o_data_bits_0_23,
  output [31:0] io_acc_o_data_bits_0_24,
  output [31:0] io_acc_o_data_bits_0_25,
  output [31:0] io_acc_o_data_bits_0_26,
  output [31:0] io_acc_o_data_bits_0_27,
  output [31:0] io_acc_o_data_bits_0_28,
  output [31:0] io_acc_o_data_bits_0_29,
  output [31:0] io_acc_o_data_bits_0_30,
  output [31:0] io_acc_o_data_bits_0_31,
  output        io_out_data_valid,
  output [7:0]  io_out_data_bits_0_0,
  output [7:0]  io_out_data_bits_0_1,
  output [7:0]  io_out_data_bits_0_2,
  output [7:0]  io_out_data_bits_0_3,
  output [7:0]  io_out_data_bits_0_4,
  output [7:0]  io_out_data_bits_0_5,
  output [7:0]  io_out_data_bits_0_6,
  output [7:0]  io_out_data_bits_0_7,
  output [7:0]  io_out_data_bits_0_8,
  output [7:0]  io_out_data_bits_0_9,
  output [7:0]  io_out_data_bits_0_10,
  output [7:0]  io_out_data_bits_0_11,
  output [7:0]  io_out_data_bits_0_12,
  output [7:0]  io_out_data_bits_0_13,
  output [7:0]  io_out_data_bits_0_14,
  output [7:0]  io_out_data_bits_0_15,
  output [7:0]  io_out_data_bits_0_16,
  output [7:0]  io_out_data_bits_0_17,
  output [7:0]  io_out_data_bits_0_18,
  output [7:0]  io_out_data_bits_0_19,
  output [7:0]  io_out_data_bits_0_20,
  output [7:0]  io_out_data_bits_0_21,
  output [7:0]  io_out_data_bits_0_22,
  output [7:0]  io_out_data_bits_0_23,
  output [7:0]  io_out_data_bits_0_24,
  output [7:0]  io_out_data_bits_0_25,
  output [7:0]  io_out_data_bits_0_26,
  output [7:0]  io_out_data_bits_0_27,
  output [7:0]  io_out_data_bits_0_28,
  output [7:0]  io_out_data_bits_0_29,
  output [7:0]  io_out_data_bits_0_30,
  output [7:0]  io_out_data_bits_0_31,
  input         io_bypass_cond
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  wire  dot_0_0_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_0_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_0_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_1_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_1_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_1_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_2_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_2_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_2_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_3_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_3_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_3_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_4_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_4_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_4_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_5_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_5_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_5_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_6_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_6_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_6_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_7_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_7_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_7_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_8_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_8_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_8_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_9_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_9_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_9_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_10_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_10_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_10_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_11_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_11_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_11_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_12_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_12_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_12_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_13_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_13_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_13_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_14_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_14_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_14_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_15_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_15_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_15_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_16_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_16_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_16_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_17_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_17_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_17_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_18_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_18_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_18_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_19_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_19_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_19_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_20_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_20_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_20_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_21_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_21_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_21_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_22_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_22_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_22_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_23_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_23_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_23_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_24_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_24_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_24_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_25_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_25_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_25_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_26_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_26_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_26_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_27_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_27_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_27_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_28_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_28_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_28_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_29_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_29_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_29_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_30_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_30_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_30_io_y; // @[TensorGemm.scala 198:11]
  wire  dot_0_31_clock; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_a_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_a_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_a_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_a_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_a_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_a_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_a_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_a_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_a_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_a_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_a_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_a_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_a_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_a_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_a_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_a_15; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_b_0; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_b_1; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_b_2; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_b_3; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_b_4; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_b_5; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_b_6; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_b_7; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_b_8; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_b_9; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_b_10; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_b_11; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_b_12; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_b_13; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_b_14; // @[TensorGemm.scala 198:11]
  wire [7:0] dot_0_31_io_b_15; // @[TensorGemm.scala 198:11]
  wire [20:0] dot_0_31_io_y; // @[TensorGemm.scala 198:11]
  reg [31:0] last_acc_write_0_0; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_1; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_2; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_3; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_4; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_5; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_6; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_7; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_8; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_9; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_10; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_11; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_12; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_13; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_14; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_15; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_16; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_17; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_18; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_19; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_20; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_21; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_22; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_23; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_24; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_25; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_26; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_27; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_28; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_29; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_30; // @[TensorGemm.scala 200:62]
  reg [31:0] last_acc_write_0_31; // @[TensorGemm.scala 200:62]
  wire [31:0] byp = io_bypass_cond ? $signed(last_acc_write_0_0) : $signed(io_acc_i_data_bits_0_0); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_0 = {{11{dot_0_0_io_y[20]}},dot_0_0_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_0 = $signed(byp) + $signed(_GEN_0); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_0_T = $signed(byp) + $signed(_GEN_0); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_1 = io_bypass_cond ? $signed(last_acc_write_0_1) : $signed(io_acc_i_data_bits_0_1); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_1 = {{11{dot_0_1_io_y[20]}},dot_0_1_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_1 = $signed(byp_1) + $signed(_GEN_1); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_1_T = $signed(byp_1) + $signed(_GEN_1); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_2 = io_bypass_cond ? $signed(last_acc_write_0_2) : $signed(io_acc_i_data_bits_0_2); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_2 = {{11{dot_0_2_io_y[20]}},dot_0_2_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_2 = $signed(byp_2) + $signed(_GEN_2); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_2_T = $signed(byp_2) + $signed(_GEN_2); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_3 = io_bypass_cond ? $signed(last_acc_write_0_3) : $signed(io_acc_i_data_bits_0_3); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_3 = {{11{dot_0_3_io_y[20]}},dot_0_3_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_3 = $signed(byp_3) + $signed(_GEN_3); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_3_T = $signed(byp_3) + $signed(_GEN_3); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_4 = io_bypass_cond ? $signed(last_acc_write_0_4) : $signed(io_acc_i_data_bits_0_4); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_4 = {{11{dot_0_4_io_y[20]}},dot_0_4_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_4 = $signed(byp_4) + $signed(_GEN_4); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_4_T = $signed(byp_4) + $signed(_GEN_4); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_5 = io_bypass_cond ? $signed(last_acc_write_0_5) : $signed(io_acc_i_data_bits_0_5); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_5 = {{11{dot_0_5_io_y[20]}},dot_0_5_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_5 = $signed(byp_5) + $signed(_GEN_5); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_5_T = $signed(byp_5) + $signed(_GEN_5); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_6 = io_bypass_cond ? $signed(last_acc_write_0_6) : $signed(io_acc_i_data_bits_0_6); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_6 = {{11{dot_0_6_io_y[20]}},dot_0_6_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_6 = $signed(byp_6) + $signed(_GEN_6); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_6_T = $signed(byp_6) + $signed(_GEN_6); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_7 = io_bypass_cond ? $signed(last_acc_write_0_7) : $signed(io_acc_i_data_bits_0_7); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_7 = {{11{dot_0_7_io_y[20]}},dot_0_7_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_7 = $signed(byp_7) + $signed(_GEN_7); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_7_T = $signed(byp_7) + $signed(_GEN_7); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_8 = io_bypass_cond ? $signed(last_acc_write_0_8) : $signed(io_acc_i_data_bits_0_8); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_8 = {{11{dot_0_8_io_y[20]}},dot_0_8_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_8 = $signed(byp_8) + $signed(_GEN_8); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_8_T = $signed(byp_8) + $signed(_GEN_8); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_9 = io_bypass_cond ? $signed(last_acc_write_0_9) : $signed(io_acc_i_data_bits_0_9); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_9 = {{11{dot_0_9_io_y[20]}},dot_0_9_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_9 = $signed(byp_9) + $signed(_GEN_9); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_9_T = $signed(byp_9) + $signed(_GEN_9); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_10 = io_bypass_cond ? $signed(last_acc_write_0_10) : $signed(io_acc_i_data_bits_0_10); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_10 = {{11{dot_0_10_io_y[20]}},dot_0_10_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_10 = $signed(byp_10) + $signed(_GEN_10); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_10_T = $signed(byp_10) + $signed(_GEN_10); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_11 = io_bypass_cond ? $signed(last_acc_write_0_11) : $signed(io_acc_i_data_bits_0_11); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_11 = {{11{dot_0_11_io_y[20]}},dot_0_11_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_11 = $signed(byp_11) + $signed(_GEN_11); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_11_T = $signed(byp_11) + $signed(_GEN_11); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_12 = io_bypass_cond ? $signed(last_acc_write_0_12) : $signed(io_acc_i_data_bits_0_12); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_12 = {{11{dot_0_12_io_y[20]}},dot_0_12_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_12 = $signed(byp_12) + $signed(_GEN_12); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_12_T = $signed(byp_12) + $signed(_GEN_12); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_13 = io_bypass_cond ? $signed(last_acc_write_0_13) : $signed(io_acc_i_data_bits_0_13); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_13 = {{11{dot_0_13_io_y[20]}},dot_0_13_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_13 = $signed(byp_13) + $signed(_GEN_13); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_13_T = $signed(byp_13) + $signed(_GEN_13); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_14 = io_bypass_cond ? $signed(last_acc_write_0_14) : $signed(io_acc_i_data_bits_0_14); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_14 = {{11{dot_0_14_io_y[20]}},dot_0_14_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_14 = $signed(byp_14) + $signed(_GEN_14); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_14_T = $signed(byp_14) + $signed(_GEN_14); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_15 = io_bypass_cond ? $signed(last_acc_write_0_15) : $signed(io_acc_i_data_bits_0_15); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_15 = {{11{dot_0_15_io_y[20]}},dot_0_15_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_15 = $signed(byp_15) + $signed(_GEN_15); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_15_T = $signed(byp_15) + $signed(_GEN_15); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_16 = io_bypass_cond ? $signed(last_acc_write_0_16) : $signed(io_acc_i_data_bits_0_16); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_16 = {{11{dot_0_16_io_y[20]}},dot_0_16_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_16 = $signed(byp_16) + $signed(_GEN_16); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_16_T = $signed(byp_16) + $signed(_GEN_16); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_17 = io_bypass_cond ? $signed(last_acc_write_0_17) : $signed(io_acc_i_data_bits_0_17); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_17 = {{11{dot_0_17_io_y[20]}},dot_0_17_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_17 = $signed(byp_17) + $signed(_GEN_17); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_17_T = $signed(byp_17) + $signed(_GEN_17); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_18 = io_bypass_cond ? $signed(last_acc_write_0_18) : $signed(io_acc_i_data_bits_0_18); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_18 = {{11{dot_0_18_io_y[20]}},dot_0_18_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_18 = $signed(byp_18) + $signed(_GEN_18); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_18_T = $signed(byp_18) + $signed(_GEN_18); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_19 = io_bypass_cond ? $signed(last_acc_write_0_19) : $signed(io_acc_i_data_bits_0_19); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_19 = {{11{dot_0_19_io_y[20]}},dot_0_19_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_19 = $signed(byp_19) + $signed(_GEN_19); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_19_T = $signed(byp_19) + $signed(_GEN_19); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_20 = io_bypass_cond ? $signed(last_acc_write_0_20) : $signed(io_acc_i_data_bits_0_20); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_20 = {{11{dot_0_20_io_y[20]}},dot_0_20_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_20 = $signed(byp_20) + $signed(_GEN_20); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_20_T = $signed(byp_20) + $signed(_GEN_20); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_21 = io_bypass_cond ? $signed(last_acc_write_0_21) : $signed(io_acc_i_data_bits_0_21); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_21 = {{11{dot_0_21_io_y[20]}},dot_0_21_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_21 = $signed(byp_21) + $signed(_GEN_21); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_21_T = $signed(byp_21) + $signed(_GEN_21); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_22 = io_bypass_cond ? $signed(last_acc_write_0_22) : $signed(io_acc_i_data_bits_0_22); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_22 = {{11{dot_0_22_io_y[20]}},dot_0_22_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_22 = $signed(byp_22) + $signed(_GEN_22); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_22_T = $signed(byp_22) + $signed(_GEN_22); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_23 = io_bypass_cond ? $signed(last_acc_write_0_23) : $signed(io_acc_i_data_bits_0_23); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_23 = {{11{dot_0_23_io_y[20]}},dot_0_23_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_23 = $signed(byp_23) + $signed(_GEN_23); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_23_T = $signed(byp_23) + $signed(_GEN_23); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_24 = io_bypass_cond ? $signed(last_acc_write_0_24) : $signed(io_acc_i_data_bits_0_24); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_24 = {{11{dot_0_24_io_y[20]}},dot_0_24_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_24 = $signed(byp_24) + $signed(_GEN_24); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_24_T = $signed(byp_24) + $signed(_GEN_24); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_25 = io_bypass_cond ? $signed(last_acc_write_0_25) : $signed(io_acc_i_data_bits_0_25); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_25 = {{11{dot_0_25_io_y[20]}},dot_0_25_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_25 = $signed(byp_25) + $signed(_GEN_25); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_25_T = $signed(byp_25) + $signed(_GEN_25); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_26 = io_bypass_cond ? $signed(last_acc_write_0_26) : $signed(io_acc_i_data_bits_0_26); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_26 = {{11{dot_0_26_io_y[20]}},dot_0_26_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_26 = $signed(byp_26) + $signed(_GEN_26); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_26_T = $signed(byp_26) + $signed(_GEN_26); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_27 = io_bypass_cond ? $signed(last_acc_write_0_27) : $signed(io_acc_i_data_bits_0_27); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_27 = {{11{dot_0_27_io_y[20]}},dot_0_27_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_27 = $signed(byp_27) + $signed(_GEN_27); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_27_T = $signed(byp_27) + $signed(_GEN_27); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_28 = io_bypass_cond ? $signed(last_acc_write_0_28) : $signed(io_acc_i_data_bits_0_28); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_28 = {{11{dot_0_28_io_y[20]}},dot_0_28_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_28 = $signed(byp_28) + $signed(_GEN_28); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_28_T = $signed(byp_28) + $signed(_GEN_28); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_29 = io_bypass_cond ? $signed(last_acc_write_0_29) : $signed(io_acc_i_data_bits_0_29); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_29 = {{11{dot_0_29_io_y[20]}},dot_0_29_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_29 = $signed(byp_29) + $signed(_GEN_29); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_29_T = $signed(byp_29) + $signed(_GEN_29); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_30 = io_bypass_cond ? $signed(last_acc_write_0_30) : $signed(io_acc_i_data_bits_0_30); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_30 = {{11{dot_0_30_io_y[20]}},dot_0_30_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_30 = $signed(byp_30) + $signed(_GEN_30); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_30_T = $signed(byp_30) + $signed(_GEN_30); // @[TensorGemm.scala 213:43]
  wire [31:0] byp_31 = io_bypass_cond ? $signed(last_acc_write_0_31) : $signed(io_acc_i_data_bits_0_31); // @[TensorGemm.scala 208:20]
  wire [31:0] _GEN_31 = {{11{dot_0_31_io_y[20]}},dot_0_31_io_y}; // @[TensorGemm.scala 209:24]
  wire [31:0] add_0_31 = $signed(byp_31) + $signed(_GEN_31); // @[TensorGemm.scala 209:24]
  wire [31:0] _io_out_data_bits_0_31_T = $signed(byp_31) + $signed(_GEN_31); // @[TensorGemm.scala 213:43]
  DotProduct dot_0_0 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_0_clock),
    .io_a_0(dot_0_0_io_a_0),
    .io_a_1(dot_0_0_io_a_1),
    .io_a_2(dot_0_0_io_a_2),
    .io_a_3(dot_0_0_io_a_3),
    .io_a_4(dot_0_0_io_a_4),
    .io_a_5(dot_0_0_io_a_5),
    .io_a_6(dot_0_0_io_a_6),
    .io_a_7(dot_0_0_io_a_7),
    .io_a_8(dot_0_0_io_a_8),
    .io_a_9(dot_0_0_io_a_9),
    .io_a_10(dot_0_0_io_a_10),
    .io_a_11(dot_0_0_io_a_11),
    .io_a_12(dot_0_0_io_a_12),
    .io_a_13(dot_0_0_io_a_13),
    .io_a_14(dot_0_0_io_a_14),
    .io_a_15(dot_0_0_io_a_15),
    .io_b_0(dot_0_0_io_b_0),
    .io_b_1(dot_0_0_io_b_1),
    .io_b_2(dot_0_0_io_b_2),
    .io_b_3(dot_0_0_io_b_3),
    .io_b_4(dot_0_0_io_b_4),
    .io_b_5(dot_0_0_io_b_5),
    .io_b_6(dot_0_0_io_b_6),
    .io_b_7(dot_0_0_io_b_7),
    .io_b_8(dot_0_0_io_b_8),
    .io_b_9(dot_0_0_io_b_9),
    .io_b_10(dot_0_0_io_b_10),
    .io_b_11(dot_0_0_io_b_11),
    .io_b_12(dot_0_0_io_b_12),
    .io_b_13(dot_0_0_io_b_13),
    .io_b_14(dot_0_0_io_b_14),
    .io_b_15(dot_0_0_io_b_15),
    .io_y(dot_0_0_io_y)
  );
  DotProduct dot_0_1 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_1_clock),
    .io_a_0(dot_0_1_io_a_0),
    .io_a_1(dot_0_1_io_a_1),
    .io_a_2(dot_0_1_io_a_2),
    .io_a_3(dot_0_1_io_a_3),
    .io_a_4(dot_0_1_io_a_4),
    .io_a_5(dot_0_1_io_a_5),
    .io_a_6(dot_0_1_io_a_6),
    .io_a_7(dot_0_1_io_a_7),
    .io_a_8(dot_0_1_io_a_8),
    .io_a_9(dot_0_1_io_a_9),
    .io_a_10(dot_0_1_io_a_10),
    .io_a_11(dot_0_1_io_a_11),
    .io_a_12(dot_0_1_io_a_12),
    .io_a_13(dot_0_1_io_a_13),
    .io_a_14(dot_0_1_io_a_14),
    .io_a_15(dot_0_1_io_a_15),
    .io_b_0(dot_0_1_io_b_0),
    .io_b_1(dot_0_1_io_b_1),
    .io_b_2(dot_0_1_io_b_2),
    .io_b_3(dot_0_1_io_b_3),
    .io_b_4(dot_0_1_io_b_4),
    .io_b_5(dot_0_1_io_b_5),
    .io_b_6(dot_0_1_io_b_6),
    .io_b_7(dot_0_1_io_b_7),
    .io_b_8(dot_0_1_io_b_8),
    .io_b_9(dot_0_1_io_b_9),
    .io_b_10(dot_0_1_io_b_10),
    .io_b_11(dot_0_1_io_b_11),
    .io_b_12(dot_0_1_io_b_12),
    .io_b_13(dot_0_1_io_b_13),
    .io_b_14(dot_0_1_io_b_14),
    .io_b_15(dot_0_1_io_b_15),
    .io_y(dot_0_1_io_y)
  );
  DotProduct dot_0_2 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_2_clock),
    .io_a_0(dot_0_2_io_a_0),
    .io_a_1(dot_0_2_io_a_1),
    .io_a_2(dot_0_2_io_a_2),
    .io_a_3(dot_0_2_io_a_3),
    .io_a_4(dot_0_2_io_a_4),
    .io_a_5(dot_0_2_io_a_5),
    .io_a_6(dot_0_2_io_a_6),
    .io_a_7(dot_0_2_io_a_7),
    .io_a_8(dot_0_2_io_a_8),
    .io_a_9(dot_0_2_io_a_9),
    .io_a_10(dot_0_2_io_a_10),
    .io_a_11(dot_0_2_io_a_11),
    .io_a_12(dot_0_2_io_a_12),
    .io_a_13(dot_0_2_io_a_13),
    .io_a_14(dot_0_2_io_a_14),
    .io_a_15(dot_0_2_io_a_15),
    .io_b_0(dot_0_2_io_b_0),
    .io_b_1(dot_0_2_io_b_1),
    .io_b_2(dot_0_2_io_b_2),
    .io_b_3(dot_0_2_io_b_3),
    .io_b_4(dot_0_2_io_b_4),
    .io_b_5(dot_0_2_io_b_5),
    .io_b_6(dot_0_2_io_b_6),
    .io_b_7(dot_0_2_io_b_7),
    .io_b_8(dot_0_2_io_b_8),
    .io_b_9(dot_0_2_io_b_9),
    .io_b_10(dot_0_2_io_b_10),
    .io_b_11(dot_0_2_io_b_11),
    .io_b_12(dot_0_2_io_b_12),
    .io_b_13(dot_0_2_io_b_13),
    .io_b_14(dot_0_2_io_b_14),
    .io_b_15(dot_0_2_io_b_15),
    .io_y(dot_0_2_io_y)
  );
  DotProduct dot_0_3 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_3_clock),
    .io_a_0(dot_0_3_io_a_0),
    .io_a_1(dot_0_3_io_a_1),
    .io_a_2(dot_0_3_io_a_2),
    .io_a_3(dot_0_3_io_a_3),
    .io_a_4(dot_0_3_io_a_4),
    .io_a_5(dot_0_3_io_a_5),
    .io_a_6(dot_0_3_io_a_6),
    .io_a_7(dot_0_3_io_a_7),
    .io_a_8(dot_0_3_io_a_8),
    .io_a_9(dot_0_3_io_a_9),
    .io_a_10(dot_0_3_io_a_10),
    .io_a_11(dot_0_3_io_a_11),
    .io_a_12(dot_0_3_io_a_12),
    .io_a_13(dot_0_3_io_a_13),
    .io_a_14(dot_0_3_io_a_14),
    .io_a_15(dot_0_3_io_a_15),
    .io_b_0(dot_0_3_io_b_0),
    .io_b_1(dot_0_3_io_b_1),
    .io_b_2(dot_0_3_io_b_2),
    .io_b_3(dot_0_3_io_b_3),
    .io_b_4(dot_0_3_io_b_4),
    .io_b_5(dot_0_3_io_b_5),
    .io_b_6(dot_0_3_io_b_6),
    .io_b_7(dot_0_3_io_b_7),
    .io_b_8(dot_0_3_io_b_8),
    .io_b_9(dot_0_3_io_b_9),
    .io_b_10(dot_0_3_io_b_10),
    .io_b_11(dot_0_3_io_b_11),
    .io_b_12(dot_0_3_io_b_12),
    .io_b_13(dot_0_3_io_b_13),
    .io_b_14(dot_0_3_io_b_14),
    .io_b_15(dot_0_3_io_b_15),
    .io_y(dot_0_3_io_y)
  );
  DotProduct dot_0_4 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_4_clock),
    .io_a_0(dot_0_4_io_a_0),
    .io_a_1(dot_0_4_io_a_1),
    .io_a_2(dot_0_4_io_a_2),
    .io_a_3(dot_0_4_io_a_3),
    .io_a_4(dot_0_4_io_a_4),
    .io_a_5(dot_0_4_io_a_5),
    .io_a_6(dot_0_4_io_a_6),
    .io_a_7(dot_0_4_io_a_7),
    .io_a_8(dot_0_4_io_a_8),
    .io_a_9(dot_0_4_io_a_9),
    .io_a_10(dot_0_4_io_a_10),
    .io_a_11(dot_0_4_io_a_11),
    .io_a_12(dot_0_4_io_a_12),
    .io_a_13(dot_0_4_io_a_13),
    .io_a_14(dot_0_4_io_a_14),
    .io_a_15(dot_0_4_io_a_15),
    .io_b_0(dot_0_4_io_b_0),
    .io_b_1(dot_0_4_io_b_1),
    .io_b_2(dot_0_4_io_b_2),
    .io_b_3(dot_0_4_io_b_3),
    .io_b_4(dot_0_4_io_b_4),
    .io_b_5(dot_0_4_io_b_5),
    .io_b_6(dot_0_4_io_b_6),
    .io_b_7(dot_0_4_io_b_7),
    .io_b_8(dot_0_4_io_b_8),
    .io_b_9(dot_0_4_io_b_9),
    .io_b_10(dot_0_4_io_b_10),
    .io_b_11(dot_0_4_io_b_11),
    .io_b_12(dot_0_4_io_b_12),
    .io_b_13(dot_0_4_io_b_13),
    .io_b_14(dot_0_4_io_b_14),
    .io_b_15(dot_0_4_io_b_15),
    .io_y(dot_0_4_io_y)
  );
  DotProduct dot_0_5 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_5_clock),
    .io_a_0(dot_0_5_io_a_0),
    .io_a_1(dot_0_5_io_a_1),
    .io_a_2(dot_0_5_io_a_2),
    .io_a_3(dot_0_5_io_a_3),
    .io_a_4(dot_0_5_io_a_4),
    .io_a_5(dot_0_5_io_a_5),
    .io_a_6(dot_0_5_io_a_6),
    .io_a_7(dot_0_5_io_a_7),
    .io_a_8(dot_0_5_io_a_8),
    .io_a_9(dot_0_5_io_a_9),
    .io_a_10(dot_0_5_io_a_10),
    .io_a_11(dot_0_5_io_a_11),
    .io_a_12(dot_0_5_io_a_12),
    .io_a_13(dot_0_5_io_a_13),
    .io_a_14(dot_0_5_io_a_14),
    .io_a_15(dot_0_5_io_a_15),
    .io_b_0(dot_0_5_io_b_0),
    .io_b_1(dot_0_5_io_b_1),
    .io_b_2(dot_0_5_io_b_2),
    .io_b_3(dot_0_5_io_b_3),
    .io_b_4(dot_0_5_io_b_4),
    .io_b_5(dot_0_5_io_b_5),
    .io_b_6(dot_0_5_io_b_6),
    .io_b_7(dot_0_5_io_b_7),
    .io_b_8(dot_0_5_io_b_8),
    .io_b_9(dot_0_5_io_b_9),
    .io_b_10(dot_0_5_io_b_10),
    .io_b_11(dot_0_5_io_b_11),
    .io_b_12(dot_0_5_io_b_12),
    .io_b_13(dot_0_5_io_b_13),
    .io_b_14(dot_0_5_io_b_14),
    .io_b_15(dot_0_5_io_b_15),
    .io_y(dot_0_5_io_y)
  );
  DotProduct dot_0_6 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_6_clock),
    .io_a_0(dot_0_6_io_a_0),
    .io_a_1(dot_0_6_io_a_1),
    .io_a_2(dot_0_6_io_a_2),
    .io_a_3(dot_0_6_io_a_3),
    .io_a_4(dot_0_6_io_a_4),
    .io_a_5(dot_0_6_io_a_5),
    .io_a_6(dot_0_6_io_a_6),
    .io_a_7(dot_0_6_io_a_7),
    .io_a_8(dot_0_6_io_a_8),
    .io_a_9(dot_0_6_io_a_9),
    .io_a_10(dot_0_6_io_a_10),
    .io_a_11(dot_0_6_io_a_11),
    .io_a_12(dot_0_6_io_a_12),
    .io_a_13(dot_0_6_io_a_13),
    .io_a_14(dot_0_6_io_a_14),
    .io_a_15(dot_0_6_io_a_15),
    .io_b_0(dot_0_6_io_b_0),
    .io_b_1(dot_0_6_io_b_1),
    .io_b_2(dot_0_6_io_b_2),
    .io_b_3(dot_0_6_io_b_3),
    .io_b_4(dot_0_6_io_b_4),
    .io_b_5(dot_0_6_io_b_5),
    .io_b_6(dot_0_6_io_b_6),
    .io_b_7(dot_0_6_io_b_7),
    .io_b_8(dot_0_6_io_b_8),
    .io_b_9(dot_0_6_io_b_9),
    .io_b_10(dot_0_6_io_b_10),
    .io_b_11(dot_0_6_io_b_11),
    .io_b_12(dot_0_6_io_b_12),
    .io_b_13(dot_0_6_io_b_13),
    .io_b_14(dot_0_6_io_b_14),
    .io_b_15(dot_0_6_io_b_15),
    .io_y(dot_0_6_io_y)
  );
  DotProduct dot_0_7 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_7_clock),
    .io_a_0(dot_0_7_io_a_0),
    .io_a_1(dot_0_7_io_a_1),
    .io_a_2(dot_0_7_io_a_2),
    .io_a_3(dot_0_7_io_a_3),
    .io_a_4(dot_0_7_io_a_4),
    .io_a_5(dot_0_7_io_a_5),
    .io_a_6(dot_0_7_io_a_6),
    .io_a_7(dot_0_7_io_a_7),
    .io_a_8(dot_0_7_io_a_8),
    .io_a_9(dot_0_7_io_a_9),
    .io_a_10(dot_0_7_io_a_10),
    .io_a_11(dot_0_7_io_a_11),
    .io_a_12(dot_0_7_io_a_12),
    .io_a_13(dot_0_7_io_a_13),
    .io_a_14(dot_0_7_io_a_14),
    .io_a_15(dot_0_7_io_a_15),
    .io_b_0(dot_0_7_io_b_0),
    .io_b_1(dot_0_7_io_b_1),
    .io_b_2(dot_0_7_io_b_2),
    .io_b_3(dot_0_7_io_b_3),
    .io_b_4(dot_0_7_io_b_4),
    .io_b_5(dot_0_7_io_b_5),
    .io_b_6(dot_0_7_io_b_6),
    .io_b_7(dot_0_7_io_b_7),
    .io_b_8(dot_0_7_io_b_8),
    .io_b_9(dot_0_7_io_b_9),
    .io_b_10(dot_0_7_io_b_10),
    .io_b_11(dot_0_7_io_b_11),
    .io_b_12(dot_0_7_io_b_12),
    .io_b_13(dot_0_7_io_b_13),
    .io_b_14(dot_0_7_io_b_14),
    .io_b_15(dot_0_7_io_b_15),
    .io_y(dot_0_7_io_y)
  );
  DotProduct dot_0_8 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_8_clock),
    .io_a_0(dot_0_8_io_a_0),
    .io_a_1(dot_0_8_io_a_1),
    .io_a_2(dot_0_8_io_a_2),
    .io_a_3(dot_0_8_io_a_3),
    .io_a_4(dot_0_8_io_a_4),
    .io_a_5(dot_0_8_io_a_5),
    .io_a_6(dot_0_8_io_a_6),
    .io_a_7(dot_0_8_io_a_7),
    .io_a_8(dot_0_8_io_a_8),
    .io_a_9(dot_0_8_io_a_9),
    .io_a_10(dot_0_8_io_a_10),
    .io_a_11(dot_0_8_io_a_11),
    .io_a_12(dot_0_8_io_a_12),
    .io_a_13(dot_0_8_io_a_13),
    .io_a_14(dot_0_8_io_a_14),
    .io_a_15(dot_0_8_io_a_15),
    .io_b_0(dot_0_8_io_b_0),
    .io_b_1(dot_0_8_io_b_1),
    .io_b_2(dot_0_8_io_b_2),
    .io_b_3(dot_0_8_io_b_3),
    .io_b_4(dot_0_8_io_b_4),
    .io_b_5(dot_0_8_io_b_5),
    .io_b_6(dot_0_8_io_b_6),
    .io_b_7(dot_0_8_io_b_7),
    .io_b_8(dot_0_8_io_b_8),
    .io_b_9(dot_0_8_io_b_9),
    .io_b_10(dot_0_8_io_b_10),
    .io_b_11(dot_0_8_io_b_11),
    .io_b_12(dot_0_8_io_b_12),
    .io_b_13(dot_0_8_io_b_13),
    .io_b_14(dot_0_8_io_b_14),
    .io_b_15(dot_0_8_io_b_15),
    .io_y(dot_0_8_io_y)
  );
  DotProduct dot_0_9 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_9_clock),
    .io_a_0(dot_0_9_io_a_0),
    .io_a_1(dot_0_9_io_a_1),
    .io_a_2(dot_0_9_io_a_2),
    .io_a_3(dot_0_9_io_a_3),
    .io_a_4(dot_0_9_io_a_4),
    .io_a_5(dot_0_9_io_a_5),
    .io_a_6(dot_0_9_io_a_6),
    .io_a_7(dot_0_9_io_a_7),
    .io_a_8(dot_0_9_io_a_8),
    .io_a_9(dot_0_9_io_a_9),
    .io_a_10(dot_0_9_io_a_10),
    .io_a_11(dot_0_9_io_a_11),
    .io_a_12(dot_0_9_io_a_12),
    .io_a_13(dot_0_9_io_a_13),
    .io_a_14(dot_0_9_io_a_14),
    .io_a_15(dot_0_9_io_a_15),
    .io_b_0(dot_0_9_io_b_0),
    .io_b_1(dot_0_9_io_b_1),
    .io_b_2(dot_0_9_io_b_2),
    .io_b_3(dot_0_9_io_b_3),
    .io_b_4(dot_0_9_io_b_4),
    .io_b_5(dot_0_9_io_b_5),
    .io_b_6(dot_0_9_io_b_6),
    .io_b_7(dot_0_9_io_b_7),
    .io_b_8(dot_0_9_io_b_8),
    .io_b_9(dot_0_9_io_b_9),
    .io_b_10(dot_0_9_io_b_10),
    .io_b_11(dot_0_9_io_b_11),
    .io_b_12(dot_0_9_io_b_12),
    .io_b_13(dot_0_9_io_b_13),
    .io_b_14(dot_0_9_io_b_14),
    .io_b_15(dot_0_9_io_b_15),
    .io_y(dot_0_9_io_y)
  );
  DotProduct dot_0_10 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_10_clock),
    .io_a_0(dot_0_10_io_a_0),
    .io_a_1(dot_0_10_io_a_1),
    .io_a_2(dot_0_10_io_a_2),
    .io_a_3(dot_0_10_io_a_3),
    .io_a_4(dot_0_10_io_a_4),
    .io_a_5(dot_0_10_io_a_5),
    .io_a_6(dot_0_10_io_a_6),
    .io_a_7(dot_0_10_io_a_7),
    .io_a_8(dot_0_10_io_a_8),
    .io_a_9(dot_0_10_io_a_9),
    .io_a_10(dot_0_10_io_a_10),
    .io_a_11(dot_0_10_io_a_11),
    .io_a_12(dot_0_10_io_a_12),
    .io_a_13(dot_0_10_io_a_13),
    .io_a_14(dot_0_10_io_a_14),
    .io_a_15(dot_0_10_io_a_15),
    .io_b_0(dot_0_10_io_b_0),
    .io_b_1(dot_0_10_io_b_1),
    .io_b_2(dot_0_10_io_b_2),
    .io_b_3(dot_0_10_io_b_3),
    .io_b_4(dot_0_10_io_b_4),
    .io_b_5(dot_0_10_io_b_5),
    .io_b_6(dot_0_10_io_b_6),
    .io_b_7(dot_0_10_io_b_7),
    .io_b_8(dot_0_10_io_b_8),
    .io_b_9(dot_0_10_io_b_9),
    .io_b_10(dot_0_10_io_b_10),
    .io_b_11(dot_0_10_io_b_11),
    .io_b_12(dot_0_10_io_b_12),
    .io_b_13(dot_0_10_io_b_13),
    .io_b_14(dot_0_10_io_b_14),
    .io_b_15(dot_0_10_io_b_15),
    .io_y(dot_0_10_io_y)
  );
  DotProduct dot_0_11 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_11_clock),
    .io_a_0(dot_0_11_io_a_0),
    .io_a_1(dot_0_11_io_a_1),
    .io_a_2(dot_0_11_io_a_2),
    .io_a_3(dot_0_11_io_a_3),
    .io_a_4(dot_0_11_io_a_4),
    .io_a_5(dot_0_11_io_a_5),
    .io_a_6(dot_0_11_io_a_6),
    .io_a_7(dot_0_11_io_a_7),
    .io_a_8(dot_0_11_io_a_8),
    .io_a_9(dot_0_11_io_a_9),
    .io_a_10(dot_0_11_io_a_10),
    .io_a_11(dot_0_11_io_a_11),
    .io_a_12(dot_0_11_io_a_12),
    .io_a_13(dot_0_11_io_a_13),
    .io_a_14(dot_0_11_io_a_14),
    .io_a_15(dot_0_11_io_a_15),
    .io_b_0(dot_0_11_io_b_0),
    .io_b_1(dot_0_11_io_b_1),
    .io_b_2(dot_0_11_io_b_2),
    .io_b_3(dot_0_11_io_b_3),
    .io_b_4(dot_0_11_io_b_4),
    .io_b_5(dot_0_11_io_b_5),
    .io_b_6(dot_0_11_io_b_6),
    .io_b_7(dot_0_11_io_b_7),
    .io_b_8(dot_0_11_io_b_8),
    .io_b_9(dot_0_11_io_b_9),
    .io_b_10(dot_0_11_io_b_10),
    .io_b_11(dot_0_11_io_b_11),
    .io_b_12(dot_0_11_io_b_12),
    .io_b_13(dot_0_11_io_b_13),
    .io_b_14(dot_0_11_io_b_14),
    .io_b_15(dot_0_11_io_b_15),
    .io_y(dot_0_11_io_y)
  );
  DotProduct dot_0_12 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_12_clock),
    .io_a_0(dot_0_12_io_a_0),
    .io_a_1(dot_0_12_io_a_1),
    .io_a_2(dot_0_12_io_a_2),
    .io_a_3(dot_0_12_io_a_3),
    .io_a_4(dot_0_12_io_a_4),
    .io_a_5(dot_0_12_io_a_5),
    .io_a_6(dot_0_12_io_a_6),
    .io_a_7(dot_0_12_io_a_7),
    .io_a_8(dot_0_12_io_a_8),
    .io_a_9(dot_0_12_io_a_9),
    .io_a_10(dot_0_12_io_a_10),
    .io_a_11(dot_0_12_io_a_11),
    .io_a_12(dot_0_12_io_a_12),
    .io_a_13(dot_0_12_io_a_13),
    .io_a_14(dot_0_12_io_a_14),
    .io_a_15(dot_0_12_io_a_15),
    .io_b_0(dot_0_12_io_b_0),
    .io_b_1(dot_0_12_io_b_1),
    .io_b_2(dot_0_12_io_b_2),
    .io_b_3(dot_0_12_io_b_3),
    .io_b_4(dot_0_12_io_b_4),
    .io_b_5(dot_0_12_io_b_5),
    .io_b_6(dot_0_12_io_b_6),
    .io_b_7(dot_0_12_io_b_7),
    .io_b_8(dot_0_12_io_b_8),
    .io_b_9(dot_0_12_io_b_9),
    .io_b_10(dot_0_12_io_b_10),
    .io_b_11(dot_0_12_io_b_11),
    .io_b_12(dot_0_12_io_b_12),
    .io_b_13(dot_0_12_io_b_13),
    .io_b_14(dot_0_12_io_b_14),
    .io_b_15(dot_0_12_io_b_15),
    .io_y(dot_0_12_io_y)
  );
  DotProduct dot_0_13 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_13_clock),
    .io_a_0(dot_0_13_io_a_0),
    .io_a_1(dot_0_13_io_a_1),
    .io_a_2(dot_0_13_io_a_2),
    .io_a_3(dot_0_13_io_a_3),
    .io_a_4(dot_0_13_io_a_4),
    .io_a_5(dot_0_13_io_a_5),
    .io_a_6(dot_0_13_io_a_6),
    .io_a_7(dot_0_13_io_a_7),
    .io_a_8(dot_0_13_io_a_8),
    .io_a_9(dot_0_13_io_a_9),
    .io_a_10(dot_0_13_io_a_10),
    .io_a_11(dot_0_13_io_a_11),
    .io_a_12(dot_0_13_io_a_12),
    .io_a_13(dot_0_13_io_a_13),
    .io_a_14(dot_0_13_io_a_14),
    .io_a_15(dot_0_13_io_a_15),
    .io_b_0(dot_0_13_io_b_0),
    .io_b_1(dot_0_13_io_b_1),
    .io_b_2(dot_0_13_io_b_2),
    .io_b_3(dot_0_13_io_b_3),
    .io_b_4(dot_0_13_io_b_4),
    .io_b_5(dot_0_13_io_b_5),
    .io_b_6(dot_0_13_io_b_6),
    .io_b_7(dot_0_13_io_b_7),
    .io_b_8(dot_0_13_io_b_8),
    .io_b_9(dot_0_13_io_b_9),
    .io_b_10(dot_0_13_io_b_10),
    .io_b_11(dot_0_13_io_b_11),
    .io_b_12(dot_0_13_io_b_12),
    .io_b_13(dot_0_13_io_b_13),
    .io_b_14(dot_0_13_io_b_14),
    .io_b_15(dot_0_13_io_b_15),
    .io_y(dot_0_13_io_y)
  );
  DotProduct dot_0_14 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_14_clock),
    .io_a_0(dot_0_14_io_a_0),
    .io_a_1(dot_0_14_io_a_1),
    .io_a_2(dot_0_14_io_a_2),
    .io_a_3(dot_0_14_io_a_3),
    .io_a_4(dot_0_14_io_a_4),
    .io_a_5(dot_0_14_io_a_5),
    .io_a_6(dot_0_14_io_a_6),
    .io_a_7(dot_0_14_io_a_7),
    .io_a_8(dot_0_14_io_a_8),
    .io_a_9(dot_0_14_io_a_9),
    .io_a_10(dot_0_14_io_a_10),
    .io_a_11(dot_0_14_io_a_11),
    .io_a_12(dot_0_14_io_a_12),
    .io_a_13(dot_0_14_io_a_13),
    .io_a_14(dot_0_14_io_a_14),
    .io_a_15(dot_0_14_io_a_15),
    .io_b_0(dot_0_14_io_b_0),
    .io_b_1(dot_0_14_io_b_1),
    .io_b_2(dot_0_14_io_b_2),
    .io_b_3(dot_0_14_io_b_3),
    .io_b_4(dot_0_14_io_b_4),
    .io_b_5(dot_0_14_io_b_5),
    .io_b_6(dot_0_14_io_b_6),
    .io_b_7(dot_0_14_io_b_7),
    .io_b_8(dot_0_14_io_b_8),
    .io_b_9(dot_0_14_io_b_9),
    .io_b_10(dot_0_14_io_b_10),
    .io_b_11(dot_0_14_io_b_11),
    .io_b_12(dot_0_14_io_b_12),
    .io_b_13(dot_0_14_io_b_13),
    .io_b_14(dot_0_14_io_b_14),
    .io_b_15(dot_0_14_io_b_15),
    .io_y(dot_0_14_io_y)
  );
  DotProduct dot_0_15 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_15_clock),
    .io_a_0(dot_0_15_io_a_0),
    .io_a_1(dot_0_15_io_a_1),
    .io_a_2(dot_0_15_io_a_2),
    .io_a_3(dot_0_15_io_a_3),
    .io_a_4(dot_0_15_io_a_4),
    .io_a_5(dot_0_15_io_a_5),
    .io_a_6(dot_0_15_io_a_6),
    .io_a_7(dot_0_15_io_a_7),
    .io_a_8(dot_0_15_io_a_8),
    .io_a_9(dot_0_15_io_a_9),
    .io_a_10(dot_0_15_io_a_10),
    .io_a_11(dot_0_15_io_a_11),
    .io_a_12(dot_0_15_io_a_12),
    .io_a_13(dot_0_15_io_a_13),
    .io_a_14(dot_0_15_io_a_14),
    .io_a_15(dot_0_15_io_a_15),
    .io_b_0(dot_0_15_io_b_0),
    .io_b_1(dot_0_15_io_b_1),
    .io_b_2(dot_0_15_io_b_2),
    .io_b_3(dot_0_15_io_b_3),
    .io_b_4(dot_0_15_io_b_4),
    .io_b_5(dot_0_15_io_b_5),
    .io_b_6(dot_0_15_io_b_6),
    .io_b_7(dot_0_15_io_b_7),
    .io_b_8(dot_0_15_io_b_8),
    .io_b_9(dot_0_15_io_b_9),
    .io_b_10(dot_0_15_io_b_10),
    .io_b_11(dot_0_15_io_b_11),
    .io_b_12(dot_0_15_io_b_12),
    .io_b_13(dot_0_15_io_b_13),
    .io_b_14(dot_0_15_io_b_14),
    .io_b_15(dot_0_15_io_b_15),
    .io_y(dot_0_15_io_y)
  );
  DotProduct dot_0_16 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_16_clock),
    .io_a_0(dot_0_16_io_a_0),
    .io_a_1(dot_0_16_io_a_1),
    .io_a_2(dot_0_16_io_a_2),
    .io_a_3(dot_0_16_io_a_3),
    .io_a_4(dot_0_16_io_a_4),
    .io_a_5(dot_0_16_io_a_5),
    .io_a_6(dot_0_16_io_a_6),
    .io_a_7(dot_0_16_io_a_7),
    .io_a_8(dot_0_16_io_a_8),
    .io_a_9(dot_0_16_io_a_9),
    .io_a_10(dot_0_16_io_a_10),
    .io_a_11(dot_0_16_io_a_11),
    .io_a_12(dot_0_16_io_a_12),
    .io_a_13(dot_0_16_io_a_13),
    .io_a_14(dot_0_16_io_a_14),
    .io_a_15(dot_0_16_io_a_15),
    .io_b_0(dot_0_16_io_b_0),
    .io_b_1(dot_0_16_io_b_1),
    .io_b_2(dot_0_16_io_b_2),
    .io_b_3(dot_0_16_io_b_3),
    .io_b_4(dot_0_16_io_b_4),
    .io_b_5(dot_0_16_io_b_5),
    .io_b_6(dot_0_16_io_b_6),
    .io_b_7(dot_0_16_io_b_7),
    .io_b_8(dot_0_16_io_b_8),
    .io_b_9(dot_0_16_io_b_9),
    .io_b_10(dot_0_16_io_b_10),
    .io_b_11(dot_0_16_io_b_11),
    .io_b_12(dot_0_16_io_b_12),
    .io_b_13(dot_0_16_io_b_13),
    .io_b_14(dot_0_16_io_b_14),
    .io_b_15(dot_0_16_io_b_15),
    .io_y(dot_0_16_io_y)
  );
  DotProduct dot_0_17 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_17_clock),
    .io_a_0(dot_0_17_io_a_0),
    .io_a_1(dot_0_17_io_a_1),
    .io_a_2(dot_0_17_io_a_2),
    .io_a_3(dot_0_17_io_a_3),
    .io_a_4(dot_0_17_io_a_4),
    .io_a_5(dot_0_17_io_a_5),
    .io_a_6(dot_0_17_io_a_6),
    .io_a_7(dot_0_17_io_a_7),
    .io_a_8(dot_0_17_io_a_8),
    .io_a_9(dot_0_17_io_a_9),
    .io_a_10(dot_0_17_io_a_10),
    .io_a_11(dot_0_17_io_a_11),
    .io_a_12(dot_0_17_io_a_12),
    .io_a_13(dot_0_17_io_a_13),
    .io_a_14(dot_0_17_io_a_14),
    .io_a_15(dot_0_17_io_a_15),
    .io_b_0(dot_0_17_io_b_0),
    .io_b_1(dot_0_17_io_b_1),
    .io_b_2(dot_0_17_io_b_2),
    .io_b_3(dot_0_17_io_b_3),
    .io_b_4(dot_0_17_io_b_4),
    .io_b_5(dot_0_17_io_b_5),
    .io_b_6(dot_0_17_io_b_6),
    .io_b_7(dot_0_17_io_b_7),
    .io_b_8(dot_0_17_io_b_8),
    .io_b_9(dot_0_17_io_b_9),
    .io_b_10(dot_0_17_io_b_10),
    .io_b_11(dot_0_17_io_b_11),
    .io_b_12(dot_0_17_io_b_12),
    .io_b_13(dot_0_17_io_b_13),
    .io_b_14(dot_0_17_io_b_14),
    .io_b_15(dot_0_17_io_b_15),
    .io_y(dot_0_17_io_y)
  );
  DotProduct dot_0_18 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_18_clock),
    .io_a_0(dot_0_18_io_a_0),
    .io_a_1(dot_0_18_io_a_1),
    .io_a_2(dot_0_18_io_a_2),
    .io_a_3(dot_0_18_io_a_3),
    .io_a_4(dot_0_18_io_a_4),
    .io_a_5(dot_0_18_io_a_5),
    .io_a_6(dot_0_18_io_a_6),
    .io_a_7(dot_0_18_io_a_7),
    .io_a_8(dot_0_18_io_a_8),
    .io_a_9(dot_0_18_io_a_9),
    .io_a_10(dot_0_18_io_a_10),
    .io_a_11(dot_0_18_io_a_11),
    .io_a_12(dot_0_18_io_a_12),
    .io_a_13(dot_0_18_io_a_13),
    .io_a_14(dot_0_18_io_a_14),
    .io_a_15(dot_0_18_io_a_15),
    .io_b_0(dot_0_18_io_b_0),
    .io_b_1(dot_0_18_io_b_1),
    .io_b_2(dot_0_18_io_b_2),
    .io_b_3(dot_0_18_io_b_3),
    .io_b_4(dot_0_18_io_b_4),
    .io_b_5(dot_0_18_io_b_5),
    .io_b_6(dot_0_18_io_b_6),
    .io_b_7(dot_0_18_io_b_7),
    .io_b_8(dot_0_18_io_b_8),
    .io_b_9(dot_0_18_io_b_9),
    .io_b_10(dot_0_18_io_b_10),
    .io_b_11(dot_0_18_io_b_11),
    .io_b_12(dot_0_18_io_b_12),
    .io_b_13(dot_0_18_io_b_13),
    .io_b_14(dot_0_18_io_b_14),
    .io_b_15(dot_0_18_io_b_15),
    .io_y(dot_0_18_io_y)
  );
  DotProduct dot_0_19 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_19_clock),
    .io_a_0(dot_0_19_io_a_0),
    .io_a_1(dot_0_19_io_a_1),
    .io_a_2(dot_0_19_io_a_2),
    .io_a_3(dot_0_19_io_a_3),
    .io_a_4(dot_0_19_io_a_4),
    .io_a_5(dot_0_19_io_a_5),
    .io_a_6(dot_0_19_io_a_6),
    .io_a_7(dot_0_19_io_a_7),
    .io_a_8(dot_0_19_io_a_8),
    .io_a_9(dot_0_19_io_a_9),
    .io_a_10(dot_0_19_io_a_10),
    .io_a_11(dot_0_19_io_a_11),
    .io_a_12(dot_0_19_io_a_12),
    .io_a_13(dot_0_19_io_a_13),
    .io_a_14(dot_0_19_io_a_14),
    .io_a_15(dot_0_19_io_a_15),
    .io_b_0(dot_0_19_io_b_0),
    .io_b_1(dot_0_19_io_b_1),
    .io_b_2(dot_0_19_io_b_2),
    .io_b_3(dot_0_19_io_b_3),
    .io_b_4(dot_0_19_io_b_4),
    .io_b_5(dot_0_19_io_b_5),
    .io_b_6(dot_0_19_io_b_6),
    .io_b_7(dot_0_19_io_b_7),
    .io_b_8(dot_0_19_io_b_8),
    .io_b_9(dot_0_19_io_b_9),
    .io_b_10(dot_0_19_io_b_10),
    .io_b_11(dot_0_19_io_b_11),
    .io_b_12(dot_0_19_io_b_12),
    .io_b_13(dot_0_19_io_b_13),
    .io_b_14(dot_0_19_io_b_14),
    .io_b_15(dot_0_19_io_b_15),
    .io_y(dot_0_19_io_y)
  );
  DotProduct dot_0_20 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_20_clock),
    .io_a_0(dot_0_20_io_a_0),
    .io_a_1(dot_0_20_io_a_1),
    .io_a_2(dot_0_20_io_a_2),
    .io_a_3(dot_0_20_io_a_3),
    .io_a_4(dot_0_20_io_a_4),
    .io_a_5(dot_0_20_io_a_5),
    .io_a_6(dot_0_20_io_a_6),
    .io_a_7(dot_0_20_io_a_7),
    .io_a_8(dot_0_20_io_a_8),
    .io_a_9(dot_0_20_io_a_9),
    .io_a_10(dot_0_20_io_a_10),
    .io_a_11(dot_0_20_io_a_11),
    .io_a_12(dot_0_20_io_a_12),
    .io_a_13(dot_0_20_io_a_13),
    .io_a_14(dot_0_20_io_a_14),
    .io_a_15(dot_0_20_io_a_15),
    .io_b_0(dot_0_20_io_b_0),
    .io_b_1(dot_0_20_io_b_1),
    .io_b_2(dot_0_20_io_b_2),
    .io_b_3(dot_0_20_io_b_3),
    .io_b_4(dot_0_20_io_b_4),
    .io_b_5(dot_0_20_io_b_5),
    .io_b_6(dot_0_20_io_b_6),
    .io_b_7(dot_0_20_io_b_7),
    .io_b_8(dot_0_20_io_b_8),
    .io_b_9(dot_0_20_io_b_9),
    .io_b_10(dot_0_20_io_b_10),
    .io_b_11(dot_0_20_io_b_11),
    .io_b_12(dot_0_20_io_b_12),
    .io_b_13(dot_0_20_io_b_13),
    .io_b_14(dot_0_20_io_b_14),
    .io_b_15(dot_0_20_io_b_15),
    .io_y(dot_0_20_io_y)
  );
  DotProduct dot_0_21 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_21_clock),
    .io_a_0(dot_0_21_io_a_0),
    .io_a_1(dot_0_21_io_a_1),
    .io_a_2(dot_0_21_io_a_2),
    .io_a_3(dot_0_21_io_a_3),
    .io_a_4(dot_0_21_io_a_4),
    .io_a_5(dot_0_21_io_a_5),
    .io_a_6(dot_0_21_io_a_6),
    .io_a_7(dot_0_21_io_a_7),
    .io_a_8(dot_0_21_io_a_8),
    .io_a_9(dot_0_21_io_a_9),
    .io_a_10(dot_0_21_io_a_10),
    .io_a_11(dot_0_21_io_a_11),
    .io_a_12(dot_0_21_io_a_12),
    .io_a_13(dot_0_21_io_a_13),
    .io_a_14(dot_0_21_io_a_14),
    .io_a_15(dot_0_21_io_a_15),
    .io_b_0(dot_0_21_io_b_0),
    .io_b_1(dot_0_21_io_b_1),
    .io_b_2(dot_0_21_io_b_2),
    .io_b_3(dot_0_21_io_b_3),
    .io_b_4(dot_0_21_io_b_4),
    .io_b_5(dot_0_21_io_b_5),
    .io_b_6(dot_0_21_io_b_6),
    .io_b_7(dot_0_21_io_b_7),
    .io_b_8(dot_0_21_io_b_8),
    .io_b_9(dot_0_21_io_b_9),
    .io_b_10(dot_0_21_io_b_10),
    .io_b_11(dot_0_21_io_b_11),
    .io_b_12(dot_0_21_io_b_12),
    .io_b_13(dot_0_21_io_b_13),
    .io_b_14(dot_0_21_io_b_14),
    .io_b_15(dot_0_21_io_b_15),
    .io_y(dot_0_21_io_y)
  );
  DotProduct dot_0_22 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_22_clock),
    .io_a_0(dot_0_22_io_a_0),
    .io_a_1(dot_0_22_io_a_1),
    .io_a_2(dot_0_22_io_a_2),
    .io_a_3(dot_0_22_io_a_3),
    .io_a_4(dot_0_22_io_a_4),
    .io_a_5(dot_0_22_io_a_5),
    .io_a_6(dot_0_22_io_a_6),
    .io_a_7(dot_0_22_io_a_7),
    .io_a_8(dot_0_22_io_a_8),
    .io_a_9(dot_0_22_io_a_9),
    .io_a_10(dot_0_22_io_a_10),
    .io_a_11(dot_0_22_io_a_11),
    .io_a_12(dot_0_22_io_a_12),
    .io_a_13(dot_0_22_io_a_13),
    .io_a_14(dot_0_22_io_a_14),
    .io_a_15(dot_0_22_io_a_15),
    .io_b_0(dot_0_22_io_b_0),
    .io_b_1(dot_0_22_io_b_1),
    .io_b_2(dot_0_22_io_b_2),
    .io_b_3(dot_0_22_io_b_3),
    .io_b_4(dot_0_22_io_b_4),
    .io_b_5(dot_0_22_io_b_5),
    .io_b_6(dot_0_22_io_b_6),
    .io_b_7(dot_0_22_io_b_7),
    .io_b_8(dot_0_22_io_b_8),
    .io_b_9(dot_0_22_io_b_9),
    .io_b_10(dot_0_22_io_b_10),
    .io_b_11(dot_0_22_io_b_11),
    .io_b_12(dot_0_22_io_b_12),
    .io_b_13(dot_0_22_io_b_13),
    .io_b_14(dot_0_22_io_b_14),
    .io_b_15(dot_0_22_io_b_15),
    .io_y(dot_0_22_io_y)
  );
  DotProduct dot_0_23 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_23_clock),
    .io_a_0(dot_0_23_io_a_0),
    .io_a_1(dot_0_23_io_a_1),
    .io_a_2(dot_0_23_io_a_2),
    .io_a_3(dot_0_23_io_a_3),
    .io_a_4(dot_0_23_io_a_4),
    .io_a_5(dot_0_23_io_a_5),
    .io_a_6(dot_0_23_io_a_6),
    .io_a_7(dot_0_23_io_a_7),
    .io_a_8(dot_0_23_io_a_8),
    .io_a_9(dot_0_23_io_a_9),
    .io_a_10(dot_0_23_io_a_10),
    .io_a_11(dot_0_23_io_a_11),
    .io_a_12(dot_0_23_io_a_12),
    .io_a_13(dot_0_23_io_a_13),
    .io_a_14(dot_0_23_io_a_14),
    .io_a_15(dot_0_23_io_a_15),
    .io_b_0(dot_0_23_io_b_0),
    .io_b_1(dot_0_23_io_b_1),
    .io_b_2(dot_0_23_io_b_2),
    .io_b_3(dot_0_23_io_b_3),
    .io_b_4(dot_0_23_io_b_4),
    .io_b_5(dot_0_23_io_b_5),
    .io_b_6(dot_0_23_io_b_6),
    .io_b_7(dot_0_23_io_b_7),
    .io_b_8(dot_0_23_io_b_8),
    .io_b_9(dot_0_23_io_b_9),
    .io_b_10(dot_0_23_io_b_10),
    .io_b_11(dot_0_23_io_b_11),
    .io_b_12(dot_0_23_io_b_12),
    .io_b_13(dot_0_23_io_b_13),
    .io_b_14(dot_0_23_io_b_14),
    .io_b_15(dot_0_23_io_b_15),
    .io_y(dot_0_23_io_y)
  );
  DotProduct dot_0_24 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_24_clock),
    .io_a_0(dot_0_24_io_a_0),
    .io_a_1(dot_0_24_io_a_1),
    .io_a_2(dot_0_24_io_a_2),
    .io_a_3(dot_0_24_io_a_3),
    .io_a_4(dot_0_24_io_a_4),
    .io_a_5(dot_0_24_io_a_5),
    .io_a_6(dot_0_24_io_a_6),
    .io_a_7(dot_0_24_io_a_7),
    .io_a_8(dot_0_24_io_a_8),
    .io_a_9(dot_0_24_io_a_9),
    .io_a_10(dot_0_24_io_a_10),
    .io_a_11(dot_0_24_io_a_11),
    .io_a_12(dot_0_24_io_a_12),
    .io_a_13(dot_0_24_io_a_13),
    .io_a_14(dot_0_24_io_a_14),
    .io_a_15(dot_0_24_io_a_15),
    .io_b_0(dot_0_24_io_b_0),
    .io_b_1(dot_0_24_io_b_1),
    .io_b_2(dot_0_24_io_b_2),
    .io_b_3(dot_0_24_io_b_3),
    .io_b_4(dot_0_24_io_b_4),
    .io_b_5(dot_0_24_io_b_5),
    .io_b_6(dot_0_24_io_b_6),
    .io_b_7(dot_0_24_io_b_7),
    .io_b_8(dot_0_24_io_b_8),
    .io_b_9(dot_0_24_io_b_9),
    .io_b_10(dot_0_24_io_b_10),
    .io_b_11(dot_0_24_io_b_11),
    .io_b_12(dot_0_24_io_b_12),
    .io_b_13(dot_0_24_io_b_13),
    .io_b_14(dot_0_24_io_b_14),
    .io_b_15(dot_0_24_io_b_15),
    .io_y(dot_0_24_io_y)
  );
  DotProduct dot_0_25 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_25_clock),
    .io_a_0(dot_0_25_io_a_0),
    .io_a_1(dot_0_25_io_a_1),
    .io_a_2(dot_0_25_io_a_2),
    .io_a_3(dot_0_25_io_a_3),
    .io_a_4(dot_0_25_io_a_4),
    .io_a_5(dot_0_25_io_a_5),
    .io_a_6(dot_0_25_io_a_6),
    .io_a_7(dot_0_25_io_a_7),
    .io_a_8(dot_0_25_io_a_8),
    .io_a_9(dot_0_25_io_a_9),
    .io_a_10(dot_0_25_io_a_10),
    .io_a_11(dot_0_25_io_a_11),
    .io_a_12(dot_0_25_io_a_12),
    .io_a_13(dot_0_25_io_a_13),
    .io_a_14(dot_0_25_io_a_14),
    .io_a_15(dot_0_25_io_a_15),
    .io_b_0(dot_0_25_io_b_0),
    .io_b_1(dot_0_25_io_b_1),
    .io_b_2(dot_0_25_io_b_2),
    .io_b_3(dot_0_25_io_b_3),
    .io_b_4(dot_0_25_io_b_4),
    .io_b_5(dot_0_25_io_b_5),
    .io_b_6(dot_0_25_io_b_6),
    .io_b_7(dot_0_25_io_b_7),
    .io_b_8(dot_0_25_io_b_8),
    .io_b_9(dot_0_25_io_b_9),
    .io_b_10(dot_0_25_io_b_10),
    .io_b_11(dot_0_25_io_b_11),
    .io_b_12(dot_0_25_io_b_12),
    .io_b_13(dot_0_25_io_b_13),
    .io_b_14(dot_0_25_io_b_14),
    .io_b_15(dot_0_25_io_b_15),
    .io_y(dot_0_25_io_y)
  );
  DotProduct dot_0_26 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_26_clock),
    .io_a_0(dot_0_26_io_a_0),
    .io_a_1(dot_0_26_io_a_1),
    .io_a_2(dot_0_26_io_a_2),
    .io_a_3(dot_0_26_io_a_3),
    .io_a_4(dot_0_26_io_a_4),
    .io_a_5(dot_0_26_io_a_5),
    .io_a_6(dot_0_26_io_a_6),
    .io_a_7(dot_0_26_io_a_7),
    .io_a_8(dot_0_26_io_a_8),
    .io_a_9(dot_0_26_io_a_9),
    .io_a_10(dot_0_26_io_a_10),
    .io_a_11(dot_0_26_io_a_11),
    .io_a_12(dot_0_26_io_a_12),
    .io_a_13(dot_0_26_io_a_13),
    .io_a_14(dot_0_26_io_a_14),
    .io_a_15(dot_0_26_io_a_15),
    .io_b_0(dot_0_26_io_b_0),
    .io_b_1(dot_0_26_io_b_1),
    .io_b_2(dot_0_26_io_b_2),
    .io_b_3(dot_0_26_io_b_3),
    .io_b_4(dot_0_26_io_b_4),
    .io_b_5(dot_0_26_io_b_5),
    .io_b_6(dot_0_26_io_b_6),
    .io_b_7(dot_0_26_io_b_7),
    .io_b_8(dot_0_26_io_b_8),
    .io_b_9(dot_0_26_io_b_9),
    .io_b_10(dot_0_26_io_b_10),
    .io_b_11(dot_0_26_io_b_11),
    .io_b_12(dot_0_26_io_b_12),
    .io_b_13(dot_0_26_io_b_13),
    .io_b_14(dot_0_26_io_b_14),
    .io_b_15(dot_0_26_io_b_15),
    .io_y(dot_0_26_io_y)
  );
  DotProduct dot_0_27 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_27_clock),
    .io_a_0(dot_0_27_io_a_0),
    .io_a_1(dot_0_27_io_a_1),
    .io_a_2(dot_0_27_io_a_2),
    .io_a_3(dot_0_27_io_a_3),
    .io_a_4(dot_0_27_io_a_4),
    .io_a_5(dot_0_27_io_a_5),
    .io_a_6(dot_0_27_io_a_6),
    .io_a_7(dot_0_27_io_a_7),
    .io_a_8(dot_0_27_io_a_8),
    .io_a_9(dot_0_27_io_a_9),
    .io_a_10(dot_0_27_io_a_10),
    .io_a_11(dot_0_27_io_a_11),
    .io_a_12(dot_0_27_io_a_12),
    .io_a_13(dot_0_27_io_a_13),
    .io_a_14(dot_0_27_io_a_14),
    .io_a_15(dot_0_27_io_a_15),
    .io_b_0(dot_0_27_io_b_0),
    .io_b_1(dot_0_27_io_b_1),
    .io_b_2(dot_0_27_io_b_2),
    .io_b_3(dot_0_27_io_b_3),
    .io_b_4(dot_0_27_io_b_4),
    .io_b_5(dot_0_27_io_b_5),
    .io_b_6(dot_0_27_io_b_6),
    .io_b_7(dot_0_27_io_b_7),
    .io_b_8(dot_0_27_io_b_8),
    .io_b_9(dot_0_27_io_b_9),
    .io_b_10(dot_0_27_io_b_10),
    .io_b_11(dot_0_27_io_b_11),
    .io_b_12(dot_0_27_io_b_12),
    .io_b_13(dot_0_27_io_b_13),
    .io_b_14(dot_0_27_io_b_14),
    .io_b_15(dot_0_27_io_b_15),
    .io_y(dot_0_27_io_y)
  );
  DotProduct dot_0_28 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_28_clock),
    .io_a_0(dot_0_28_io_a_0),
    .io_a_1(dot_0_28_io_a_1),
    .io_a_2(dot_0_28_io_a_2),
    .io_a_3(dot_0_28_io_a_3),
    .io_a_4(dot_0_28_io_a_4),
    .io_a_5(dot_0_28_io_a_5),
    .io_a_6(dot_0_28_io_a_6),
    .io_a_7(dot_0_28_io_a_7),
    .io_a_8(dot_0_28_io_a_8),
    .io_a_9(dot_0_28_io_a_9),
    .io_a_10(dot_0_28_io_a_10),
    .io_a_11(dot_0_28_io_a_11),
    .io_a_12(dot_0_28_io_a_12),
    .io_a_13(dot_0_28_io_a_13),
    .io_a_14(dot_0_28_io_a_14),
    .io_a_15(dot_0_28_io_a_15),
    .io_b_0(dot_0_28_io_b_0),
    .io_b_1(dot_0_28_io_b_1),
    .io_b_2(dot_0_28_io_b_2),
    .io_b_3(dot_0_28_io_b_3),
    .io_b_4(dot_0_28_io_b_4),
    .io_b_5(dot_0_28_io_b_5),
    .io_b_6(dot_0_28_io_b_6),
    .io_b_7(dot_0_28_io_b_7),
    .io_b_8(dot_0_28_io_b_8),
    .io_b_9(dot_0_28_io_b_9),
    .io_b_10(dot_0_28_io_b_10),
    .io_b_11(dot_0_28_io_b_11),
    .io_b_12(dot_0_28_io_b_12),
    .io_b_13(dot_0_28_io_b_13),
    .io_b_14(dot_0_28_io_b_14),
    .io_b_15(dot_0_28_io_b_15),
    .io_y(dot_0_28_io_y)
  );
  DotProduct dot_0_29 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_29_clock),
    .io_a_0(dot_0_29_io_a_0),
    .io_a_1(dot_0_29_io_a_1),
    .io_a_2(dot_0_29_io_a_2),
    .io_a_3(dot_0_29_io_a_3),
    .io_a_4(dot_0_29_io_a_4),
    .io_a_5(dot_0_29_io_a_5),
    .io_a_6(dot_0_29_io_a_6),
    .io_a_7(dot_0_29_io_a_7),
    .io_a_8(dot_0_29_io_a_8),
    .io_a_9(dot_0_29_io_a_9),
    .io_a_10(dot_0_29_io_a_10),
    .io_a_11(dot_0_29_io_a_11),
    .io_a_12(dot_0_29_io_a_12),
    .io_a_13(dot_0_29_io_a_13),
    .io_a_14(dot_0_29_io_a_14),
    .io_a_15(dot_0_29_io_a_15),
    .io_b_0(dot_0_29_io_b_0),
    .io_b_1(dot_0_29_io_b_1),
    .io_b_2(dot_0_29_io_b_2),
    .io_b_3(dot_0_29_io_b_3),
    .io_b_4(dot_0_29_io_b_4),
    .io_b_5(dot_0_29_io_b_5),
    .io_b_6(dot_0_29_io_b_6),
    .io_b_7(dot_0_29_io_b_7),
    .io_b_8(dot_0_29_io_b_8),
    .io_b_9(dot_0_29_io_b_9),
    .io_b_10(dot_0_29_io_b_10),
    .io_b_11(dot_0_29_io_b_11),
    .io_b_12(dot_0_29_io_b_12),
    .io_b_13(dot_0_29_io_b_13),
    .io_b_14(dot_0_29_io_b_14),
    .io_b_15(dot_0_29_io_b_15),
    .io_y(dot_0_29_io_y)
  );
  DotProduct dot_0_30 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_30_clock),
    .io_a_0(dot_0_30_io_a_0),
    .io_a_1(dot_0_30_io_a_1),
    .io_a_2(dot_0_30_io_a_2),
    .io_a_3(dot_0_30_io_a_3),
    .io_a_4(dot_0_30_io_a_4),
    .io_a_5(dot_0_30_io_a_5),
    .io_a_6(dot_0_30_io_a_6),
    .io_a_7(dot_0_30_io_a_7),
    .io_a_8(dot_0_30_io_a_8),
    .io_a_9(dot_0_30_io_a_9),
    .io_a_10(dot_0_30_io_a_10),
    .io_a_11(dot_0_30_io_a_11),
    .io_a_12(dot_0_30_io_a_12),
    .io_a_13(dot_0_30_io_a_13),
    .io_a_14(dot_0_30_io_a_14),
    .io_a_15(dot_0_30_io_a_15),
    .io_b_0(dot_0_30_io_b_0),
    .io_b_1(dot_0_30_io_b_1),
    .io_b_2(dot_0_30_io_b_2),
    .io_b_3(dot_0_30_io_b_3),
    .io_b_4(dot_0_30_io_b_4),
    .io_b_5(dot_0_30_io_b_5),
    .io_b_6(dot_0_30_io_b_6),
    .io_b_7(dot_0_30_io_b_7),
    .io_b_8(dot_0_30_io_b_8),
    .io_b_9(dot_0_30_io_b_9),
    .io_b_10(dot_0_30_io_b_10),
    .io_b_11(dot_0_30_io_b_11),
    .io_b_12(dot_0_30_io_b_12),
    .io_b_13(dot_0_30_io_b_13),
    .io_b_14(dot_0_30_io_b_14),
    .io_b_15(dot_0_30_io_b_15),
    .io_y(dot_0_30_io_y)
  );
  DotProduct dot_0_31 ( // @[TensorGemm.scala 198:11]
    .clock(dot_0_31_clock),
    .io_a_0(dot_0_31_io_a_0),
    .io_a_1(dot_0_31_io_a_1),
    .io_a_2(dot_0_31_io_a_2),
    .io_a_3(dot_0_31_io_a_3),
    .io_a_4(dot_0_31_io_a_4),
    .io_a_5(dot_0_31_io_a_5),
    .io_a_6(dot_0_31_io_a_6),
    .io_a_7(dot_0_31_io_a_7),
    .io_a_8(dot_0_31_io_a_8),
    .io_a_9(dot_0_31_io_a_9),
    .io_a_10(dot_0_31_io_a_10),
    .io_a_11(dot_0_31_io_a_11),
    .io_a_12(dot_0_31_io_a_12),
    .io_a_13(dot_0_31_io_a_13),
    .io_a_14(dot_0_31_io_a_14),
    .io_a_15(dot_0_31_io_a_15),
    .io_b_0(dot_0_31_io_b_0),
    .io_b_1(dot_0_31_io_b_1),
    .io_b_2(dot_0_31_io_b_2),
    .io_b_3(dot_0_31_io_b_3),
    .io_b_4(dot_0_31_io_b_4),
    .io_b_5(dot_0_31_io_b_5),
    .io_b_6(dot_0_31_io_b_6),
    .io_b_7(dot_0_31_io_b_7),
    .io_b_8(dot_0_31_io_b_8),
    .io_b_9(dot_0_31_io_b_9),
    .io_b_10(dot_0_31_io_b_10),
    .io_b_11(dot_0_31_io_b_11),
    .io_b_12(dot_0_31_io_b_12),
    .io_b_13(dot_0_31_io_b_13),
    .io_b_14(dot_0_31_io_b_14),
    .io_b_15(dot_0_31_io_b_15),
    .io_y(dot_0_31_io_y)
  );
  assign io_acc_o_data_valid = io_acc_i_data_valid | io_valid_reset; // @[TensorGemm.scala 216:46]
  assign io_acc_o_data_bits_0_0 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_0); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_1 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_1); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_2 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_2); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_3 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_3); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_4 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_4); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_5 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_5); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_6 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_6); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_7 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_7); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_8 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_8); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_9 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_9); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_10 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_10); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_11 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_11); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_12 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_12); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_13 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_13); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_14 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_14); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_15 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_15); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_16 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_16); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_17 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_17); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_18 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_18); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_19 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_19); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_20 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_20); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_21 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_21); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_22 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_22); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_23 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_23); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_24 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_24); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_25 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_25); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_26 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_26); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_27 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_27); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_28 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_28); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_29 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_29); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_30 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_30); // @[TensorGemm.scala 211:39]
  assign io_acc_o_data_bits_0_31 = io_valid_reset ? $signed(32'sh0) : $signed(add_0_31); // @[TensorGemm.scala 211:39]
  assign io_out_data_valid = io_acc_i_data_valid & ~io_valid_reset; // @[TensorGemm.scala 217:44]
  assign io_out_data_bits_0_0 = _io_out_data_bits_0_0_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_1 = _io_out_data_bits_0_1_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_2 = _io_out_data_bits_0_2_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_3 = _io_out_data_bits_0_3_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_4 = _io_out_data_bits_0_4_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_5 = _io_out_data_bits_0_5_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_6 = _io_out_data_bits_0_6_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_7 = _io_out_data_bits_0_7_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_8 = _io_out_data_bits_0_8_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_9 = _io_out_data_bits_0_9_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_10 = _io_out_data_bits_0_10_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_11 = _io_out_data_bits_0_11_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_12 = _io_out_data_bits_0_12_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_13 = _io_out_data_bits_0_13_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_14 = _io_out_data_bits_0_14_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_15 = _io_out_data_bits_0_15_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_16 = _io_out_data_bits_0_16_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_17 = _io_out_data_bits_0_17_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_18 = _io_out_data_bits_0_18_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_19 = _io_out_data_bits_0_19_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_20 = _io_out_data_bits_0_20_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_21 = _io_out_data_bits_0_21_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_22 = _io_out_data_bits_0_22_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_23 = _io_out_data_bits_0_23_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_24 = _io_out_data_bits_0_24_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_25 = _io_out_data_bits_0_25_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_26 = _io_out_data_bits_0_26_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_27 = _io_out_data_bits_0_27_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_28 = _io_out_data_bits_0_28_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_29 = _io_out_data_bits_0_29_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_30 = _io_out_data_bits_0_30_T[7:0]; // @[TensorGemm.scala 213:30]
  assign io_out_data_bits_0_31 = _io_out_data_bits_0_31_T[7:0]; // @[TensorGemm.scala 213:30]
  assign dot_0_0_clock = clock;
  assign dot_0_0_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_0_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_0_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_0_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_0_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_0_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_0_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_0_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_0_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_0_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_0_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_0_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_0_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_0_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_0_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_0_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_0_io_b_0 = io_wgt_data_bits_0_0; // @[TensorGemm.scala 206:53]
  assign dot_0_0_io_b_1 = io_wgt_data_bits_0_1; // @[TensorGemm.scala 206:53]
  assign dot_0_0_io_b_2 = io_wgt_data_bits_0_2; // @[TensorGemm.scala 206:53]
  assign dot_0_0_io_b_3 = io_wgt_data_bits_0_3; // @[TensorGemm.scala 206:53]
  assign dot_0_0_io_b_4 = io_wgt_data_bits_0_4; // @[TensorGemm.scala 206:53]
  assign dot_0_0_io_b_5 = io_wgt_data_bits_0_5; // @[TensorGemm.scala 206:53]
  assign dot_0_0_io_b_6 = io_wgt_data_bits_0_6; // @[TensorGemm.scala 206:53]
  assign dot_0_0_io_b_7 = io_wgt_data_bits_0_7; // @[TensorGemm.scala 206:53]
  assign dot_0_0_io_b_8 = io_wgt_data_bits_0_8; // @[TensorGemm.scala 206:53]
  assign dot_0_0_io_b_9 = io_wgt_data_bits_0_9; // @[TensorGemm.scala 206:53]
  assign dot_0_0_io_b_10 = io_wgt_data_bits_0_10; // @[TensorGemm.scala 206:53]
  assign dot_0_0_io_b_11 = io_wgt_data_bits_0_11; // @[TensorGemm.scala 206:53]
  assign dot_0_0_io_b_12 = io_wgt_data_bits_0_12; // @[TensorGemm.scala 206:53]
  assign dot_0_0_io_b_13 = io_wgt_data_bits_0_13; // @[TensorGemm.scala 206:53]
  assign dot_0_0_io_b_14 = io_wgt_data_bits_0_14; // @[TensorGemm.scala 206:53]
  assign dot_0_0_io_b_15 = io_wgt_data_bits_0_15; // @[TensorGemm.scala 206:53]
  assign dot_0_1_clock = clock;
  assign dot_0_1_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_1_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_1_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_1_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_1_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_1_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_1_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_1_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_1_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_1_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_1_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_1_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_1_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_1_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_1_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_1_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_1_io_b_0 = io_wgt_data_bits_1_0; // @[TensorGemm.scala 206:53]
  assign dot_0_1_io_b_1 = io_wgt_data_bits_1_1; // @[TensorGemm.scala 206:53]
  assign dot_0_1_io_b_2 = io_wgt_data_bits_1_2; // @[TensorGemm.scala 206:53]
  assign dot_0_1_io_b_3 = io_wgt_data_bits_1_3; // @[TensorGemm.scala 206:53]
  assign dot_0_1_io_b_4 = io_wgt_data_bits_1_4; // @[TensorGemm.scala 206:53]
  assign dot_0_1_io_b_5 = io_wgt_data_bits_1_5; // @[TensorGemm.scala 206:53]
  assign dot_0_1_io_b_6 = io_wgt_data_bits_1_6; // @[TensorGemm.scala 206:53]
  assign dot_0_1_io_b_7 = io_wgt_data_bits_1_7; // @[TensorGemm.scala 206:53]
  assign dot_0_1_io_b_8 = io_wgt_data_bits_1_8; // @[TensorGemm.scala 206:53]
  assign dot_0_1_io_b_9 = io_wgt_data_bits_1_9; // @[TensorGemm.scala 206:53]
  assign dot_0_1_io_b_10 = io_wgt_data_bits_1_10; // @[TensorGemm.scala 206:53]
  assign dot_0_1_io_b_11 = io_wgt_data_bits_1_11; // @[TensorGemm.scala 206:53]
  assign dot_0_1_io_b_12 = io_wgt_data_bits_1_12; // @[TensorGemm.scala 206:53]
  assign dot_0_1_io_b_13 = io_wgt_data_bits_1_13; // @[TensorGemm.scala 206:53]
  assign dot_0_1_io_b_14 = io_wgt_data_bits_1_14; // @[TensorGemm.scala 206:53]
  assign dot_0_1_io_b_15 = io_wgt_data_bits_1_15; // @[TensorGemm.scala 206:53]
  assign dot_0_2_clock = clock;
  assign dot_0_2_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_2_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_2_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_2_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_2_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_2_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_2_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_2_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_2_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_2_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_2_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_2_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_2_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_2_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_2_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_2_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_2_io_b_0 = io_wgt_data_bits_2_0; // @[TensorGemm.scala 206:53]
  assign dot_0_2_io_b_1 = io_wgt_data_bits_2_1; // @[TensorGemm.scala 206:53]
  assign dot_0_2_io_b_2 = io_wgt_data_bits_2_2; // @[TensorGemm.scala 206:53]
  assign dot_0_2_io_b_3 = io_wgt_data_bits_2_3; // @[TensorGemm.scala 206:53]
  assign dot_0_2_io_b_4 = io_wgt_data_bits_2_4; // @[TensorGemm.scala 206:53]
  assign dot_0_2_io_b_5 = io_wgt_data_bits_2_5; // @[TensorGemm.scala 206:53]
  assign dot_0_2_io_b_6 = io_wgt_data_bits_2_6; // @[TensorGemm.scala 206:53]
  assign dot_0_2_io_b_7 = io_wgt_data_bits_2_7; // @[TensorGemm.scala 206:53]
  assign dot_0_2_io_b_8 = io_wgt_data_bits_2_8; // @[TensorGemm.scala 206:53]
  assign dot_0_2_io_b_9 = io_wgt_data_bits_2_9; // @[TensorGemm.scala 206:53]
  assign dot_0_2_io_b_10 = io_wgt_data_bits_2_10; // @[TensorGemm.scala 206:53]
  assign dot_0_2_io_b_11 = io_wgt_data_bits_2_11; // @[TensorGemm.scala 206:53]
  assign dot_0_2_io_b_12 = io_wgt_data_bits_2_12; // @[TensorGemm.scala 206:53]
  assign dot_0_2_io_b_13 = io_wgt_data_bits_2_13; // @[TensorGemm.scala 206:53]
  assign dot_0_2_io_b_14 = io_wgt_data_bits_2_14; // @[TensorGemm.scala 206:53]
  assign dot_0_2_io_b_15 = io_wgt_data_bits_2_15; // @[TensorGemm.scala 206:53]
  assign dot_0_3_clock = clock;
  assign dot_0_3_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_3_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_3_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_3_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_3_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_3_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_3_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_3_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_3_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_3_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_3_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_3_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_3_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_3_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_3_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_3_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_3_io_b_0 = io_wgt_data_bits_3_0; // @[TensorGemm.scala 206:53]
  assign dot_0_3_io_b_1 = io_wgt_data_bits_3_1; // @[TensorGemm.scala 206:53]
  assign dot_0_3_io_b_2 = io_wgt_data_bits_3_2; // @[TensorGemm.scala 206:53]
  assign dot_0_3_io_b_3 = io_wgt_data_bits_3_3; // @[TensorGemm.scala 206:53]
  assign dot_0_3_io_b_4 = io_wgt_data_bits_3_4; // @[TensorGemm.scala 206:53]
  assign dot_0_3_io_b_5 = io_wgt_data_bits_3_5; // @[TensorGemm.scala 206:53]
  assign dot_0_3_io_b_6 = io_wgt_data_bits_3_6; // @[TensorGemm.scala 206:53]
  assign dot_0_3_io_b_7 = io_wgt_data_bits_3_7; // @[TensorGemm.scala 206:53]
  assign dot_0_3_io_b_8 = io_wgt_data_bits_3_8; // @[TensorGemm.scala 206:53]
  assign dot_0_3_io_b_9 = io_wgt_data_bits_3_9; // @[TensorGemm.scala 206:53]
  assign dot_0_3_io_b_10 = io_wgt_data_bits_3_10; // @[TensorGemm.scala 206:53]
  assign dot_0_3_io_b_11 = io_wgt_data_bits_3_11; // @[TensorGemm.scala 206:53]
  assign dot_0_3_io_b_12 = io_wgt_data_bits_3_12; // @[TensorGemm.scala 206:53]
  assign dot_0_3_io_b_13 = io_wgt_data_bits_3_13; // @[TensorGemm.scala 206:53]
  assign dot_0_3_io_b_14 = io_wgt_data_bits_3_14; // @[TensorGemm.scala 206:53]
  assign dot_0_3_io_b_15 = io_wgt_data_bits_3_15; // @[TensorGemm.scala 206:53]
  assign dot_0_4_clock = clock;
  assign dot_0_4_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_4_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_4_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_4_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_4_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_4_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_4_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_4_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_4_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_4_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_4_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_4_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_4_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_4_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_4_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_4_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_4_io_b_0 = io_wgt_data_bits_4_0; // @[TensorGemm.scala 206:53]
  assign dot_0_4_io_b_1 = io_wgt_data_bits_4_1; // @[TensorGemm.scala 206:53]
  assign dot_0_4_io_b_2 = io_wgt_data_bits_4_2; // @[TensorGemm.scala 206:53]
  assign dot_0_4_io_b_3 = io_wgt_data_bits_4_3; // @[TensorGemm.scala 206:53]
  assign dot_0_4_io_b_4 = io_wgt_data_bits_4_4; // @[TensorGemm.scala 206:53]
  assign dot_0_4_io_b_5 = io_wgt_data_bits_4_5; // @[TensorGemm.scala 206:53]
  assign dot_0_4_io_b_6 = io_wgt_data_bits_4_6; // @[TensorGemm.scala 206:53]
  assign dot_0_4_io_b_7 = io_wgt_data_bits_4_7; // @[TensorGemm.scala 206:53]
  assign dot_0_4_io_b_8 = io_wgt_data_bits_4_8; // @[TensorGemm.scala 206:53]
  assign dot_0_4_io_b_9 = io_wgt_data_bits_4_9; // @[TensorGemm.scala 206:53]
  assign dot_0_4_io_b_10 = io_wgt_data_bits_4_10; // @[TensorGemm.scala 206:53]
  assign dot_0_4_io_b_11 = io_wgt_data_bits_4_11; // @[TensorGemm.scala 206:53]
  assign dot_0_4_io_b_12 = io_wgt_data_bits_4_12; // @[TensorGemm.scala 206:53]
  assign dot_0_4_io_b_13 = io_wgt_data_bits_4_13; // @[TensorGemm.scala 206:53]
  assign dot_0_4_io_b_14 = io_wgt_data_bits_4_14; // @[TensorGemm.scala 206:53]
  assign dot_0_4_io_b_15 = io_wgt_data_bits_4_15; // @[TensorGemm.scala 206:53]
  assign dot_0_5_clock = clock;
  assign dot_0_5_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_5_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_5_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_5_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_5_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_5_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_5_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_5_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_5_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_5_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_5_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_5_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_5_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_5_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_5_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_5_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_5_io_b_0 = io_wgt_data_bits_5_0; // @[TensorGemm.scala 206:53]
  assign dot_0_5_io_b_1 = io_wgt_data_bits_5_1; // @[TensorGemm.scala 206:53]
  assign dot_0_5_io_b_2 = io_wgt_data_bits_5_2; // @[TensorGemm.scala 206:53]
  assign dot_0_5_io_b_3 = io_wgt_data_bits_5_3; // @[TensorGemm.scala 206:53]
  assign dot_0_5_io_b_4 = io_wgt_data_bits_5_4; // @[TensorGemm.scala 206:53]
  assign dot_0_5_io_b_5 = io_wgt_data_bits_5_5; // @[TensorGemm.scala 206:53]
  assign dot_0_5_io_b_6 = io_wgt_data_bits_5_6; // @[TensorGemm.scala 206:53]
  assign dot_0_5_io_b_7 = io_wgt_data_bits_5_7; // @[TensorGemm.scala 206:53]
  assign dot_0_5_io_b_8 = io_wgt_data_bits_5_8; // @[TensorGemm.scala 206:53]
  assign dot_0_5_io_b_9 = io_wgt_data_bits_5_9; // @[TensorGemm.scala 206:53]
  assign dot_0_5_io_b_10 = io_wgt_data_bits_5_10; // @[TensorGemm.scala 206:53]
  assign dot_0_5_io_b_11 = io_wgt_data_bits_5_11; // @[TensorGemm.scala 206:53]
  assign dot_0_5_io_b_12 = io_wgt_data_bits_5_12; // @[TensorGemm.scala 206:53]
  assign dot_0_5_io_b_13 = io_wgt_data_bits_5_13; // @[TensorGemm.scala 206:53]
  assign dot_0_5_io_b_14 = io_wgt_data_bits_5_14; // @[TensorGemm.scala 206:53]
  assign dot_0_5_io_b_15 = io_wgt_data_bits_5_15; // @[TensorGemm.scala 206:53]
  assign dot_0_6_clock = clock;
  assign dot_0_6_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_6_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_6_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_6_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_6_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_6_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_6_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_6_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_6_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_6_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_6_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_6_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_6_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_6_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_6_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_6_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_6_io_b_0 = io_wgt_data_bits_6_0; // @[TensorGemm.scala 206:53]
  assign dot_0_6_io_b_1 = io_wgt_data_bits_6_1; // @[TensorGemm.scala 206:53]
  assign dot_0_6_io_b_2 = io_wgt_data_bits_6_2; // @[TensorGemm.scala 206:53]
  assign dot_0_6_io_b_3 = io_wgt_data_bits_6_3; // @[TensorGemm.scala 206:53]
  assign dot_0_6_io_b_4 = io_wgt_data_bits_6_4; // @[TensorGemm.scala 206:53]
  assign dot_0_6_io_b_5 = io_wgt_data_bits_6_5; // @[TensorGemm.scala 206:53]
  assign dot_0_6_io_b_6 = io_wgt_data_bits_6_6; // @[TensorGemm.scala 206:53]
  assign dot_0_6_io_b_7 = io_wgt_data_bits_6_7; // @[TensorGemm.scala 206:53]
  assign dot_0_6_io_b_8 = io_wgt_data_bits_6_8; // @[TensorGemm.scala 206:53]
  assign dot_0_6_io_b_9 = io_wgt_data_bits_6_9; // @[TensorGemm.scala 206:53]
  assign dot_0_6_io_b_10 = io_wgt_data_bits_6_10; // @[TensorGemm.scala 206:53]
  assign dot_0_6_io_b_11 = io_wgt_data_bits_6_11; // @[TensorGemm.scala 206:53]
  assign dot_0_6_io_b_12 = io_wgt_data_bits_6_12; // @[TensorGemm.scala 206:53]
  assign dot_0_6_io_b_13 = io_wgt_data_bits_6_13; // @[TensorGemm.scala 206:53]
  assign dot_0_6_io_b_14 = io_wgt_data_bits_6_14; // @[TensorGemm.scala 206:53]
  assign dot_0_6_io_b_15 = io_wgt_data_bits_6_15; // @[TensorGemm.scala 206:53]
  assign dot_0_7_clock = clock;
  assign dot_0_7_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_7_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_7_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_7_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_7_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_7_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_7_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_7_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_7_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_7_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_7_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_7_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_7_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_7_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_7_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_7_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_7_io_b_0 = io_wgt_data_bits_7_0; // @[TensorGemm.scala 206:53]
  assign dot_0_7_io_b_1 = io_wgt_data_bits_7_1; // @[TensorGemm.scala 206:53]
  assign dot_0_7_io_b_2 = io_wgt_data_bits_7_2; // @[TensorGemm.scala 206:53]
  assign dot_0_7_io_b_3 = io_wgt_data_bits_7_3; // @[TensorGemm.scala 206:53]
  assign dot_0_7_io_b_4 = io_wgt_data_bits_7_4; // @[TensorGemm.scala 206:53]
  assign dot_0_7_io_b_5 = io_wgt_data_bits_7_5; // @[TensorGemm.scala 206:53]
  assign dot_0_7_io_b_6 = io_wgt_data_bits_7_6; // @[TensorGemm.scala 206:53]
  assign dot_0_7_io_b_7 = io_wgt_data_bits_7_7; // @[TensorGemm.scala 206:53]
  assign dot_0_7_io_b_8 = io_wgt_data_bits_7_8; // @[TensorGemm.scala 206:53]
  assign dot_0_7_io_b_9 = io_wgt_data_bits_7_9; // @[TensorGemm.scala 206:53]
  assign dot_0_7_io_b_10 = io_wgt_data_bits_7_10; // @[TensorGemm.scala 206:53]
  assign dot_0_7_io_b_11 = io_wgt_data_bits_7_11; // @[TensorGemm.scala 206:53]
  assign dot_0_7_io_b_12 = io_wgt_data_bits_7_12; // @[TensorGemm.scala 206:53]
  assign dot_0_7_io_b_13 = io_wgt_data_bits_7_13; // @[TensorGemm.scala 206:53]
  assign dot_0_7_io_b_14 = io_wgt_data_bits_7_14; // @[TensorGemm.scala 206:53]
  assign dot_0_7_io_b_15 = io_wgt_data_bits_7_15; // @[TensorGemm.scala 206:53]
  assign dot_0_8_clock = clock;
  assign dot_0_8_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_8_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_8_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_8_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_8_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_8_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_8_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_8_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_8_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_8_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_8_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_8_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_8_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_8_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_8_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_8_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_8_io_b_0 = io_wgt_data_bits_8_0; // @[TensorGemm.scala 206:53]
  assign dot_0_8_io_b_1 = io_wgt_data_bits_8_1; // @[TensorGemm.scala 206:53]
  assign dot_0_8_io_b_2 = io_wgt_data_bits_8_2; // @[TensorGemm.scala 206:53]
  assign dot_0_8_io_b_3 = io_wgt_data_bits_8_3; // @[TensorGemm.scala 206:53]
  assign dot_0_8_io_b_4 = io_wgt_data_bits_8_4; // @[TensorGemm.scala 206:53]
  assign dot_0_8_io_b_5 = io_wgt_data_bits_8_5; // @[TensorGemm.scala 206:53]
  assign dot_0_8_io_b_6 = io_wgt_data_bits_8_6; // @[TensorGemm.scala 206:53]
  assign dot_0_8_io_b_7 = io_wgt_data_bits_8_7; // @[TensorGemm.scala 206:53]
  assign dot_0_8_io_b_8 = io_wgt_data_bits_8_8; // @[TensorGemm.scala 206:53]
  assign dot_0_8_io_b_9 = io_wgt_data_bits_8_9; // @[TensorGemm.scala 206:53]
  assign dot_0_8_io_b_10 = io_wgt_data_bits_8_10; // @[TensorGemm.scala 206:53]
  assign dot_0_8_io_b_11 = io_wgt_data_bits_8_11; // @[TensorGemm.scala 206:53]
  assign dot_0_8_io_b_12 = io_wgt_data_bits_8_12; // @[TensorGemm.scala 206:53]
  assign dot_0_8_io_b_13 = io_wgt_data_bits_8_13; // @[TensorGemm.scala 206:53]
  assign dot_0_8_io_b_14 = io_wgt_data_bits_8_14; // @[TensorGemm.scala 206:53]
  assign dot_0_8_io_b_15 = io_wgt_data_bits_8_15; // @[TensorGemm.scala 206:53]
  assign dot_0_9_clock = clock;
  assign dot_0_9_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_9_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_9_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_9_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_9_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_9_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_9_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_9_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_9_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_9_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_9_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_9_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_9_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_9_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_9_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_9_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_9_io_b_0 = io_wgt_data_bits_9_0; // @[TensorGemm.scala 206:53]
  assign dot_0_9_io_b_1 = io_wgt_data_bits_9_1; // @[TensorGemm.scala 206:53]
  assign dot_0_9_io_b_2 = io_wgt_data_bits_9_2; // @[TensorGemm.scala 206:53]
  assign dot_0_9_io_b_3 = io_wgt_data_bits_9_3; // @[TensorGemm.scala 206:53]
  assign dot_0_9_io_b_4 = io_wgt_data_bits_9_4; // @[TensorGemm.scala 206:53]
  assign dot_0_9_io_b_5 = io_wgt_data_bits_9_5; // @[TensorGemm.scala 206:53]
  assign dot_0_9_io_b_6 = io_wgt_data_bits_9_6; // @[TensorGemm.scala 206:53]
  assign dot_0_9_io_b_7 = io_wgt_data_bits_9_7; // @[TensorGemm.scala 206:53]
  assign dot_0_9_io_b_8 = io_wgt_data_bits_9_8; // @[TensorGemm.scala 206:53]
  assign dot_0_9_io_b_9 = io_wgt_data_bits_9_9; // @[TensorGemm.scala 206:53]
  assign dot_0_9_io_b_10 = io_wgt_data_bits_9_10; // @[TensorGemm.scala 206:53]
  assign dot_0_9_io_b_11 = io_wgt_data_bits_9_11; // @[TensorGemm.scala 206:53]
  assign dot_0_9_io_b_12 = io_wgt_data_bits_9_12; // @[TensorGemm.scala 206:53]
  assign dot_0_9_io_b_13 = io_wgt_data_bits_9_13; // @[TensorGemm.scala 206:53]
  assign dot_0_9_io_b_14 = io_wgt_data_bits_9_14; // @[TensorGemm.scala 206:53]
  assign dot_0_9_io_b_15 = io_wgt_data_bits_9_15; // @[TensorGemm.scala 206:53]
  assign dot_0_10_clock = clock;
  assign dot_0_10_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_10_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_10_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_10_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_10_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_10_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_10_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_10_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_10_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_10_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_10_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_10_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_10_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_10_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_10_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_10_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_10_io_b_0 = io_wgt_data_bits_10_0; // @[TensorGemm.scala 206:53]
  assign dot_0_10_io_b_1 = io_wgt_data_bits_10_1; // @[TensorGemm.scala 206:53]
  assign dot_0_10_io_b_2 = io_wgt_data_bits_10_2; // @[TensorGemm.scala 206:53]
  assign dot_0_10_io_b_3 = io_wgt_data_bits_10_3; // @[TensorGemm.scala 206:53]
  assign dot_0_10_io_b_4 = io_wgt_data_bits_10_4; // @[TensorGemm.scala 206:53]
  assign dot_0_10_io_b_5 = io_wgt_data_bits_10_5; // @[TensorGemm.scala 206:53]
  assign dot_0_10_io_b_6 = io_wgt_data_bits_10_6; // @[TensorGemm.scala 206:53]
  assign dot_0_10_io_b_7 = io_wgt_data_bits_10_7; // @[TensorGemm.scala 206:53]
  assign dot_0_10_io_b_8 = io_wgt_data_bits_10_8; // @[TensorGemm.scala 206:53]
  assign dot_0_10_io_b_9 = io_wgt_data_bits_10_9; // @[TensorGemm.scala 206:53]
  assign dot_0_10_io_b_10 = io_wgt_data_bits_10_10; // @[TensorGemm.scala 206:53]
  assign dot_0_10_io_b_11 = io_wgt_data_bits_10_11; // @[TensorGemm.scala 206:53]
  assign dot_0_10_io_b_12 = io_wgt_data_bits_10_12; // @[TensorGemm.scala 206:53]
  assign dot_0_10_io_b_13 = io_wgt_data_bits_10_13; // @[TensorGemm.scala 206:53]
  assign dot_0_10_io_b_14 = io_wgt_data_bits_10_14; // @[TensorGemm.scala 206:53]
  assign dot_0_10_io_b_15 = io_wgt_data_bits_10_15; // @[TensorGemm.scala 206:53]
  assign dot_0_11_clock = clock;
  assign dot_0_11_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_11_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_11_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_11_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_11_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_11_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_11_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_11_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_11_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_11_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_11_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_11_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_11_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_11_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_11_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_11_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_11_io_b_0 = io_wgt_data_bits_11_0; // @[TensorGemm.scala 206:53]
  assign dot_0_11_io_b_1 = io_wgt_data_bits_11_1; // @[TensorGemm.scala 206:53]
  assign dot_0_11_io_b_2 = io_wgt_data_bits_11_2; // @[TensorGemm.scala 206:53]
  assign dot_0_11_io_b_3 = io_wgt_data_bits_11_3; // @[TensorGemm.scala 206:53]
  assign dot_0_11_io_b_4 = io_wgt_data_bits_11_4; // @[TensorGemm.scala 206:53]
  assign dot_0_11_io_b_5 = io_wgt_data_bits_11_5; // @[TensorGemm.scala 206:53]
  assign dot_0_11_io_b_6 = io_wgt_data_bits_11_6; // @[TensorGemm.scala 206:53]
  assign dot_0_11_io_b_7 = io_wgt_data_bits_11_7; // @[TensorGemm.scala 206:53]
  assign dot_0_11_io_b_8 = io_wgt_data_bits_11_8; // @[TensorGemm.scala 206:53]
  assign dot_0_11_io_b_9 = io_wgt_data_bits_11_9; // @[TensorGemm.scala 206:53]
  assign dot_0_11_io_b_10 = io_wgt_data_bits_11_10; // @[TensorGemm.scala 206:53]
  assign dot_0_11_io_b_11 = io_wgt_data_bits_11_11; // @[TensorGemm.scala 206:53]
  assign dot_0_11_io_b_12 = io_wgt_data_bits_11_12; // @[TensorGemm.scala 206:53]
  assign dot_0_11_io_b_13 = io_wgt_data_bits_11_13; // @[TensorGemm.scala 206:53]
  assign dot_0_11_io_b_14 = io_wgt_data_bits_11_14; // @[TensorGemm.scala 206:53]
  assign dot_0_11_io_b_15 = io_wgt_data_bits_11_15; // @[TensorGemm.scala 206:53]
  assign dot_0_12_clock = clock;
  assign dot_0_12_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_12_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_12_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_12_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_12_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_12_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_12_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_12_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_12_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_12_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_12_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_12_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_12_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_12_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_12_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_12_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_12_io_b_0 = io_wgt_data_bits_12_0; // @[TensorGemm.scala 206:53]
  assign dot_0_12_io_b_1 = io_wgt_data_bits_12_1; // @[TensorGemm.scala 206:53]
  assign dot_0_12_io_b_2 = io_wgt_data_bits_12_2; // @[TensorGemm.scala 206:53]
  assign dot_0_12_io_b_3 = io_wgt_data_bits_12_3; // @[TensorGemm.scala 206:53]
  assign dot_0_12_io_b_4 = io_wgt_data_bits_12_4; // @[TensorGemm.scala 206:53]
  assign dot_0_12_io_b_5 = io_wgt_data_bits_12_5; // @[TensorGemm.scala 206:53]
  assign dot_0_12_io_b_6 = io_wgt_data_bits_12_6; // @[TensorGemm.scala 206:53]
  assign dot_0_12_io_b_7 = io_wgt_data_bits_12_7; // @[TensorGemm.scala 206:53]
  assign dot_0_12_io_b_8 = io_wgt_data_bits_12_8; // @[TensorGemm.scala 206:53]
  assign dot_0_12_io_b_9 = io_wgt_data_bits_12_9; // @[TensorGemm.scala 206:53]
  assign dot_0_12_io_b_10 = io_wgt_data_bits_12_10; // @[TensorGemm.scala 206:53]
  assign dot_0_12_io_b_11 = io_wgt_data_bits_12_11; // @[TensorGemm.scala 206:53]
  assign dot_0_12_io_b_12 = io_wgt_data_bits_12_12; // @[TensorGemm.scala 206:53]
  assign dot_0_12_io_b_13 = io_wgt_data_bits_12_13; // @[TensorGemm.scala 206:53]
  assign dot_0_12_io_b_14 = io_wgt_data_bits_12_14; // @[TensorGemm.scala 206:53]
  assign dot_0_12_io_b_15 = io_wgt_data_bits_12_15; // @[TensorGemm.scala 206:53]
  assign dot_0_13_clock = clock;
  assign dot_0_13_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_13_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_13_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_13_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_13_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_13_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_13_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_13_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_13_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_13_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_13_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_13_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_13_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_13_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_13_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_13_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_13_io_b_0 = io_wgt_data_bits_13_0; // @[TensorGemm.scala 206:53]
  assign dot_0_13_io_b_1 = io_wgt_data_bits_13_1; // @[TensorGemm.scala 206:53]
  assign dot_0_13_io_b_2 = io_wgt_data_bits_13_2; // @[TensorGemm.scala 206:53]
  assign dot_0_13_io_b_3 = io_wgt_data_bits_13_3; // @[TensorGemm.scala 206:53]
  assign dot_0_13_io_b_4 = io_wgt_data_bits_13_4; // @[TensorGemm.scala 206:53]
  assign dot_0_13_io_b_5 = io_wgt_data_bits_13_5; // @[TensorGemm.scala 206:53]
  assign dot_0_13_io_b_6 = io_wgt_data_bits_13_6; // @[TensorGemm.scala 206:53]
  assign dot_0_13_io_b_7 = io_wgt_data_bits_13_7; // @[TensorGemm.scala 206:53]
  assign dot_0_13_io_b_8 = io_wgt_data_bits_13_8; // @[TensorGemm.scala 206:53]
  assign dot_0_13_io_b_9 = io_wgt_data_bits_13_9; // @[TensorGemm.scala 206:53]
  assign dot_0_13_io_b_10 = io_wgt_data_bits_13_10; // @[TensorGemm.scala 206:53]
  assign dot_0_13_io_b_11 = io_wgt_data_bits_13_11; // @[TensorGemm.scala 206:53]
  assign dot_0_13_io_b_12 = io_wgt_data_bits_13_12; // @[TensorGemm.scala 206:53]
  assign dot_0_13_io_b_13 = io_wgt_data_bits_13_13; // @[TensorGemm.scala 206:53]
  assign dot_0_13_io_b_14 = io_wgt_data_bits_13_14; // @[TensorGemm.scala 206:53]
  assign dot_0_13_io_b_15 = io_wgt_data_bits_13_15; // @[TensorGemm.scala 206:53]
  assign dot_0_14_clock = clock;
  assign dot_0_14_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_14_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_14_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_14_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_14_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_14_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_14_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_14_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_14_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_14_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_14_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_14_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_14_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_14_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_14_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_14_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_14_io_b_0 = io_wgt_data_bits_14_0; // @[TensorGemm.scala 206:53]
  assign dot_0_14_io_b_1 = io_wgt_data_bits_14_1; // @[TensorGemm.scala 206:53]
  assign dot_0_14_io_b_2 = io_wgt_data_bits_14_2; // @[TensorGemm.scala 206:53]
  assign dot_0_14_io_b_3 = io_wgt_data_bits_14_3; // @[TensorGemm.scala 206:53]
  assign dot_0_14_io_b_4 = io_wgt_data_bits_14_4; // @[TensorGemm.scala 206:53]
  assign dot_0_14_io_b_5 = io_wgt_data_bits_14_5; // @[TensorGemm.scala 206:53]
  assign dot_0_14_io_b_6 = io_wgt_data_bits_14_6; // @[TensorGemm.scala 206:53]
  assign dot_0_14_io_b_7 = io_wgt_data_bits_14_7; // @[TensorGemm.scala 206:53]
  assign dot_0_14_io_b_8 = io_wgt_data_bits_14_8; // @[TensorGemm.scala 206:53]
  assign dot_0_14_io_b_9 = io_wgt_data_bits_14_9; // @[TensorGemm.scala 206:53]
  assign dot_0_14_io_b_10 = io_wgt_data_bits_14_10; // @[TensorGemm.scala 206:53]
  assign dot_0_14_io_b_11 = io_wgt_data_bits_14_11; // @[TensorGemm.scala 206:53]
  assign dot_0_14_io_b_12 = io_wgt_data_bits_14_12; // @[TensorGemm.scala 206:53]
  assign dot_0_14_io_b_13 = io_wgt_data_bits_14_13; // @[TensorGemm.scala 206:53]
  assign dot_0_14_io_b_14 = io_wgt_data_bits_14_14; // @[TensorGemm.scala 206:53]
  assign dot_0_14_io_b_15 = io_wgt_data_bits_14_15; // @[TensorGemm.scala 206:53]
  assign dot_0_15_clock = clock;
  assign dot_0_15_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_15_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_15_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_15_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_15_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_15_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_15_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_15_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_15_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_15_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_15_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_15_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_15_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_15_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_15_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_15_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_15_io_b_0 = io_wgt_data_bits_15_0; // @[TensorGemm.scala 206:53]
  assign dot_0_15_io_b_1 = io_wgt_data_bits_15_1; // @[TensorGemm.scala 206:53]
  assign dot_0_15_io_b_2 = io_wgt_data_bits_15_2; // @[TensorGemm.scala 206:53]
  assign dot_0_15_io_b_3 = io_wgt_data_bits_15_3; // @[TensorGemm.scala 206:53]
  assign dot_0_15_io_b_4 = io_wgt_data_bits_15_4; // @[TensorGemm.scala 206:53]
  assign dot_0_15_io_b_5 = io_wgt_data_bits_15_5; // @[TensorGemm.scala 206:53]
  assign dot_0_15_io_b_6 = io_wgt_data_bits_15_6; // @[TensorGemm.scala 206:53]
  assign dot_0_15_io_b_7 = io_wgt_data_bits_15_7; // @[TensorGemm.scala 206:53]
  assign dot_0_15_io_b_8 = io_wgt_data_bits_15_8; // @[TensorGemm.scala 206:53]
  assign dot_0_15_io_b_9 = io_wgt_data_bits_15_9; // @[TensorGemm.scala 206:53]
  assign dot_0_15_io_b_10 = io_wgt_data_bits_15_10; // @[TensorGemm.scala 206:53]
  assign dot_0_15_io_b_11 = io_wgt_data_bits_15_11; // @[TensorGemm.scala 206:53]
  assign dot_0_15_io_b_12 = io_wgt_data_bits_15_12; // @[TensorGemm.scala 206:53]
  assign dot_0_15_io_b_13 = io_wgt_data_bits_15_13; // @[TensorGemm.scala 206:53]
  assign dot_0_15_io_b_14 = io_wgt_data_bits_15_14; // @[TensorGemm.scala 206:53]
  assign dot_0_15_io_b_15 = io_wgt_data_bits_15_15; // @[TensorGemm.scala 206:53]
  assign dot_0_16_clock = clock;
  assign dot_0_16_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_16_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_16_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_16_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_16_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_16_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_16_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_16_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_16_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_16_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_16_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_16_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_16_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_16_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_16_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_16_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_16_io_b_0 = io_wgt_data_bits_16_0; // @[TensorGemm.scala 206:53]
  assign dot_0_16_io_b_1 = io_wgt_data_bits_16_1; // @[TensorGemm.scala 206:53]
  assign dot_0_16_io_b_2 = io_wgt_data_bits_16_2; // @[TensorGemm.scala 206:53]
  assign dot_0_16_io_b_3 = io_wgt_data_bits_16_3; // @[TensorGemm.scala 206:53]
  assign dot_0_16_io_b_4 = io_wgt_data_bits_16_4; // @[TensorGemm.scala 206:53]
  assign dot_0_16_io_b_5 = io_wgt_data_bits_16_5; // @[TensorGemm.scala 206:53]
  assign dot_0_16_io_b_6 = io_wgt_data_bits_16_6; // @[TensorGemm.scala 206:53]
  assign dot_0_16_io_b_7 = io_wgt_data_bits_16_7; // @[TensorGemm.scala 206:53]
  assign dot_0_16_io_b_8 = io_wgt_data_bits_16_8; // @[TensorGemm.scala 206:53]
  assign dot_0_16_io_b_9 = io_wgt_data_bits_16_9; // @[TensorGemm.scala 206:53]
  assign dot_0_16_io_b_10 = io_wgt_data_bits_16_10; // @[TensorGemm.scala 206:53]
  assign dot_0_16_io_b_11 = io_wgt_data_bits_16_11; // @[TensorGemm.scala 206:53]
  assign dot_0_16_io_b_12 = io_wgt_data_bits_16_12; // @[TensorGemm.scala 206:53]
  assign dot_0_16_io_b_13 = io_wgt_data_bits_16_13; // @[TensorGemm.scala 206:53]
  assign dot_0_16_io_b_14 = io_wgt_data_bits_16_14; // @[TensorGemm.scala 206:53]
  assign dot_0_16_io_b_15 = io_wgt_data_bits_16_15; // @[TensorGemm.scala 206:53]
  assign dot_0_17_clock = clock;
  assign dot_0_17_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_17_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_17_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_17_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_17_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_17_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_17_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_17_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_17_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_17_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_17_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_17_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_17_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_17_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_17_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_17_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_17_io_b_0 = io_wgt_data_bits_17_0; // @[TensorGemm.scala 206:53]
  assign dot_0_17_io_b_1 = io_wgt_data_bits_17_1; // @[TensorGemm.scala 206:53]
  assign dot_0_17_io_b_2 = io_wgt_data_bits_17_2; // @[TensorGemm.scala 206:53]
  assign dot_0_17_io_b_3 = io_wgt_data_bits_17_3; // @[TensorGemm.scala 206:53]
  assign dot_0_17_io_b_4 = io_wgt_data_bits_17_4; // @[TensorGemm.scala 206:53]
  assign dot_0_17_io_b_5 = io_wgt_data_bits_17_5; // @[TensorGemm.scala 206:53]
  assign dot_0_17_io_b_6 = io_wgt_data_bits_17_6; // @[TensorGemm.scala 206:53]
  assign dot_0_17_io_b_7 = io_wgt_data_bits_17_7; // @[TensorGemm.scala 206:53]
  assign dot_0_17_io_b_8 = io_wgt_data_bits_17_8; // @[TensorGemm.scala 206:53]
  assign dot_0_17_io_b_9 = io_wgt_data_bits_17_9; // @[TensorGemm.scala 206:53]
  assign dot_0_17_io_b_10 = io_wgt_data_bits_17_10; // @[TensorGemm.scala 206:53]
  assign dot_0_17_io_b_11 = io_wgt_data_bits_17_11; // @[TensorGemm.scala 206:53]
  assign dot_0_17_io_b_12 = io_wgt_data_bits_17_12; // @[TensorGemm.scala 206:53]
  assign dot_0_17_io_b_13 = io_wgt_data_bits_17_13; // @[TensorGemm.scala 206:53]
  assign dot_0_17_io_b_14 = io_wgt_data_bits_17_14; // @[TensorGemm.scala 206:53]
  assign dot_0_17_io_b_15 = io_wgt_data_bits_17_15; // @[TensorGemm.scala 206:53]
  assign dot_0_18_clock = clock;
  assign dot_0_18_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_18_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_18_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_18_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_18_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_18_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_18_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_18_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_18_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_18_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_18_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_18_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_18_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_18_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_18_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_18_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_18_io_b_0 = io_wgt_data_bits_18_0; // @[TensorGemm.scala 206:53]
  assign dot_0_18_io_b_1 = io_wgt_data_bits_18_1; // @[TensorGemm.scala 206:53]
  assign dot_0_18_io_b_2 = io_wgt_data_bits_18_2; // @[TensorGemm.scala 206:53]
  assign dot_0_18_io_b_3 = io_wgt_data_bits_18_3; // @[TensorGemm.scala 206:53]
  assign dot_0_18_io_b_4 = io_wgt_data_bits_18_4; // @[TensorGemm.scala 206:53]
  assign dot_0_18_io_b_5 = io_wgt_data_bits_18_5; // @[TensorGemm.scala 206:53]
  assign dot_0_18_io_b_6 = io_wgt_data_bits_18_6; // @[TensorGemm.scala 206:53]
  assign dot_0_18_io_b_7 = io_wgt_data_bits_18_7; // @[TensorGemm.scala 206:53]
  assign dot_0_18_io_b_8 = io_wgt_data_bits_18_8; // @[TensorGemm.scala 206:53]
  assign dot_0_18_io_b_9 = io_wgt_data_bits_18_9; // @[TensorGemm.scala 206:53]
  assign dot_0_18_io_b_10 = io_wgt_data_bits_18_10; // @[TensorGemm.scala 206:53]
  assign dot_0_18_io_b_11 = io_wgt_data_bits_18_11; // @[TensorGemm.scala 206:53]
  assign dot_0_18_io_b_12 = io_wgt_data_bits_18_12; // @[TensorGemm.scala 206:53]
  assign dot_0_18_io_b_13 = io_wgt_data_bits_18_13; // @[TensorGemm.scala 206:53]
  assign dot_0_18_io_b_14 = io_wgt_data_bits_18_14; // @[TensorGemm.scala 206:53]
  assign dot_0_18_io_b_15 = io_wgt_data_bits_18_15; // @[TensorGemm.scala 206:53]
  assign dot_0_19_clock = clock;
  assign dot_0_19_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_19_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_19_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_19_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_19_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_19_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_19_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_19_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_19_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_19_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_19_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_19_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_19_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_19_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_19_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_19_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_19_io_b_0 = io_wgt_data_bits_19_0; // @[TensorGemm.scala 206:53]
  assign dot_0_19_io_b_1 = io_wgt_data_bits_19_1; // @[TensorGemm.scala 206:53]
  assign dot_0_19_io_b_2 = io_wgt_data_bits_19_2; // @[TensorGemm.scala 206:53]
  assign dot_0_19_io_b_3 = io_wgt_data_bits_19_3; // @[TensorGemm.scala 206:53]
  assign dot_0_19_io_b_4 = io_wgt_data_bits_19_4; // @[TensorGemm.scala 206:53]
  assign dot_0_19_io_b_5 = io_wgt_data_bits_19_5; // @[TensorGemm.scala 206:53]
  assign dot_0_19_io_b_6 = io_wgt_data_bits_19_6; // @[TensorGemm.scala 206:53]
  assign dot_0_19_io_b_7 = io_wgt_data_bits_19_7; // @[TensorGemm.scala 206:53]
  assign dot_0_19_io_b_8 = io_wgt_data_bits_19_8; // @[TensorGemm.scala 206:53]
  assign dot_0_19_io_b_9 = io_wgt_data_bits_19_9; // @[TensorGemm.scala 206:53]
  assign dot_0_19_io_b_10 = io_wgt_data_bits_19_10; // @[TensorGemm.scala 206:53]
  assign dot_0_19_io_b_11 = io_wgt_data_bits_19_11; // @[TensorGemm.scala 206:53]
  assign dot_0_19_io_b_12 = io_wgt_data_bits_19_12; // @[TensorGemm.scala 206:53]
  assign dot_0_19_io_b_13 = io_wgt_data_bits_19_13; // @[TensorGemm.scala 206:53]
  assign dot_0_19_io_b_14 = io_wgt_data_bits_19_14; // @[TensorGemm.scala 206:53]
  assign dot_0_19_io_b_15 = io_wgt_data_bits_19_15; // @[TensorGemm.scala 206:53]
  assign dot_0_20_clock = clock;
  assign dot_0_20_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_20_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_20_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_20_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_20_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_20_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_20_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_20_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_20_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_20_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_20_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_20_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_20_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_20_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_20_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_20_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_20_io_b_0 = io_wgt_data_bits_20_0; // @[TensorGemm.scala 206:53]
  assign dot_0_20_io_b_1 = io_wgt_data_bits_20_1; // @[TensorGemm.scala 206:53]
  assign dot_0_20_io_b_2 = io_wgt_data_bits_20_2; // @[TensorGemm.scala 206:53]
  assign dot_0_20_io_b_3 = io_wgt_data_bits_20_3; // @[TensorGemm.scala 206:53]
  assign dot_0_20_io_b_4 = io_wgt_data_bits_20_4; // @[TensorGemm.scala 206:53]
  assign dot_0_20_io_b_5 = io_wgt_data_bits_20_5; // @[TensorGemm.scala 206:53]
  assign dot_0_20_io_b_6 = io_wgt_data_bits_20_6; // @[TensorGemm.scala 206:53]
  assign dot_0_20_io_b_7 = io_wgt_data_bits_20_7; // @[TensorGemm.scala 206:53]
  assign dot_0_20_io_b_8 = io_wgt_data_bits_20_8; // @[TensorGemm.scala 206:53]
  assign dot_0_20_io_b_9 = io_wgt_data_bits_20_9; // @[TensorGemm.scala 206:53]
  assign dot_0_20_io_b_10 = io_wgt_data_bits_20_10; // @[TensorGemm.scala 206:53]
  assign dot_0_20_io_b_11 = io_wgt_data_bits_20_11; // @[TensorGemm.scala 206:53]
  assign dot_0_20_io_b_12 = io_wgt_data_bits_20_12; // @[TensorGemm.scala 206:53]
  assign dot_0_20_io_b_13 = io_wgt_data_bits_20_13; // @[TensorGemm.scala 206:53]
  assign dot_0_20_io_b_14 = io_wgt_data_bits_20_14; // @[TensorGemm.scala 206:53]
  assign dot_0_20_io_b_15 = io_wgt_data_bits_20_15; // @[TensorGemm.scala 206:53]
  assign dot_0_21_clock = clock;
  assign dot_0_21_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_21_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_21_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_21_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_21_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_21_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_21_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_21_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_21_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_21_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_21_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_21_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_21_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_21_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_21_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_21_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_21_io_b_0 = io_wgt_data_bits_21_0; // @[TensorGemm.scala 206:53]
  assign dot_0_21_io_b_1 = io_wgt_data_bits_21_1; // @[TensorGemm.scala 206:53]
  assign dot_0_21_io_b_2 = io_wgt_data_bits_21_2; // @[TensorGemm.scala 206:53]
  assign dot_0_21_io_b_3 = io_wgt_data_bits_21_3; // @[TensorGemm.scala 206:53]
  assign dot_0_21_io_b_4 = io_wgt_data_bits_21_4; // @[TensorGemm.scala 206:53]
  assign dot_0_21_io_b_5 = io_wgt_data_bits_21_5; // @[TensorGemm.scala 206:53]
  assign dot_0_21_io_b_6 = io_wgt_data_bits_21_6; // @[TensorGemm.scala 206:53]
  assign dot_0_21_io_b_7 = io_wgt_data_bits_21_7; // @[TensorGemm.scala 206:53]
  assign dot_0_21_io_b_8 = io_wgt_data_bits_21_8; // @[TensorGemm.scala 206:53]
  assign dot_0_21_io_b_9 = io_wgt_data_bits_21_9; // @[TensorGemm.scala 206:53]
  assign dot_0_21_io_b_10 = io_wgt_data_bits_21_10; // @[TensorGemm.scala 206:53]
  assign dot_0_21_io_b_11 = io_wgt_data_bits_21_11; // @[TensorGemm.scala 206:53]
  assign dot_0_21_io_b_12 = io_wgt_data_bits_21_12; // @[TensorGemm.scala 206:53]
  assign dot_0_21_io_b_13 = io_wgt_data_bits_21_13; // @[TensorGemm.scala 206:53]
  assign dot_0_21_io_b_14 = io_wgt_data_bits_21_14; // @[TensorGemm.scala 206:53]
  assign dot_0_21_io_b_15 = io_wgt_data_bits_21_15; // @[TensorGemm.scala 206:53]
  assign dot_0_22_clock = clock;
  assign dot_0_22_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_22_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_22_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_22_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_22_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_22_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_22_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_22_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_22_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_22_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_22_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_22_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_22_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_22_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_22_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_22_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_22_io_b_0 = io_wgt_data_bits_22_0; // @[TensorGemm.scala 206:53]
  assign dot_0_22_io_b_1 = io_wgt_data_bits_22_1; // @[TensorGemm.scala 206:53]
  assign dot_0_22_io_b_2 = io_wgt_data_bits_22_2; // @[TensorGemm.scala 206:53]
  assign dot_0_22_io_b_3 = io_wgt_data_bits_22_3; // @[TensorGemm.scala 206:53]
  assign dot_0_22_io_b_4 = io_wgt_data_bits_22_4; // @[TensorGemm.scala 206:53]
  assign dot_0_22_io_b_5 = io_wgt_data_bits_22_5; // @[TensorGemm.scala 206:53]
  assign dot_0_22_io_b_6 = io_wgt_data_bits_22_6; // @[TensorGemm.scala 206:53]
  assign dot_0_22_io_b_7 = io_wgt_data_bits_22_7; // @[TensorGemm.scala 206:53]
  assign dot_0_22_io_b_8 = io_wgt_data_bits_22_8; // @[TensorGemm.scala 206:53]
  assign dot_0_22_io_b_9 = io_wgt_data_bits_22_9; // @[TensorGemm.scala 206:53]
  assign dot_0_22_io_b_10 = io_wgt_data_bits_22_10; // @[TensorGemm.scala 206:53]
  assign dot_0_22_io_b_11 = io_wgt_data_bits_22_11; // @[TensorGemm.scala 206:53]
  assign dot_0_22_io_b_12 = io_wgt_data_bits_22_12; // @[TensorGemm.scala 206:53]
  assign dot_0_22_io_b_13 = io_wgt_data_bits_22_13; // @[TensorGemm.scala 206:53]
  assign dot_0_22_io_b_14 = io_wgt_data_bits_22_14; // @[TensorGemm.scala 206:53]
  assign dot_0_22_io_b_15 = io_wgt_data_bits_22_15; // @[TensorGemm.scala 206:53]
  assign dot_0_23_clock = clock;
  assign dot_0_23_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_23_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_23_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_23_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_23_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_23_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_23_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_23_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_23_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_23_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_23_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_23_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_23_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_23_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_23_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_23_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_23_io_b_0 = io_wgt_data_bits_23_0; // @[TensorGemm.scala 206:53]
  assign dot_0_23_io_b_1 = io_wgt_data_bits_23_1; // @[TensorGemm.scala 206:53]
  assign dot_0_23_io_b_2 = io_wgt_data_bits_23_2; // @[TensorGemm.scala 206:53]
  assign dot_0_23_io_b_3 = io_wgt_data_bits_23_3; // @[TensorGemm.scala 206:53]
  assign dot_0_23_io_b_4 = io_wgt_data_bits_23_4; // @[TensorGemm.scala 206:53]
  assign dot_0_23_io_b_5 = io_wgt_data_bits_23_5; // @[TensorGemm.scala 206:53]
  assign dot_0_23_io_b_6 = io_wgt_data_bits_23_6; // @[TensorGemm.scala 206:53]
  assign dot_0_23_io_b_7 = io_wgt_data_bits_23_7; // @[TensorGemm.scala 206:53]
  assign dot_0_23_io_b_8 = io_wgt_data_bits_23_8; // @[TensorGemm.scala 206:53]
  assign dot_0_23_io_b_9 = io_wgt_data_bits_23_9; // @[TensorGemm.scala 206:53]
  assign dot_0_23_io_b_10 = io_wgt_data_bits_23_10; // @[TensorGemm.scala 206:53]
  assign dot_0_23_io_b_11 = io_wgt_data_bits_23_11; // @[TensorGemm.scala 206:53]
  assign dot_0_23_io_b_12 = io_wgt_data_bits_23_12; // @[TensorGemm.scala 206:53]
  assign dot_0_23_io_b_13 = io_wgt_data_bits_23_13; // @[TensorGemm.scala 206:53]
  assign dot_0_23_io_b_14 = io_wgt_data_bits_23_14; // @[TensorGemm.scala 206:53]
  assign dot_0_23_io_b_15 = io_wgt_data_bits_23_15; // @[TensorGemm.scala 206:53]
  assign dot_0_24_clock = clock;
  assign dot_0_24_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_24_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_24_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_24_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_24_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_24_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_24_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_24_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_24_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_24_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_24_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_24_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_24_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_24_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_24_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_24_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_24_io_b_0 = io_wgt_data_bits_24_0; // @[TensorGemm.scala 206:53]
  assign dot_0_24_io_b_1 = io_wgt_data_bits_24_1; // @[TensorGemm.scala 206:53]
  assign dot_0_24_io_b_2 = io_wgt_data_bits_24_2; // @[TensorGemm.scala 206:53]
  assign dot_0_24_io_b_3 = io_wgt_data_bits_24_3; // @[TensorGemm.scala 206:53]
  assign dot_0_24_io_b_4 = io_wgt_data_bits_24_4; // @[TensorGemm.scala 206:53]
  assign dot_0_24_io_b_5 = io_wgt_data_bits_24_5; // @[TensorGemm.scala 206:53]
  assign dot_0_24_io_b_6 = io_wgt_data_bits_24_6; // @[TensorGemm.scala 206:53]
  assign dot_0_24_io_b_7 = io_wgt_data_bits_24_7; // @[TensorGemm.scala 206:53]
  assign dot_0_24_io_b_8 = io_wgt_data_bits_24_8; // @[TensorGemm.scala 206:53]
  assign dot_0_24_io_b_9 = io_wgt_data_bits_24_9; // @[TensorGemm.scala 206:53]
  assign dot_0_24_io_b_10 = io_wgt_data_bits_24_10; // @[TensorGemm.scala 206:53]
  assign dot_0_24_io_b_11 = io_wgt_data_bits_24_11; // @[TensorGemm.scala 206:53]
  assign dot_0_24_io_b_12 = io_wgt_data_bits_24_12; // @[TensorGemm.scala 206:53]
  assign dot_0_24_io_b_13 = io_wgt_data_bits_24_13; // @[TensorGemm.scala 206:53]
  assign dot_0_24_io_b_14 = io_wgt_data_bits_24_14; // @[TensorGemm.scala 206:53]
  assign dot_0_24_io_b_15 = io_wgt_data_bits_24_15; // @[TensorGemm.scala 206:53]
  assign dot_0_25_clock = clock;
  assign dot_0_25_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_25_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_25_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_25_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_25_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_25_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_25_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_25_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_25_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_25_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_25_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_25_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_25_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_25_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_25_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_25_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_25_io_b_0 = io_wgt_data_bits_25_0; // @[TensorGemm.scala 206:53]
  assign dot_0_25_io_b_1 = io_wgt_data_bits_25_1; // @[TensorGemm.scala 206:53]
  assign dot_0_25_io_b_2 = io_wgt_data_bits_25_2; // @[TensorGemm.scala 206:53]
  assign dot_0_25_io_b_3 = io_wgt_data_bits_25_3; // @[TensorGemm.scala 206:53]
  assign dot_0_25_io_b_4 = io_wgt_data_bits_25_4; // @[TensorGemm.scala 206:53]
  assign dot_0_25_io_b_5 = io_wgt_data_bits_25_5; // @[TensorGemm.scala 206:53]
  assign dot_0_25_io_b_6 = io_wgt_data_bits_25_6; // @[TensorGemm.scala 206:53]
  assign dot_0_25_io_b_7 = io_wgt_data_bits_25_7; // @[TensorGemm.scala 206:53]
  assign dot_0_25_io_b_8 = io_wgt_data_bits_25_8; // @[TensorGemm.scala 206:53]
  assign dot_0_25_io_b_9 = io_wgt_data_bits_25_9; // @[TensorGemm.scala 206:53]
  assign dot_0_25_io_b_10 = io_wgt_data_bits_25_10; // @[TensorGemm.scala 206:53]
  assign dot_0_25_io_b_11 = io_wgt_data_bits_25_11; // @[TensorGemm.scala 206:53]
  assign dot_0_25_io_b_12 = io_wgt_data_bits_25_12; // @[TensorGemm.scala 206:53]
  assign dot_0_25_io_b_13 = io_wgt_data_bits_25_13; // @[TensorGemm.scala 206:53]
  assign dot_0_25_io_b_14 = io_wgt_data_bits_25_14; // @[TensorGemm.scala 206:53]
  assign dot_0_25_io_b_15 = io_wgt_data_bits_25_15; // @[TensorGemm.scala 206:53]
  assign dot_0_26_clock = clock;
  assign dot_0_26_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_26_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_26_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_26_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_26_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_26_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_26_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_26_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_26_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_26_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_26_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_26_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_26_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_26_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_26_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_26_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_26_io_b_0 = io_wgt_data_bits_26_0; // @[TensorGemm.scala 206:53]
  assign dot_0_26_io_b_1 = io_wgt_data_bits_26_1; // @[TensorGemm.scala 206:53]
  assign dot_0_26_io_b_2 = io_wgt_data_bits_26_2; // @[TensorGemm.scala 206:53]
  assign dot_0_26_io_b_3 = io_wgt_data_bits_26_3; // @[TensorGemm.scala 206:53]
  assign dot_0_26_io_b_4 = io_wgt_data_bits_26_4; // @[TensorGemm.scala 206:53]
  assign dot_0_26_io_b_5 = io_wgt_data_bits_26_5; // @[TensorGemm.scala 206:53]
  assign dot_0_26_io_b_6 = io_wgt_data_bits_26_6; // @[TensorGemm.scala 206:53]
  assign dot_0_26_io_b_7 = io_wgt_data_bits_26_7; // @[TensorGemm.scala 206:53]
  assign dot_0_26_io_b_8 = io_wgt_data_bits_26_8; // @[TensorGemm.scala 206:53]
  assign dot_0_26_io_b_9 = io_wgt_data_bits_26_9; // @[TensorGemm.scala 206:53]
  assign dot_0_26_io_b_10 = io_wgt_data_bits_26_10; // @[TensorGemm.scala 206:53]
  assign dot_0_26_io_b_11 = io_wgt_data_bits_26_11; // @[TensorGemm.scala 206:53]
  assign dot_0_26_io_b_12 = io_wgt_data_bits_26_12; // @[TensorGemm.scala 206:53]
  assign dot_0_26_io_b_13 = io_wgt_data_bits_26_13; // @[TensorGemm.scala 206:53]
  assign dot_0_26_io_b_14 = io_wgt_data_bits_26_14; // @[TensorGemm.scala 206:53]
  assign dot_0_26_io_b_15 = io_wgt_data_bits_26_15; // @[TensorGemm.scala 206:53]
  assign dot_0_27_clock = clock;
  assign dot_0_27_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_27_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_27_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_27_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_27_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_27_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_27_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_27_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_27_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_27_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_27_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_27_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_27_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_27_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_27_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_27_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_27_io_b_0 = io_wgt_data_bits_27_0; // @[TensorGemm.scala 206:53]
  assign dot_0_27_io_b_1 = io_wgt_data_bits_27_1; // @[TensorGemm.scala 206:53]
  assign dot_0_27_io_b_2 = io_wgt_data_bits_27_2; // @[TensorGemm.scala 206:53]
  assign dot_0_27_io_b_3 = io_wgt_data_bits_27_3; // @[TensorGemm.scala 206:53]
  assign dot_0_27_io_b_4 = io_wgt_data_bits_27_4; // @[TensorGemm.scala 206:53]
  assign dot_0_27_io_b_5 = io_wgt_data_bits_27_5; // @[TensorGemm.scala 206:53]
  assign dot_0_27_io_b_6 = io_wgt_data_bits_27_6; // @[TensorGemm.scala 206:53]
  assign dot_0_27_io_b_7 = io_wgt_data_bits_27_7; // @[TensorGemm.scala 206:53]
  assign dot_0_27_io_b_8 = io_wgt_data_bits_27_8; // @[TensorGemm.scala 206:53]
  assign dot_0_27_io_b_9 = io_wgt_data_bits_27_9; // @[TensorGemm.scala 206:53]
  assign dot_0_27_io_b_10 = io_wgt_data_bits_27_10; // @[TensorGemm.scala 206:53]
  assign dot_0_27_io_b_11 = io_wgt_data_bits_27_11; // @[TensorGemm.scala 206:53]
  assign dot_0_27_io_b_12 = io_wgt_data_bits_27_12; // @[TensorGemm.scala 206:53]
  assign dot_0_27_io_b_13 = io_wgt_data_bits_27_13; // @[TensorGemm.scala 206:53]
  assign dot_0_27_io_b_14 = io_wgt_data_bits_27_14; // @[TensorGemm.scala 206:53]
  assign dot_0_27_io_b_15 = io_wgt_data_bits_27_15; // @[TensorGemm.scala 206:53]
  assign dot_0_28_clock = clock;
  assign dot_0_28_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_28_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_28_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_28_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_28_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_28_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_28_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_28_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_28_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_28_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_28_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_28_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_28_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_28_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_28_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_28_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_28_io_b_0 = io_wgt_data_bits_28_0; // @[TensorGemm.scala 206:53]
  assign dot_0_28_io_b_1 = io_wgt_data_bits_28_1; // @[TensorGemm.scala 206:53]
  assign dot_0_28_io_b_2 = io_wgt_data_bits_28_2; // @[TensorGemm.scala 206:53]
  assign dot_0_28_io_b_3 = io_wgt_data_bits_28_3; // @[TensorGemm.scala 206:53]
  assign dot_0_28_io_b_4 = io_wgt_data_bits_28_4; // @[TensorGemm.scala 206:53]
  assign dot_0_28_io_b_5 = io_wgt_data_bits_28_5; // @[TensorGemm.scala 206:53]
  assign dot_0_28_io_b_6 = io_wgt_data_bits_28_6; // @[TensorGemm.scala 206:53]
  assign dot_0_28_io_b_7 = io_wgt_data_bits_28_7; // @[TensorGemm.scala 206:53]
  assign dot_0_28_io_b_8 = io_wgt_data_bits_28_8; // @[TensorGemm.scala 206:53]
  assign dot_0_28_io_b_9 = io_wgt_data_bits_28_9; // @[TensorGemm.scala 206:53]
  assign dot_0_28_io_b_10 = io_wgt_data_bits_28_10; // @[TensorGemm.scala 206:53]
  assign dot_0_28_io_b_11 = io_wgt_data_bits_28_11; // @[TensorGemm.scala 206:53]
  assign dot_0_28_io_b_12 = io_wgt_data_bits_28_12; // @[TensorGemm.scala 206:53]
  assign dot_0_28_io_b_13 = io_wgt_data_bits_28_13; // @[TensorGemm.scala 206:53]
  assign dot_0_28_io_b_14 = io_wgt_data_bits_28_14; // @[TensorGemm.scala 206:53]
  assign dot_0_28_io_b_15 = io_wgt_data_bits_28_15; // @[TensorGemm.scala 206:53]
  assign dot_0_29_clock = clock;
  assign dot_0_29_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_29_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_29_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_29_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_29_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_29_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_29_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_29_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_29_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_29_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_29_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_29_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_29_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_29_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_29_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_29_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_29_io_b_0 = io_wgt_data_bits_29_0; // @[TensorGemm.scala 206:53]
  assign dot_0_29_io_b_1 = io_wgt_data_bits_29_1; // @[TensorGemm.scala 206:53]
  assign dot_0_29_io_b_2 = io_wgt_data_bits_29_2; // @[TensorGemm.scala 206:53]
  assign dot_0_29_io_b_3 = io_wgt_data_bits_29_3; // @[TensorGemm.scala 206:53]
  assign dot_0_29_io_b_4 = io_wgt_data_bits_29_4; // @[TensorGemm.scala 206:53]
  assign dot_0_29_io_b_5 = io_wgt_data_bits_29_5; // @[TensorGemm.scala 206:53]
  assign dot_0_29_io_b_6 = io_wgt_data_bits_29_6; // @[TensorGemm.scala 206:53]
  assign dot_0_29_io_b_7 = io_wgt_data_bits_29_7; // @[TensorGemm.scala 206:53]
  assign dot_0_29_io_b_8 = io_wgt_data_bits_29_8; // @[TensorGemm.scala 206:53]
  assign dot_0_29_io_b_9 = io_wgt_data_bits_29_9; // @[TensorGemm.scala 206:53]
  assign dot_0_29_io_b_10 = io_wgt_data_bits_29_10; // @[TensorGemm.scala 206:53]
  assign dot_0_29_io_b_11 = io_wgt_data_bits_29_11; // @[TensorGemm.scala 206:53]
  assign dot_0_29_io_b_12 = io_wgt_data_bits_29_12; // @[TensorGemm.scala 206:53]
  assign dot_0_29_io_b_13 = io_wgt_data_bits_29_13; // @[TensorGemm.scala 206:53]
  assign dot_0_29_io_b_14 = io_wgt_data_bits_29_14; // @[TensorGemm.scala 206:53]
  assign dot_0_29_io_b_15 = io_wgt_data_bits_29_15; // @[TensorGemm.scala 206:53]
  assign dot_0_30_clock = clock;
  assign dot_0_30_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_30_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_30_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_30_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_30_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_30_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_30_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_30_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_30_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_30_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_30_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_30_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_30_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_30_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_30_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_30_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_30_io_b_0 = io_wgt_data_bits_30_0; // @[TensorGemm.scala 206:53]
  assign dot_0_30_io_b_1 = io_wgt_data_bits_30_1; // @[TensorGemm.scala 206:53]
  assign dot_0_30_io_b_2 = io_wgt_data_bits_30_2; // @[TensorGemm.scala 206:53]
  assign dot_0_30_io_b_3 = io_wgt_data_bits_30_3; // @[TensorGemm.scala 206:53]
  assign dot_0_30_io_b_4 = io_wgt_data_bits_30_4; // @[TensorGemm.scala 206:53]
  assign dot_0_30_io_b_5 = io_wgt_data_bits_30_5; // @[TensorGemm.scala 206:53]
  assign dot_0_30_io_b_6 = io_wgt_data_bits_30_6; // @[TensorGemm.scala 206:53]
  assign dot_0_30_io_b_7 = io_wgt_data_bits_30_7; // @[TensorGemm.scala 206:53]
  assign dot_0_30_io_b_8 = io_wgt_data_bits_30_8; // @[TensorGemm.scala 206:53]
  assign dot_0_30_io_b_9 = io_wgt_data_bits_30_9; // @[TensorGemm.scala 206:53]
  assign dot_0_30_io_b_10 = io_wgt_data_bits_30_10; // @[TensorGemm.scala 206:53]
  assign dot_0_30_io_b_11 = io_wgt_data_bits_30_11; // @[TensorGemm.scala 206:53]
  assign dot_0_30_io_b_12 = io_wgt_data_bits_30_12; // @[TensorGemm.scala 206:53]
  assign dot_0_30_io_b_13 = io_wgt_data_bits_30_13; // @[TensorGemm.scala 206:53]
  assign dot_0_30_io_b_14 = io_wgt_data_bits_30_14; // @[TensorGemm.scala 206:53]
  assign dot_0_30_io_b_15 = io_wgt_data_bits_30_15; // @[TensorGemm.scala 206:53]
  assign dot_0_31_clock = clock;
  assign dot_0_31_io_a_0 = io_inp_data_bits_0_0; // @[TensorGemm.scala 205:53]
  assign dot_0_31_io_a_1 = io_inp_data_bits_0_1; // @[TensorGemm.scala 205:53]
  assign dot_0_31_io_a_2 = io_inp_data_bits_0_2; // @[TensorGemm.scala 205:53]
  assign dot_0_31_io_a_3 = io_inp_data_bits_0_3; // @[TensorGemm.scala 205:53]
  assign dot_0_31_io_a_4 = io_inp_data_bits_0_4; // @[TensorGemm.scala 205:53]
  assign dot_0_31_io_a_5 = io_inp_data_bits_0_5; // @[TensorGemm.scala 205:53]
  assign dot_0_31_io_a_6 = io_inp_data_bits_0_6; // @[TensorGemm.scala 205:53]
  assign dot_0_31_io_a_7 = io_inp_data_bits_0_7; // @[TensorGemm.scala 205:53]
  assign dot_0_31_io_a_8 = io_inp_data_bits_0_8; // @[TensorGemm.scala 205:53]
  assign dot_0_31_io_a_9 = io_inp_data_bits_0_9; // @[TensorGemm.scala 205:53]
  assign dot_0_31_io_a_10 = io_inp_data_bits_0_10; // @[TensorGemm.scala 205:53]
  assign dot_0_31_io_a_11 = io_inp_data_bits_0_11; // @[TensorGemm.scala 205:53]
  assign dot_0_31_io_a_12 = io_inp_data_bits_0_12; // @[TensorGemm.scala 205:53]
  assign dot_0_31_io_a_13 = io_inp_data_bits_0_13; // @[TensorGemm.scala 205:53]
  assign dot_0_31_io_a_14 = io_inp_data_bits_0_14; // @[TensorGemm.scala 205:53]
  assign dot_0_31_io_a_15 = io_inp_data_bits_0_15; // @[TensorGemm.scala 205:53]
  assign dot_0_31_io_b_0 = io_wgt_data_bits_31_0; // @[TensorGemm.scala 206:53]
  assign dot_0_31_io_b_1 = io_wgt_data_bits_31_1; // @[TensorGemm.scala 206:53]
  assign dot_0_31_io_b_2 = io_wgt_data_bits_31_2; // @[TensorGemm.scala 206:53]
  assign dot_0_31_io_b_3 = io_wgt_data_bits_31_3; // @[TensorGemm.scala 206:53]
  assign dot_0_31_io_b_4 = io_wgt_data_bits_31_4; // @[TensorGemm.scala 206:53]
  assign dot_0_31_io_b_5 = io_wgt_data_bits_31_5; // @[TensorGemm.scala 206:53]
  assign dot_0_31_io_b_6 = io_wgt_data_bits_31_6; // @[TensorGemm.scala 206:53]
  assign dot_0_31_io_b_7 = io_wgt_data_bits_31_7; // @[TensorGemm.scala 206:53]
  assign dot_0_31_io_b_8 = io_wgt_data_bits_31_8; // @[TensorGemm.scala 206:53]
  assign dot_0_31_io_b_9 = io_wgt_data_bits_31_9; // @[TensorGemm.scala 206:53]
  assign dot_0_31_io_b_10 = io_wgt_data_bits_31_10; // @[TensorGemm.scala 206:53]
  assign dot_0_31_io_b_11 = io_wgt_data_bits_31_11; // @[TensorGemm.scala 206:53]
  assign dot_0_31_io_b_12 = io_wgt_data_bits_31_12; // @[TensorGemm.scala 206:53]
  assign dot_0_31_io_b_13 = io_wgt_data_bits_31_13; // @[TensorGemm.scala 206:53]
  assign dot_0_31_io_b_14 = io_wgt_data_bits_31_14; // @[TensorGemm.scala 206:53]
  assign dot_0_31_io_b_15 = io_wgt_data_bits_31_15; // @[TensorGemm.scala 206:53]
  always @(posedge clock) begin
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_0 <= 32'sh0;
    end else begin
      last_acc_write_0_0 <= add_0_0;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_1 <= 32'sh0;
    end else begin
      last_acc_write_0_1 <= add_0_1;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_2 <= 32'sh0;
    end else begin
      last_acc_write_0_2 <= add_0_2;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_3 <= 32'sh0;
    end else begin
      last_acc_write_0_3 <= add_0_3;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_4 <= 32'sh0;
    end else begin
      last_acc_write_0_4 <= add_0_4;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_5 <= 32'sh0;
    end else begin
      last_acc_write_0_5 <= add_0_5;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_6 <= 32'sh0;
    end else begin
      last_acc_write_0_6 <= add_0_6;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_7 <= 32'sh0;
    end else begin
      last_acc_write_0_7 <= add_0_7;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_8 <= 32'sh0;
    end else begin
      last_acc_write_0_8 <= add_0_8;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_9 <= 32'sh0;
    end else begin
      last_acc_write_0_9 <= add_0_9;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_10 <= 32'sh0;
    end else begin
      last_acc_write_0_10 <= add_0_10;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_11 <= 32'sh0;
    end else begin
      last_acc_write_0_11 <= add_0_11;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_12 <= 32'sh0;
    end else begin
      last_acc_write_0_12 <= add_0_12;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_13 <= 32'sh0;
    end else begin
      last_acc_write_0_13 <= add_0_13;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_14 <= 32'sh0;
    end else begin
      last_acc_write_0_14 <= add_0_14;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_15 <= 32'sh0;
    end else begin
      last_acc_write_0_15 <= add_0_15;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_16 <= 32'sh0;
    end else begin
      last_acc_write_0_16 <= add_0_16;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_17 <= 32'sh0;
    end else begin
      last_acc_write_0_17 <= add_0_17;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_18 <= 32'sh0;
    end else begin
      last_acc_write_0_18 <= add_0_18;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_19 <= 32'sh0;
    end else begin
      last_acc_write_0_19 <= add_0_19;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_20 <= 32'sh0;
    end else begin
      last_acc_write_0_20 <= add_0_20;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_21 <= 32'sh0;
    end else begin
      last_acc_write_0_21 <= add_0_21;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_22 <= 32'sh0;
    end else begin
      last_acc_write_0_22 <= add_0_22;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_23 <= 32'sh0;
    end else begin
      last_acc_write_0_23 <= add_0_23;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_24 <= 32'sh0;
    end else begin
      last_acc_write_0_24 <= add_0_24;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_25 <= 32'sh0;
    end else begin
      last_acc_write_0_25 <= add_0_25;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_26 <= 32'sh0;
    end else begin
      last_acc_write_0_26 <= add_0_26;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_27 <= 32'sh0;
    end else begin
      last_acc_write_0_27 <= add_0_27;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_28 <= 32'sh0;
    end else begin
      last_acc_write_0_28 <= add_0_28;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_29 <= 32'sh0;
    end else begin
      last_acc_write_0_29 <= add_0_29;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_30 <= 32'sh0;
    end else begin
      last_acc_write_0_30 <= add_0_30;
    end
    if (io_valid_reset) begin // @[TensorGemm.scala 210:20]
      last_acc_write_0_31 <= 32'sh0;
    end else begin
      last_acc_write_0_31 <= add_0_31;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  last_acc_write_0_0 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  last_acc_write_0_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  last_acc_write_0_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  last_acc_write_0_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  last_acc_write_0_4 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  last_acc_write_0_5 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  last_acc_write_0_6 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  last_acc_write_0_7 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  last_acc_write_0_8 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  last_acc_write_0_9 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  last_acc_write_0_10 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  last_acc_write_0_11 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  last_acc_write_0_12 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  last_acc_write_0_13 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  last_acc_write_0_14 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  last_acc_write_0_15 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  last_acc_write_0_16 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  last_acc_write_0_17 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  last_acc_write_0_18 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  last_acc_write_0_19 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  last_acc_write_0_20 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  last_acc_write_0_21 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  last_acc_write_0_22 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  last_acc_write_0_23 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  last_acc_write_0_24 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  last_acc_write_0_25 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  last_acc_write_0_26 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  last_acc_write_0_27 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  last_acc_write_0_28 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  last_acc_write_0_29 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  last_acc_write_0_30 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  last_acc_write_0_31 = _RAND_31[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module TensorGemm(
  input         clock,
  input         reset,
  input         io_start,
  output        io_done,
  input  [9:0]  io_dec_wgt_1,
  input  [9:0]  io_dec_wgt_0,
  input  [10:0] io_dec_inp_1,
  input  [10:0] io_dec_inp_0,
  input  [10:0] io_dec_acc_1,
  input  [10:0] io_dec_acc_0,
  input         io_dec_empty_0,
  input  [13:0] io_dec_lp_1,
  input  [13:0] io_dec_lp_0,
  input  [13:0] io_dec_uop_end,
  input  [12:0] io_dec_uop_begin,
  input         io_dec_reset,
  input         io_dec_push_next,
  input         io_dec_push_prev,
  input         io_dec_pop_next,
  input         io_dec_pop_prev,
  input  [2:0]  io_dec_op,
  output        io_uop_idx_valid,
  output [6:0]  io_uop_idx_bits,
  input         io_uop_data_valid,
  input  [9:0]  io_uop_data_bits_u2,
  input  [10:0] io_uop_data_bits_u1,
  input  [10:0] io_uop_data_bits_u0,
  output        io_inp_rd_0_idx_valid,
  output [6:0]  io_inp_rd_0_idx_bits,
  input         io_inp_rd_0_data_valid,
  input  [7:0]  io_inp_rd_0_data_bits_0_0,
  input  [7:0]  io_inp_rd_0_data_bits_0_1,
  input  [7:0]  io_inp_rd_0_data_bits_0_2,
  input  [7:0]  io_inp_rd_0_data_bits_0_3,
  input  [7:0]  io_inp_rd_0_data_bits_0_4,
  input  [7:0]  io_inp_rd_0_data_bits_0_5,
  input  [7:0]  io_inp_rd_0_data_bits_0_6,
  input  [7:0]  io_inp_rd_0_data_bits_0_7,
  input  [7:0]  io_inp_rd_0_data_bits_0_8,
  input  [7:0]  io_inp_rd_0_data_bits_0_9,
  input  [7:0]  io_inp_rd_0_data_bits_0_10,
  input  [7:0]  io_inp_rd_0_data_bits_0_11,
  input  [7:0]  io_inp_rd_0_data_bits_0_12,
  input  [7:0]  io_inp_rd_0_data_bits_0_13,
  input  [7:0]  io_inp_rd_0_data_bits_0_14,
  input  [7:0]  io_inp_rd_0_data_bits_0_15,
  output        io_wgt_rd_0_idx_valid,
  output [5:0]  io_wgt_rd_0_idx_bits,
  input         io_wgt_rd_0_data_valid,
  input  [7:0]  io_wgt_rd_0_data_bits_0_0,
  input  [7:0]  io_wgt_rd_0_data_bits_0_1,
  input  [7:0]  io_wgt_rd_0_data_bits_0_2,
  input  [7:0]  io_wgt_rd_0_data_bits_0_3,
  input  [7:0]  io_wgt_rd_0_data_bits_0_4,
  input  [7:0]  io_wgt_rd_0_data_bits_0_5,
  input  [7:0]  io_wgt_rd_0_data_bits_0_6,
  input  [7:0]  io_wgt_rd_0_data_bits_0_7,
  input  [7:0]  io_wgt_rd_0_data_bits_0_8,
  input  [7:0]  io_wgt_rd_0_data_bits_0_9,
  input  [7:0]  io_wgt_rd_0_data_bits_0_10,
  input  [7:0]  io_wgt_rd_0_data_bits_0_11,
  input  [7:0]  io_wgt_rd_0_data_bits_0_12,
  input  [7:0]  io_wgt_rd_0_data_bits_0_13,
  input  [7:0]  io_wgt_rd_0_data_bits_0_14,
  input  [7:0]  io_wgt_rd_0_data_bits_0_15,
  input  [7:0]  io_wgt_rd_0_data_bits_1_0,
  input  [7:0]  io_wgt_rd_0_data_bits_1_1,
  input  [7:0]  io_wgt_rd_0_data_bits_1_2,
  input  [7:0]  io_wgt_rd_0_data_bits_1_3,
  input  [7:0]  io_wgt_rd_0_data_bits_1_4,
  input  [7:0]  io_wgt_rd_0_data_bits_1_5,
  input  [7:0]  io_wgt_rd_0_data_bits_1_6,
  input  [7:0]  io_wgt_rd_0_data_bits_1_7,
  input  [7:0]  io_wgt_rd_0_data_bits_1_8,
  input  [7:0]  io_wgt_rd_0_data_bits_1_9,
  input  [7:0]  io_wgt_rd_0_data_bits_1_10,
  input  [7:0]  io_wgt_rd_0_data_bits_1_11,
  input  [7:0]  io_wgt_rd_0_data_bits_1_12,
  input  [7:0]  io_wgt_rd_0_data_bits_1_13,
  input  [7:0]  io_wgt_rd_0_data_bits_1_14,
  input  [7:0]  io_wgt_rd_0_data_bits_1_15,
  input  [7:0]  io_wgt_rd_0_data_bits_2_0,
  input  [7:0]  io_wgt_rd_0_data_bits_2_1,
  input  [7:0]  io_wgt_rd_0_data_bits_2_2,
  input  [7:0]  io_wgt_rd_0_data_bits_2_3,
  input  [7:0]  io_wgt_rd_0_data_bits_2_4,
  input  [7:0]  io_wgt_rd_0_data_bits_2_5,
  input  [7:0]  io_wgt_rd_0_data_bits_2_6,
  input  [7:0]  io_wgt_rd_0_data_bits_2_7,
  input  [7:0]  io_wgt_rd_0_data_bits_2_8,
  input  [7:0]  io_wgt_rd_0_data_bits_2_9,
  input  [7:0]  io_wgt_rd_0_data_bits_2_10,
  input  [7:0]  io_wgt_rd_0_data_bits_2_11,
  input  [7:0]  io_wgt_rd_0_data_bits_2_12,
  input  [7:0]  io_wgt_rd_0_data_bits_2_13,
  input  [7:0]  io_wgt_rd_0_data_bits_2_14,
  input  [7:0]  io_wgt_rd_0_data_bits_2_15,
  input  [7:0]  io_wgt_rd_0_data_bits_3_0,
  input  [7:0]  io_wgt_rd_0_data_bits_3_1,
  input  [7:0]  io_wgt_rd_0_data_bits_3_2,
  input  [7:0]  io_wgt_rd_0_data_bits_3_3,
  input  [7:0]  io_wgt_rd_0_data_bits_3_4,
  input  [7:0]  io_wgt_rd_0_data_bits_3_5,
  input  [7:0]  io_wgt_rd_0_data_bits_3_6,
  input  [7:0]  io_wgt_rd_0_data_bits_3_7,
  input  [7:0]  io_wgt_rd_0_data_bits_3_8,
  input  [7:0]  io_wgt_rd_0_data_bits_3_9,
  input  [7:0]  io_wgt_rd_0_data_bits_3_10,
  input  [7:0]  io_wgt_rd_0_data_bits_3_11,
  input  [7:0]  io_wgt_rd_0_data_bits_3_12,
  input  [7:0]  io_wgt_rd_0_data_bits_3_13,
  input  [7:0]  io_wgt_rd_0_data_bits_3_14,
  input  [7:0]  io_wgt_rd_0_data_bits_3_15,
  input  [7:0]  io_wgt_rd_0_data_bits_4_0,
  input  [7:0]  io_wgt_rd_0_data_bits_4_1,
  input  [7:0]  io_wgt_rd_0_data_bits_4_2,
  input  [7:0]  io_wgt_rd_0_data_bits_4_3,
  input  [7:0]  io_wgt_rd_0_data_bits_4_4,
  input  [7:0]  io_wgt_rd_0_data_bits_4_5,
  input  [7:0]  io_wgt_rd_0_data_bits_4_6,
  input  [7:0]  io_wgt_rd_0_data_bits_4_7,
  input  [7:0]  io_wgt_rd_0_data_bits_4_8,
  input  [7:0]  io_wgt_rd_0_data_bits_4_9,
  input  [7:0]  io_wgt_rd_0_data_bits_4_10,
  input  [7:0]  io_wgt_rd_0_data_bits_4_11,
  input  [7:0]  io_wgt_rd_0_data_bits_4_12,
  input  [7:0]  io_wgt_rd_0_data_bits_4_13,
  input  [7:0]  io_wgt_rd_0_data_bits_4_14,
  input  [7:0]  io_wgt_rd_0_data_bits_4_15,
  input  [7:0]  io_wgt_rd_0_data_bits_5_0,
  input  [7:0]  io_wgt_rd_0_data_bits_5_1,
  input  [7:0]  io_wgt_rd_0_data_bits_5_2,
  input  [7:0]  io_wgt_rd_0_data_bits_5_3,
  input  [7:0]  io_wgt_rd_0_data_bits_5_4,
  input  [7:0]  io_wgt_rd_0_data_bits_5_5,
  input  [7:0]  io_wgt_rd_0_data_bits_5_6,
  input  [7:0]  io_wgt_rd_0_data_bits_5_7,
  input  [7:0]  io_wgt_rd_0_data_bits_5_8,
  input  [7:0]  io_wgt_rd_0_data_bits_5_9,
  input  [7:0]  io_wgt_rd_0_data_bits_5_10,
  input  [7:0]  io_wgt_rd_0_data_bits_5_11,
  input  [7:0]  io_wgt_rd_0_data_bits_5_12,
  input  [7:0]  io_wgt_rd_0_data_bits_5_13,
  input  [7:0]  io_wgt_rd_0_data_bits_5_14,
  input  [7:0]  io_wgt_rd_0_data_bits_5_15,
  input  [7:0]  io_wgt_rd_0_data_bits_6_0,
  input  [7:0]  io_wgt_rd_0_data_bits_6_1,
  input  [7:0]  io_wgt_rd_0_data_bits_6_2,
  input  [7:0]  io_wgt_rd_0_data_bits_6_3,
  input  [7:0]  io_wgt_rd_0_data_bits_6_4,
  input  [7:0]  io_wgt_rd_0_data_bits_6_5,
  input  [7:0]  io_wgt_rd_0_data_bits_6_6,
  input  [7:0]  io_wgt_rd_0_data_bits_6_7,
  input  [7:0]  io_wgt_rd_0_data_bits_6_8,
  input  [7:0]  io_wgt_rd_0_data_bits_6_9,
  input  [7:0]  io_wgt_rd_0_data_bits_6_10,
  input  [7:0]  io_wgt_rd_0_data_bits_6_11,
  input  [7:0]  io_wgt_rd_0_data_bits_6_12,
  input  [7:0]  io_wgt_rd_0_data_bits_6_13,
  input  [7:0]  io_wgt_rd_0_data_bits_6_14,
  input  [7:0]  io_wgt_rd_0_data_bits_6_15,
  input  [7:0]  io_wgt_rd_0_data_bits_7_0,
  input  [7:0]  io_wgt_rd_0_data_bits_7_1,
  input  [7:0]  io_wgt_rd_0_data_bits_7_2,
  input  [7:0]  io_wgt_rd_0_data_bits_7_3,
  input  [7:0]  io_wgt_rd_0_data_bits_7_4,
  input  [7:0]  io_wgt_rd_0_data_bits_7_5,
  input  [7:0]  io_wgt_rd_0_data_bits_7_6,
  input  [7:0]  io_wgt_rd_0_data_bits_7_7,
  input  [7:0]  io_wgt_rd_0_data_bits_7_8,
  input  [7:0]  io_wgt_rd_0_data_bits_7_9,
  input  [7:0]  io_wgt_rd_0_data_bits_7_10,
  input  [7:0]  io_wgt_rd_0_data_bits_7_11,
  input  [7:0]  io_wgt_rd_0_data_bits_7_12,
  input  [7:0]  io_wgt_rd_0_data_bits_7_13,
  input  [7:0]  io_wgt_rd_0_data_bits_7_14,
  input  [7:0]  io_wgt_rd_0_data_bits_7_15,
  input  [7:0]  io_wgt_rd_0_data_bits_8_0,
  input  [7:0]  io_wgt_rd_0_data_bits_8_1,
  input  [7:0]  io_wgt_rd_0_data_bits_8_2,
  input  [7:0]  io_wgt_rd_0_data_bits_8_3,
  input  [7:0]  io_wgt_rd_0_data_bits_8_4,
  input  [7:0]  io_wgt_rd_0_data_bits_8_5,
  input  [7:0]  io_wgt_rd_0_data_bits_8_6,
  input  [7:0]  io_wgt_rd_0_data_bits_8_7,
  input  [7:0]  io_wgt_rd_0_data_bits_8_8,
  input  [7:0]  io_wgt_rd_0_data_bits_8_9,
  input  [7:0]  io_wgt_rd_0_data_bits_8_10,
  input  [7:0]  io_wgt_rd_0_data_bits_8_11,
  input  [7:0]  io_wgt_rd_0_data_bits_8_12,
  input  [7:0]  io_wgt_rd_0_data_bits_8_13,
  input  [7:0]  io_wgt_rd_0_data_bits_8_14,
  input  [7:0]  io_wgt_rd_0_data_bits_8_15,
  input  [7:0]  io_wgt_rd_0_data_bits_9_0,
  input  [7:0]  io_wgt_rd_0_data_bits_9_1,
  input  [7:0]  io_wgt_rd_0_data_bits_9_2,
  input  [7:0]  io_wgt_rd_0_data_bits_9_3,
  input  [7:0]  io_wgt_rd_0_data_bits_9_4,
  input  [7:0]  io_wgt_rd_0_data_bits_9_5,
  input  [7:0]  io_wgt_rd_0_data_bits_9_6,
  input  [7:0]  io_wgt_rd_0_data_bits_9_7,
  input  [7:0]  io_wgt_rd_0_data_bits_9_8,
  input  [7:0]  io_wgt_rd_0_data_bits_9_9,
  input  [7:0]  io_wgt_rd_0_data_bits_9_10,
  input  [7:0]  io_wgt_rd_0_data_bits_9_11,
  input  [7:0]  io_wgt_rd_0_data_bits_9_12,
  input  [7:0]  io_wgt_rd_0_data_bits_9_13,
  input  [7:0]  io_wgt_rd_0_data_bits_9_14,
  input  [7:0]  io_wgt_rd_0_data_bits_9_15,
  input  [7:0]  io_wgt_rd_0_data_bits_10_0,
  input  [7:0]  io_wgt_rd_0_data_bits_10_1,
  input  [7:0]  io_wgt_rd_0_data_bits_10_2,
  input  [7:0]  io_wgt_rd_0_data_bits_10_3,
  input  [7:0]  io_wgt_rd_0_data_bits_10_4,
  input  [7:0]  io_wgt_rd_0_data_bits_10_5,
  input  [7:0]  io_wgt_rd_0_data_bits_10_6,
  input  [7:0]  io_wgt_rd_0_data_bits_10_7,
  input  [7:0]  io_wgt_rd_0_data_bits_10_8,
  input  [7:0]  io_wgt_rd_0_data_bits_10_9,
  input  [7:0]  io_wgt_rd_0_data_bits_10_10,
  input  [7:0]  io_wgt_rd_0_data_bits_10_11,
  input  [7:0]  io_wgt_rd_0_data_bits_10_12,
  input  [7:0]  io_wgt_rd_0_data_bits_10_13,
  input  [7:0]  io_wgt_rd_0_data_bits_10_14,
  input  [7:0]  io_wgt_rd_0_data_bits_10_15,
  input  [7:0]  io_wgt_rd_0_data_bits_11_0,
  input  [7:0]  io_wgt_rd_0_data_bits_11_1,
  input  [7:0]  io_wgt_rd_0_data_bits_11_2,
  input  [7:0]  io_wgt_rd_0_data_bits_11_3,
  input  [7:0]  io_wgt_rd_0_data_bits_11_4,
  input  [7:0]  io_wgt_rd_0_data_bits_11_5,
  input  [7:0]  io_wgt_rd_0_data_bits_11_6,
  input  [7:0]  io_wgt_rd_0_data_bits_11_7,
  input  [7:0]  io_wgt_rd_0_data_bits_11_8,
  input  [7:0]  io_wgt_rd_0_data_bits_11_9,
  input  [7:0]  io_wgt_rd_0_data_bits_11_10,
  input  [7:0]  io_wgt_rd_0_data_bits_11_11,
  input  [7:0]  io_wgt_rd_0_data_bits_11_12,
  input  [7:0]  io_wgt_rd_0_data_bits_11_13,
  input  [7:0]  io_wgt_rd_0_data_bits_11_14,
  input  [7:0]  io_wgt_rd_0_data_bits_11_15,
  input  [7:0]  io_wgt_rd_0_data_bits_12_0,
  input  [7:0]  io_wgt_rd_0_data_bits_12_1,
  input  [7:0]  io_wgt_rd_0_data_bits_12_2,
  input  [7:0]  io_wgt_rd_0_data_bits_12_3,
  input  [7:0]  io_wgt_rd_0_data_bits_12_4,
  input  [7:0]  io_wgt_rd_0_data_bits_12_5,
  input  [7:0]  io_wgt_rd_0_data_bits_12_6,
  input  [7:0]  io_wgt_rd_0_data_bits_12_7,
  input  [7:0]  io_wgt_rd_0_data_bits_12_8,
  input  [7:0]  io_wgt_rd_0_data_bits_12_9,
  input  [7:0]  io_wgt_rd_0_data_bits_12_10,
  input  [7:0]  io_wgt_rd_0_data_bits_12_11,
  input  [7:0]  io_wgt_rd_0_data_bits_12_12,
  input  [7:0]  io_wgt_rd_0_data_bits_12_13,
  input  [7:0]  io_wgt_rd_0_data_bits_12_14,
  input  [7:0]  io_wgt_rd_0_data_bits_12_15,
  input  [7:0]  io_wgt_rd_0_data_bits_13_0,
  input  [7:0]  io_wgt_rd_0_data_bits_13_1,
  input  [7:0]  io_wgt_rd_0_data_bits_13_2,
  input  [7:0]  io_wgt_rd_0_data_bits_13_3,
  input  [7:0]  io_wgt_rd_0_data_bits_13_4,
  input  [7:0]  io_wgt_rd_0_data_bits_13_5,
  input  [7:0]  io_wgt_rd_0_data_bits_13_6,
  input  [7:0]  io_wgt_rd_0_data_bits_13_7,
  input  [7:0]  io_wgt_rd_0_data_bits_13_8,
  input  [7:0]  io_wgt_rd_0_data_bits_13_9,
  input  [7:0]  io_wgt_rd_0_data_bits_13_10,
  input  [7:0]  io_wgt_rd_0_data_bits_13_11,
  input  [7:0]  io_wgt_rd_0_data_bits_13_12,
  input  [7:0]  io_wgt_rd_0_data_bits_13_13,
  input  [7:0]  io_wgt_rd_0_data_bits_13_14,
  input  [7:0]  io_wgt_rd_0_data_bits_13_15,
  input  [7:0]  io_wgt_rd_0_data_bits_14_0,
  input  [7:0]  io_wgt_rd_0_data_bits_14_1,
  input  [7:0]  io_wgt_rd_0_data_bits_14_2,
  input  [7:0]  io_wgt_rd_0_data_bits_14_3,
  input  [7:0]  io_wgt_rd_0_data_bits_14_4,
  input  [7:0]  io_wgt_rd_0_data_bits_14_5,
  input  [7:0]  io_wgt_rd_0_data_bits_14_6,
  input  [7:0]  io_wgt_rd_0_data_bits_14_7,
  input  [7:0]  io_wgt_rd_0_data_bits_14_8,
  input  [7:0]  io_wgt_rd_0_data_bits_14_9,
  input  [7:0]  io_wgt_rd_0_data_bits_14_10,
  input  [7:0]  io_wgt_rd_0_data_bits_14_11,
  input  [7:0]  io_wgt_rd_0_data_bits_14_12,
  input  [7:0]  io_wgt_rd_0_data_bits_14_13,
  input  [7:0]  io_wgt_rd_0_data_bits_14_14,
  input  [7:0]  io_wgt_rd_0_data_bits_14_15,
  input  [7:0]  io_wgt_rd_0_data_bits_15_0,
  input  [7:0]  io_wgt_rd_0_data_bits_15_1,
  input  [7:0]  io_wgt_rd_0_data_bits_15_2,
  input  [7:0]  io_wgt_rd_0_data_bits_15_3,
  input  [7:0]  io_wgt_rd_0_data_bits_15_4,
  input  [7:0]  io_wgt_rd_0_data_bits_15_5,
  input  [7:0]  io_wgt_rd_0_data_bits_15_6,
  input  [7:0]  io_wgt_rd_0_data_bits_15_7,
  input  [7:0]  io_wgt_rd_0_data_bits_15_8,
  input  [7:0]  io_wgt_rd_0_data_bits_15_9,
  input  [7:0]  io_wgt_rd_0_data_bits_15_10,
  input  [7:0]  io_wgt_rd_0_data_bits_15_11,
  input  [7:0]  io_wgt_rd_0_data_bits_15_12,
  input  [7:0]  io_wgt_rd_0_data_bits_15_13,
  input  [7:0]  io_wgt_rd_0_data_bits_15_14,
  input  [7:0]  io_wgt_rd_0_data_bits_15_15,
  input  [7:0]  io_wgt_rd_0_data_bits_16_0,
  input  [7:0]  io_wgt_rd_0_data_bits_16_1,
  input  [7:0]  io_wgt_rd_0_data_bits_16_2,
  input  [7:0]  io_wgt_rd_0_data_bits_16_3,
  input  [7:0]  io_wgt_rd_0_data_bits_16_4,
  input  [7:0]  io_wgt_rd_0_data_bits_16_5,
  input  [7:0]  io_wgt_rd_0_data_bits_16_6,
  input  [7:0]  io_wgt_rd_0_data_bits_16_7,
  input  [7:0]  io_wgt_rd_0_data_bits_16_8,
  input  [7:0]  io_wgt_rd_0_data_bits_16_9,
  input  [7:0]  io_wgt_rd_0_data_bits_16_10,
  input  [7:0]  io_wgt_rd_0_data_bits_16_11,
  input  [7:0]  io_wgt_rd_0_data_bits_16_12,
  input  [7:0]  io_wgt_rd_0_data_bits_16_13,
  input  [7:0]  io_wgt_rd_0_data_bits_16_14,
  input  [7:0]  io_wgt_rd_0_data_bits_16_15,
  input  [7:0]  io_wgt_rd_0_data_bits_17_0,
  input  [7:0]  io_wgt_rd_0_data_bits_17_1,
  input  [7:0]  io_wgt_rd_0_data_bits_17_2,
  input  [7:0]  io_wgt_rd_0_data_bits_17_3,
  input  [7:0]  io_wgt_rd_0_data_bits_17_4,
  input  [7:0]  io_wgt_rd_0_data_bits_17_5,
  input  [7:0]  io_wgt_rd_0_data_bits_17_6,
  input  [7:0]  io_wgt_rd_0_data_bits_17_7,
  input  [7:0]  io_wgt_rd_0_data_bits_17_8,
  input  [7:0]  io_wgt_rd_0_data_bits_17_9,
  input  [7:0]  io_wgt_rd_0_data_bits_17_10,
  input  [7:0]  io_wgt_rd_0_data_bits_17_11,
  input  [7:0]  io_wgt_rd_0_data_bits_17_12,
  input  [7:0]  io_wgt_rd_0_data_bits_17_13,
  input  [7:0]  io_wgt_rd_0_data_bits_17_14,
  input  [7:0]  io_wgt_rd_0_data_bits_17_15,
  input  [7:0]  io_wgt_rd_0_data_bits_18_0,
  input  [7:0]  io_wgt_rd_0_data_bits_18_1,
  input  [7:0]  io_wgt_rd_0_data_bits_18_2,
  input  [7:0]  io_wgt_rd_0_data_bits_18_3,
  input  [7:0]  io_wgt_rd_0_data_bits_18_4,
  input  [7:0]  io_wgt_rd_0_data_bits_18_5,
  input  [7:0]  io_wgt_rd_0_data_bits_18_6,
  input  [7:0]  io_wgt_rd_0_data_bits_18_7,
  input  [7:0]  io_wgt_rd_0_data_bits_18_8,
  input  [7:0]  io_wgt_rd_0_data_bits_18_9,
  input  [7:0]  io_wgt_rd_0_data_bits_18_10,
  input  [7:0]  io_wgt_rd_0_data_bits_18_11,
  input  [7:0]  io_wgt_rd_0_data_bits_18_12,
  input  [7:0]  io_wgt_rd_0_data_bits_18_13,
  input  [7:0]  io_wgt_rd_0_data_bits_18_14,
  input  [7:0]  io_wgt_rd_0_data_bits_18_15,
  input  [7:0]  io_wgt_rd_0_data_bits_19_0,
  input  [7:0]  io_wgt_rd_0_data_bits_19_1,
  input  [7:0]  io_wgt_rd_0_data_bits_19_2,
  input  [7:0]  io_wgt_rd_0_data_bits_19_3,
  input  [7:0]  io_wgt_rd_0_data_bits_19_4,
  input  [7:0]  io_wgt_rd_0_data_bits_19_5,
  input  [7:0]  io_wgt_rd_0_data_bits_19_6,
  input  [7:0]  io_wgt_rd_0_data_bits_19_7,
  input  [7:0]  io_wgt_rd_0_data_bits_19_8,
  input  [7:0]  io_wgt_rd_0_data_bits_19_9,
  input  [7:0]  io_wgt_rd_0_data_bits_19_10,
  input  [7:0]  io_wgt_rd_0_data_bits_19_11,
  input  [7:0]  io_wgt_rd_0_data_bits_19_12,
  input  [7:0]  io_wgt_rd_0_data_bits_19_13,
  input  [7:0]  io_wgt_rd_0_data_bits_19_14,
  input  [7:0]  io_wgt_rd_0_data_bits_19_15,
  input  [7:0]  io_wgt_rd_0_data_bits_20_0,
  input  [7:0]  io_wgt_rd_0_data_bits_20_1,
  input  [7:0]  io_wgt_rd_0_data_bits_20_2,
  input  [7:0]  io_wgt_rd_0_data_bits_20_3,
  input  [7:0]  io_wgt_rd_0_data_bits_20_4,
  input  [7:0]  io_wgt_rd_0_data_bits_20_5,
  input  [7:0]  io_wgt_rd_0_data_bits_20_6,
  input  [7:0]  io_wgt_rd_0_data_bits_20_7,
  input  [7:0]  io_wgt_rd_0_data_bits_20_8,
  input  [7:0]  io_wgt_rd_0_data_bits_20_9,
  input  [7:0]  io_wgt_rd_0_data_bits_20_10,
  input  [7:0]  io_wgt_rd_0_data_bits_20_11,
  input  [7:0]  io_wgt_rd_0_data_bits_20_12,
  input  [7:0]  io_wgt_rd_0_data_bits_20_13,
  input  [7:0]  io_wgt_rd_0_data_bits_20_14,
  input  [7:0]  io_wgt_rd_0_data_bits_20_15,
  input  [7:0]  io_wgt_rd_0_data_bits_21_0,
  input  [7:0]  io_wgt_rd_0_data_bits_21_1,
  input  [7:0]  io_wgt_rd_0_data_bits_21_2,
  input  [7:0]  io_wgt_rd_0_data_bits_21_3,
  input  [7:0]  io_wgt_rd_0_data_bits_21_4,
  input  [7:0]  io_wgt_rd_0_data_bits_21_5,
  input  [7:0]  io_wgt_rd_0_data_bits_21_6,
  input  [7:0]  io_wgt_rd_0_data_bits_21_7,
  input  [7:0]  io_wgt_rd_0_data_bits_21_8,
  input  [7:0]  io_wgt_rd_0_data_bits_21_9,
  input  [7:0]  io_wgt_rd_0_data_bits_21_10,
  input  [7:0]  io_wgt_rd_0_data_bits_21_11,
  input  [7:0]  io_wgt_rd_0_data_bits_21_12,
  input  [7:0]  io_wgt_rd_0_data_bits_21_13,
  input  [7:0]  io_wgt_rd_0_data_bits_21_14,
  input  [7:0]  io_wgt_rd_0_data_bits_21_15,
  input  [7:0]  io_wgt_rd_0_data_bits_22_0,
  input  [7:0]  io_wgt_rd_0_data_bits_22_1,
  input  [7:0]  io_wgt_rd_0_data_bits_22_2,
  input  [7:0]  io_wgt_rd_0_data_bits_22_3,
  input  [7:0]  io_wgt_rd_0_data_bits_22_4,
  input  [7:0]  io_wgt_rd_0_data_bits_22_5,
  input  [7:0]  io_wgt_rd_0_data_bits_22_6,
  input  [7:0]  io_wgt_rd_0_data_bits_22_7,
  input  [7:0]  io_wgt_rd_0_data_bits_22_8,
  input  [7:0]  io_wgt_rd_0_data_bits_22_9,
  input  [7:0]  io_wgt_rd_0_data_bits_22_10,
  input  [7:0]  io_wgt_rd_0_data_bits_22_11,
  input  [7:0]  io_wgt_rd_0_data_bits_22_12,
  input  [7:0]  io_wgt_rd_0_data_bits_22_13,
  input  [7:0]  io_wgt_rd_0_data_bits_22_14,
  input  [7:0]  io_wgt_rd_0_data_bits_22_15,
  input  [7:0]  io_wgt_rd_0_data_bits_23_0,
  input  [7:0]  io_wgt_rd_0_data_bits_23_1,
  input  [7:0]  io_wgt_rd_0_data_bits_23_2,
  input  [7:0]  io_wgt_rd_0_data_bits_23_3,
  input  [7:0]  io_wgt_rd_0_data_bits_23_4,
  input  [7:0]  io_wgt_rd_0_data_bits_23_5,
  input  [7:0]  io_wgt_rd_0_data_bits_23_6,
  input  [7:0]  io_wgt_rd_0_data_bits_23_7,
  input  [7:0]  io_wgt_rd_0_data_bits_23_8,
  input  [7:0]  io_wgt_rd_0_data_bits_23_9,
  input  [7:0]  io_wgt_rd_0_data_bits_23_10,
  input  [7:0]  io_wgt_rd_0_data_bits_23_11,
  input  [7:0]  io_wgt_rd_0_data_bits_23_12,
  input  [7:0]  io_wgt_rd_0_data_bits_23_13,
  input  [7:0]  io_wgt_rd_0_data_bits_23_14,
  input  [7:0]  io_wgt_rd_0_data_bits_23_15,
  input  [7:0]  io_wgt_rd_0_data_bits_24_0,
  input  [7:0]  io_wgt_rd_0_data_bits_24_1,
  input  [7:0]  io_wgt_rd_0_data_bits_24_2,
  input  [7:0]  io_wgt_rd_0_data_bits_24_3,
  input  [7:0]  io_wgt_rd_0_data_bits_24_4,
  input  [7:0]  io_wgt_rd_0_data_bits_24_5,
  input  [7:0]  io_wgt_rd_0_data_bits_24_6,
  input  [7:0]  io_wgt_rd_0_data_bits_24_7,
  input  [7:0]  io_wgt_rd_0_data_bits_24_8,
  input  [7:0]  io_wgt_rd_0_data_bits_24_9,
  input  [7:0]  io_wgt_rd_0_data_bits_24_10,
  input  [7:0]  io_wgt_rd_0_data_bits_24_11,
  input  [7:0]  io_wgt_rd_0_data_bits_24_12,
  input  [7:0]  io_wgt_rd_0_data_bits_24_13,
  input  [7:0]  io_wgt_rd_0_data_bits_24_14,
  input  [7:0]  io_wgt_rd_0_data_bits_24_15,
  input  [7:0]  io_wgt_rd_0_data_bits_25_0,
  input  [7:0]  io_wgt_rd_0_data_bits_25_1,
  input  [7:0]  io_wgt_rd_0_data_bits_25_2,
  input  [7:0]  io_wgt_rd_0_data_bits_25_3,
  input  [7:0]  io_wgt_rd_0_data_bits_25_4,
  input  [7:0]  io_wgt_rd_0_data_bits_25_5,
  input  [7:0]  io_wgt_rd_0_data_bits_25_6,
  input  [7:0]  io_wgt_rd_0_data_bits_25_7,
  input  [7:0]  io_wgt_rd_0_data_bits_25_8,
  input  [7:0]  io_wgt_rd_0_data_bits_25_9,
  input  [7:0]  io_wgt_rd_0_data_bits_25_10,
  input  [7:0]  io_wgt_rd_0_data_bits_25_11,
  input  [7:0]  io_wgt_rd_0_data_bits_25_12,
  input  [7:0]  io_wgt_rd_0_data_bits_25_13,
  input  [7:0]  io_wgt_rd_0_data_bits_25_14,
  input  [7:0]  io_wgt_rd_0_data_bits_25_15,
  input  [7:0]  io_wgt_rd_0_data_bits_26_0,
  input  [7:0]  io_wgt_rd_0_data_bits_26_1,
  input  [7:0]  io_wgt_rd_0_data_bits_26_2,
  input  [7:0]  io_wgt_rd_0_data_bits_26_3,
  input  [7:0]  io_wgt_rd_0_data_bits_26_4,
  input  [7:0]  io_wgt_rd_0_data_bits_26_5,
  input  [7:0]  io_wgt_rd_0_data_bits_26_6,
  input  [7:0]  io_wgt_rd_0_data_bits_26_7,
  input  [7:0]  io_wgt_rd_0_data_bits_26_8,
  input  [7:0]  io_wgt_rd_0_data_bits_26_9,
  input  [7:0]  io_wgt_rd_0_data_bits_26_10,
  input  [7:0]  io_wgt_rd_0_data_bits_26_11,
  input  [7:0]  io_wgt_rd_0_data_bits_26_12,
  input  [7:0]  io_wgt_rd_0_data_bits_26_13,
  input  [7:0]  io_wgt_rd_0_data_bits_26_14,
  input  [7:0]  io_wgt_rd_0_data_bits_26_15,
  input  [7:0]  io_wgt_rd_0_data_bits_27_0,
  input  [7:0]  io_wgt_rd_0_data_bits_27_1,
  input  [7:0]  io_wgt_rd_0_data_bits_27_2,
  input  [7:0]  io_wgt_rd_0_data_bits_27_3,
  input  [7:0]  io_wgt_rd_0_data_bits_27_4,
  input  [7:0]  io_wgt_rd_0_data_bits_27_5,
  input  [7:0]  io_wgt_rd_0_data_bits_27_6,
  input  [7:0]  io_wgt_rd_0_data_bits_27_7,
  input  [7:0]  io_wgt_rd_0_data_bits_27_8,
  input  [7:0]  io_wgt_rd_0_data_bits_27_9,
  input  [7:0]  io_wgt_rd_0_data_bits_27_10,
  input  [7:0]  io_wgt_rd_0_data_bits_27_11,
  input  [7:0]  io_wgt_rd_0_data_bits_27_12,
  input  [7:0]  io_wgt_rd_0_data_bits_27_13,
  input  [7:0]  io_wgt_rd_0_data_bits_27_14,
  input  [7:0]  io_wgt_rd_0_data_bits_27_15,
  input  [7:0]  io_wgt_rd_0_data_bits_28_0,
  input  [7:0]  io_wgt_rd_0_data_bits_28_1,
  input  [7:0]  io_wgt_rd_0_data_bits_28_2,
  input  [7:0]  io_wgt_rd_0_data_bits_28_3,
  input  [7:0]  io_wgt_rd_0_data_bits_28_4,
  input  [7:0]  io_wgt_rd_0_data_bits_28_5,
  input  [7:0]  io_wgt_rd_0_data_bits_28_6,
  input  [7:0]  io_wgt_rd_0_data_bits_28_7,
  input  [7:0]  io_wgt_rd_0_data_bits_28_8,
  input  [7:0]  io_wgt_rd_0_data_bits_28_9,
  input  [7:0]  io_wgt_rd_0_data_bits_28_10,
  input  [7:0]  io_wgt_rd_0_data_bits_28_11,
  input  [7:0]  io_wgt_rd_0_data_bits_28_12,
  input  [7:0]  io_wgt_rd_0_data_bits_28_13,
  input  [7:0]  io_wgt_rd_0_data_bits_28_14,
  input  [7:0]  io_wgt_rd_0_data_bits_28_15,
  input  [7:0]  io_wgt_rd_0_data_bits_29_0,
  input  [7:0]  io_wgt_rd_0_data_bits_29_1,
  input  [7:0]  io_wgt_rd_0_data_bits_29_2,
  input  [7:0]  io_wgt_rd_0_data_bits_29_3,
  input  [7:0]  io_wgt_rd_0_data_bits_29_4,
  input  [7:0]  io_wgt_rd_0_data_bits_29_5,
  input  [7:0]  io_wgt_rd_0_data_bits_29_6,
  input  [7:0]  io_wgt_rd_0_data_bits_29_7,
  input  [7:0]  io_wgt_rd_0_data_bits_29_8,
  input  [7:0]  io_wgt_rd_0_data_bits_29_9,
  input  [7:0]  io_wgt_rd_0_data_bits_29_10,
  input  [7:0]  io_wgt_rd_0_data_bits_29_11,
  input  [7:0]  io_wgt_rd_0_data_bits_29_12,
  input  [7:0]  io_wgt_rd_0_data_bits_29_13,
  input  [7:0]  io_wgt_rd_0_data_bits_29_14,
  input  [7:0]  io_wgt_rd_0_data_bits_29_15,
  input  [7:0]  io_wgt_rd_0_data_bits_30_0,
  input  [7:0]  io_wgt_rd_0_data_bits_30_1,
  input  [7:0]  io_wgt_rd_0_data_bits_30_2,
  input  [7:0]  io_wgt_rd_0_data_bits_30_3,
  input  [7:0]  io_wgt_rd_0_data_bits_30_4,
  input  [7:0]  io_wgt_rd_0_data_bits_30_5,
  input  [7:0]  io_wgt_rd_0_data_bits_30_6,
  input  [7:0]  io_wgt_rd_0_data_bits_30_7,
  input  [7:0]  io_wgt_rd_0_data_bits_30_8,
  input  [7:0]  io_wgt_rd_0_data_bits_30_9,
  input  [7:0]  io_wgt_rd_0_data_bits_30_10,
  input  [7:0]  io_wgt_rd_0_data_bits_30_11,
  input  [7:0]  io_wgt_rd_0_data_bits_30_12,
  input  [7:0]  io_wgt_rd_0_data_bits_30_13,
  input  [7:0]  io_wgt_rd_0_data_bits_30_14,
  input  [7:0]  io_wgt_rd_0_data_bits_30_15,
  input  [7:0]  io_wgt_rd_0_data_bits_31_0,
  input  [7:0]  io_wgt_rd_0_data_bits_31_1,
  input  [7:0]  io_wgt_rd_0_data_bits_31_2,
  input  [7:0]  io_wgt_rd_0_data_bits_31_3,
  input  [7:0]  io_wgt_rd_0_data_bits_31_4,
  input  [7:0]  io_wgt_rd_0_data_bits_31_5,
  input  [7:0]  io_wgt_rd_0_data_bits_31_6,
  input  [7:0]  io_wgt_rd_0_data_bits_31_7,
  input  [7:0]  io_wgt_rd_0_data_bits_31_8,
  input  [7:0]  io_wgt_rd_0_data_bits_31_9,
  input  [7:0]  io_wgt_rd_0_data_bits_31_10,
  input  [7:0]  io_wgt_rd_0_data_bits_31_11,
  input  [7:0]  io_wgt_rd_0_data_bits_31_12,
  input  [7:0]  io_wgt_rd_0_data_bits_31_13,
  input  [7:0]  io_wgt_rd_0_data_bits_31_14,
  input  [7:0]  io_wgt_rd_0_data_bits_31_15,
  output        io_acc_rd_0_idx_valid,
  output [6:0]  io_acc_rd_0_idx_bits,
  input         io_acc_rd_0_data_valid,
  input  [31:0] io_acc_rd_0_data_bits_0_0,
  input  [31:0] io_acc_rd_0_data_bits_0_1,
  input  [31:0] io_acc_rd_0_data_bits_0_2,
  input  [31:0] io_acc_rd_0_data_bits_0_3,
  input  [31:0] io_acc_rd_0_data_bits_0_4,
  input  [31:0] io_acc_rd_0_data_bits_0_5,
  input  [31:0] io_acc_rd_0_data_bits_0_6,
  input  [31:0] io_acc_rd_0_data_bits_0_7,
  input  [31:0] io_acc_rd_0_data_bits_0_8,
  input  [31:0] io_acc_rd_0_data_bits_0_9,
  input  [31:0] io_acc_rd_0_data_bits_0_10,
  input  [31:0] io_acc_rd_0_data_bits_0_11,
  input  [31:0] io_acc_rd_0_data_bits_0_12,
  input  [31:0] io_acc_rd_0_data_bits_0_13,
  input  [31:0] io_acc_rd_0_data_bits_0_14,
  input  [31:0] io_acc_rd_0_data_bits_0_15,
  input  [31:0] io_acc_rd_0_data_bits_0_16,
  input  [31:0] io_acc_rd_0_data_bits_0_17,
  input  [31:0] io_acc_rd_0_data_bits_0_18,
  input  [31:0] io_acc_rd_0_data_bits_0_19,
  input  [31:0] io_acc_rd_0_data_bits_0_20,
  input  [31:0] io_acc_rd_0_data_bits_0_21,
  input  [31:0] io_acc_rd_0_data_bits_0_22,
  input  [31:0] io_acc_rd_0_data_bits_0_23,
  input  [31:0] io_acc_rd_0_data_bits_0_24,
  input  [31:0] io_acc_rd_0_data_bits_0_25,
  input  [31:0] io_acc_rd_0_data_bits_0_26,
  input  [31:0] io_acc_rd_0_data_bits_0_27,
  input  [31:0] io_acc_rd_0_data_bits_0_28,
  input  [31:0] io_acc_rd_0_data_bits_0_29,
  input  [31:0] io_acc_rd_0_data_bits_0_30,
  input  [31:0] io_acc_rd_0_data_bits_0_31,
  output        io_acc_wr_0_valid,
  output [6:0]  io_acc_wr_0_bits_idx,
  output [31:0] io_acc_wr_0_bits_data_0_0,
  output [31:0] io_acc_wr_0_bits_data_0_1,
  output [31:0] io_acc_wr_0_bits_data_0_2,
  output [31:0] io_acc_wr_0_bits_data_0_3,
  output [31:0] io_acc_wr_0_bits_data_0_4,
  output [31:0] io_acc_wr_0_bits_data_0_5,
  output [31:0] io_acc_wr_0_bits_data_0_6,
  output [31:0] io_acc_wr_0_bits_data_0_7,
  output [31:0] io_acc_wr_0_bits_data_0_8,
  output [31:0] io_acc_wr_0_bits_data_0_9,
  output [31:0] io_acc_wr_0_bits_data_0_10,
  output [31:0] io_acc_wr_0_bits_data_0_11,
  output [31:0] io_acc_wr_0_bits_data_0_12,
  output [31:0] io_acc_wr_0_bits_data_0_13,
  output [31:0] io_acc_wr_0_bits_data_0_14,
  output [31:0] io_acc_wr_0_bits_data_0_15,
  output [31:0] io_acc_wr_0_bits_data_0_16,
  output [31:0] io_acc_wr_0_bits_data_0_17,
  output [31:0] io_acc_wr_0_bits_data_0_18,
  output [31:0] io_acc_wr_0_bits_data_0_19,
  output [31:0] io_acc_wr_0_bits_data_0_20,
  output [31:0] io_acc_wr_0_bits_data_0_21,
  output [31:0] io_acc_wr_0_bits_data_0_22,
  output [31:0] io_acc_wr_0_bits_data_0_23,
  output [31:0] io_acc_wr_0_bits_data_0_24,
  output [31:0] io_acc_wr_0_bits_data_0_25,
  output [31:0] io_acc_wr_0_bits_data_0_26,
  output [31:0] io_acc_wr_0_bits_data_0_27,
  output [31:0] io_acc_wr_0_bits_data_0_28,
  output [31:0] io_acc_wr_0_bits_data_0_29,
  output [31:0] io_acc_wr_0_bits_data_0_30,
  output [31:0] io_acc_wr_0_bits_data_0_31,
  input         io_out_rd_0_data_valid,
  output        io_out_wr_0_valid,
  output [6:0]  io_out_wr_0_bits_idx,
  output [7:0]  io_out_wr_0_bits_data_0_0,
  output [7:0]  io_out_wr_0_bits_data_0_1,
  output [7:0]  io_out_wr_0_bits_data_0_2,
  output [7:0]  io_out_wr_0_bits_data_0_3,
  output [7:0]  io_out_wr_0_bits_data_0_4,
  output [7:0]  io_out_wr_0_bits_data_0_5,
  output [7:0]  io_out_wr_0_bits_data_0_6,
  output [7:0]  io_out_wr_0_bits_data_0_7,
  output [7:0]  io_out_wr_0_bits_data_0_8,
  output [7:0]  io_out_wr_0_bits_data_0_9,
  output [7:0]  io_out_wr_0_bits_data_0_10,
  output [7:0]  io_out_wr_0_bits_data_0_11,
  output [7:0]  io_out_wr_0_bits_data_0_12,
  output [7:0]  io_out_wr_0_bits_data_0_13,
  output [7:0]  io_out_wr_0_bits_data_0_14,
  output [7:0]  io_out_wr_0_bits_data_0_15,
  output [7:0]  io_out_wr_0_bits_data_0_16,
  output [7:0]  io_out_wr_0_bits_data_0_17,
  output [7:0]  io_out_wr_0_bits_data_0_18,
  output [7:0]  io_out_wr_0_bits_data_0_19,
  output [7:0]  io_out_wr_0_bits_data_0_20,
  output [7:0]  io_out_wr_0_bits_data_0_21,
  output [7:0]  io_out_wr_0_bits_data_0_22,
  output [7:0]  io_out_wr_0_bits_data_0_23,
  output [7:0]  io_out_wr_0_bits_data_0_24,
  output [7:0]  io_out_wr_0_bits_data_0_25,
  output [7:0]  io_out_wr_0_bits_data_0_26,
  output [7:0]  io_out_wr_0_bits_data_0_27,
  output [7:0]  io_out_wr_0_bits_data_0_28,
  output [7:0]  io_out_wr_0_bits_data_0_29,
  output [7:0]  io_out_wr_0_bits_data_0_30,
  output [7:0]  io_out_wr_0_bits_data_0_31
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
`endif // RANDOMIZE_REG_INIT
  wire  m_clock; // @[TensorGemm.scala 554:17]
  wire  m_reset; // @[TensorGemm.scala 554:17]
  wire  m_io_start; // @[TensorGemm.scala 554:17]
  wire  m_io_last; // @[TensorGemm.scala 554:17]
  wire [9:0] m_io_dec_wgt_1; // @[TensorGemm.scala 554:17]
  wire [9:0] m_io_dec_wgt_0; // @[TensorGemm.scala 554:17]
  wire [10:0] m_io_dec_inp_1; // @[TensorGemm.scala 554:17]
  wire [10:0] m_io_dec_inp_0; // @[TensorGemm.scala 554:17]
  wire [10:0] m_io_dec_acc_1; // @[TensorGemm.scala 554:17]
  wire [10:0] m_io_dec_acc_0; // @[TensorGemm.scala 554:17]
  wire [13:0] m_io_dec_lp_1; // @[TensorGemm.scala 554:17]
  wire [13:0] m_io_dec_lp_0; // @[TensorGemm.scala 554:17]
  wire [13:0] m_io_dec_uop_end; // @[TensorGemm.scala 554:17]
  wire [12:0] m_io_dec_uop_begin; // @[TensorGemm.scala 554:17]
  wire [6:0] m_io_acc_i; // @[TensorGemm.scala 554:17]
  wire [6:0] m_io_inp_i; // @[TensorGemm.scala 554:17]
  wire [5:0] m_io_wgt_i; // @[TensorGemm.scala 554:17]
  wire [6:0] m_io_uop_idx; // @[TensorGemm.scala 554:17]
  wire  m_io_valid; // @[TensorGemm.scala 554:17]
  wire  reset_pipe_clock; // @[TensorGemm.scala 603:26]
  wire  reset_pipe_reset; // @[TensorGemm.scala 603:26]
  wire  reset_pipe_io_enq_valid; // @[TensorGemm.scala 603:26]
  wire  reset_pipe_io_enq_bits; // @[TensorGemm.scala 603:26]
  wire  reset_pipe_io_deq_valid; // @[TensorGemm.scala 603:26]
  wire  reset_pipe_io_deq_bits; // @[TensorGemm.scala 603:26]
  wire  acc_idx_pipe_clock; // @[TensorGemm.scala 610:28]
  wire  acc_idx_pipe_reset; // @[TensorGemm.scala 610:28]
  wire  acc_idx_pipe_io_enq_valid; // @[TensorGemm.scala 610:28]
  wire [6:0] acc_idx_pipe_io_enq_bits; // @[TensorGemm.scala 610:28]
  wire  acc_idx_pipe_io_deq_valid; // @[TensorGemm.scala 610:28]
  wire [6:0] acc_idx_pipe_io_deq_bits; // @[TensorGemm.scala 610:28]
  wire  wrpipe0_clock; // @[TensorGemm.scala 637:23]
  wire  wrpipe0_reset; // @[TensorGemm.scala 637:23]
  wire  wrpipe0_io_enq_valid; // @[TensorGemm.scala 637:23]
  wire [6:0] wrpipe0_io_enq_bits; // @[TensorGemm.scala 637:23]
  wire  wrpipe0_io_deq_valid; // @[TensorGemm.scala 637:23]
  wire [6:0] wrpipe0_io_deq_bits; // @[TensorGemm.scala 637:23]
  wire  wrpipeNs_clock; // @[TensorGemm.scala 641:24]
  wire  wrpipeNs_reset; // @[TensorGemm.scala 641:24]
  wire  wrpipeNs_io_enq_valid; // @[TensorGemm.scala 641:24]
  wire [6:0] wrpipeNs_io_enq_bits; // @[TensorGemm.scala 641:24]
  wire  wrpipeNs_io_deq_valid; // @[TensorGemm.scala 641:24]
  wire [6:0] wrpipeNs_io_deq_bits; // @[TensorGemm.scala 641:24]
  wire  wrpipe_0_clock; // @[TensorGemm.scala 645:22]
  wire  wrpipe_0_reset; // @[TensorGemm.scala 645:22]
  wire  wrpipe_0_io_enq_valid; // @[TensorGemm.scala 645:22]
  wire [6:0] wrpipe_0_io_enq_bits; // @[TensorGemm.scala 645:22]
  wire  wrpipe_0_io_deq_valid; // @[TensorGemm.scala 645:22]
  wire [6:0] wrpipe_0_io_deq_bits; // @[TensorGemm.scala 645:22]
  wire  mvc_0_clock; // @[TensorGemm.scala 686:55]
  wire  mvc_0_io_valid_reset; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_inp_data_bits_0_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_inp_data_bits_0_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_inp_data_bits_0_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_inp_data_bits_0_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_inp_data_bits_0_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_inp_data_bits_0_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_inp_data_bits_0_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_inp_data_bits_0_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_inp_data_bits_0_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_inp_data_bits_0_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_inp_data_bits_0_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_inp_data_bits_0_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_inp_data_bits_0_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_inp_data_bits_0_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_inp_data_bits_0_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_inp_data_bits_0_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_0_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_0_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_0_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_0_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_0_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_0_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_0_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_0_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_0_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_0_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_0_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_0_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_0_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_0_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_0_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_0_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_1_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_1_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_1_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_1_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_1_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_1_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_1_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_1_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_1_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_1_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_1_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_1_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_1_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_1_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_1_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_1_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_2_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_2_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_2_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_2_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_2_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_2_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_2_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_2_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_2_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_2_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_2_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_2_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_2_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_2_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_2_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_2_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_3_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_3_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_3_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_3_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_3_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_3_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_3_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_3_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_3_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_3_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_3_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_3_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_3_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_3_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_3_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_3_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_4_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_4_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_4_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_4_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_4_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_4_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_4_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_4_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_4_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_4_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_4_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_4_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_4_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_4_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_4_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_4_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_5_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_5_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_5_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_5_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_5_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_5_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_5_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_5_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_5_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_5_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_5_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_5_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_5_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_5_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_5_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_5_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_6_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_6_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_6_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_6_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_6_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_6_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_6_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_6_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_6_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_6_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_6_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_6_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_6_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_6_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_6_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_6_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_7_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_7_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_7_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_7_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_7_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_7_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_7_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_7_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_7_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_7_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_7_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_7_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_7_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_7_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_7_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_7_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_8_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_8_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_8_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_8_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_8_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_8_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_8_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_8_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_8_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_8_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_8_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_8_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_8_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_8_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_8_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_8_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_9_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_9_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_9_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_9_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_9_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_9_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_9_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_9_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_9_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_9_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_9_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_9_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_9_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_9_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_9_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_9_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_10_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_10_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_10_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_10_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_10_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_10_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_10_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_10_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_10_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_10_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_10_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_10_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_10_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_10_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_10_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_10_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_11_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_11_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_11_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_11_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_11_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_11_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_11_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_11_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_11_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_11_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_11_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_11_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_11_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_11_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_11_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_11_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_12_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_12_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_12_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_12_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_12_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_12_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_12_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_12_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_12_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_12_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_12_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_12_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_12_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_12_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_12_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_12_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_13_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_13_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_13_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_13_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_13_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_13_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_13_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_13_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_13_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_13_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_13_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_13_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_13_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_13_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_13_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_13_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_14_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_14_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_14_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_14_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_14_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_14_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_14_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_14_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_14_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_14_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_14_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_14_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_14_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_14_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_14_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_14_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_15_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_15_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_15_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_15_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_15_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_15_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_15_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_15_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_15_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_15_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_15_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_15_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_15_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_15_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_15_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_15_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_16_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_16_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_16_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_16_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_16_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_16_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_16_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_16_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_16_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_16_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_16_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_16_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_16_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_16_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_16_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_16_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_17_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_17_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_17_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_17_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_17_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_17_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_17_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_17_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_17_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_17_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_17_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_17_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_17_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_17_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_17_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_17_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_18_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_18_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_18_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_18_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_18_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_18_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_18_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_18_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_18_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_18_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_18_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_18_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_18_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_18_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_18_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_18_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_19_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_19_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_19_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_19_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_19_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_19_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_19_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_19_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_19_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_19_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_19_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_19_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_19_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_19_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_19_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_19_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_20_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_20_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_20_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_20_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_20_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_20_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_20_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_20_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_20_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_20_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_20_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_20_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_20_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_20_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_20_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_20_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_21_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_21_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_21_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_21_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_21_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_21_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_21_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_21_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_21_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_21_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_21_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_21_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_21_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_21_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_21_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_21_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_22_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_22_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_22_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_22_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_22_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_22_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_22_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_22_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_22_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_22_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_22_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_22_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_22_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_22_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_22_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_22_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_23_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_23_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_23_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_23_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_23_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_23_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_23_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_23_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_23_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_23_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_23_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_23_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_23_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_23_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_23_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_23_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_24_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_24_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_24_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_24_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_24_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_24_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_24_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_24_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_24_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_24_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_24_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_24_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_24_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_24_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_24_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_24_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_25_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_25_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_25_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_25_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_25_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_25_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_25_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_25_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_25_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_25_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_25_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_25_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_25_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_25_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_25_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_25_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_26_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_26_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_26_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_26_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_26_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_26_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_26_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_26_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_26_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_26_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_26_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_26_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_26_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_26_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_26_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_26_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_27_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_27_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_27_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_27_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_27_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_27_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_27_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_27_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_27_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_27_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_27_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_27_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_27_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_27_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_27_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_27_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_28_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_28_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_28_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_28_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_28_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_28_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_28_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_28_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_28_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_28_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_28_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_28_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_28_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_28_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_28_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_28_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_29_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_29_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_29_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_29_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_29_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_29_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_29_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_29_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_29_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_29_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_29_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_29_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_29_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_29_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_29_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_29_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_30_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_30_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_30_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_30_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_30_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_30_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_30_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_30_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_30_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_30_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_30_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_30_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_30_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_30_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_30_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_30_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_31_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_31_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_31_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_31_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_31_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_31_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_31_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_31_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_31_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_31_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_31_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_31_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_31_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_31_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_31_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_wgt_data_bits_31_15; // @[TensorGemm.scala 686:55]
  wire  mvc_0_io_acc_i_data_valid; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_0; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_1; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_2; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_3; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_4; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_5; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_6; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_7; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_8; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_9; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_10; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_11; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_12; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_13; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_14; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_15; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_16; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_17; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_18; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_19; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_20; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_21; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_22; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_23; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_24; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_25; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_26; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_27; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_28; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_29; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_30; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_i_data_bits_0_31; // @[TensorGemm.scala 686:55]
  wire  mvc_0_io_acc_o_data_valid; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_0; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_1; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_2; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_3; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_4; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_5; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_6; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_7; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_8; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_9; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_10; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_11; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_12; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_13; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_14; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_15; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_16; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_17; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_18; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_19; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_20; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_21; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_22; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_23; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_24; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_25; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_26; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_27; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_28; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_29; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_30; // @[TensorGemm.scala 686:55]
  wire [31:0] mvc_0_io_acc_o_data_bits_0_31; // @[TensorGemm.scala 686:55]
  wire  mvc_0_io_out_data_valid; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_0; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_1; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_2; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_3; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_4; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_5; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_6; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_7; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_8; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_9; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_10; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_11; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_12; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_13; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_14; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_15; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_16; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_17; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_18; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_19; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_20; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_21; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_22; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_23; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_24; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_25; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_26; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_27; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_28; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_29; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_30; // @[TensorGemm.scala 686:55]
  wire [7:0] mvc_0_io_out_data_bits_0_31; // @[TensorGemm.scala 686:55]
  wire  mvc_0_io_bypass_cond; // @[TensorGemm.scala 686:55]
  wire  wrpipe2_clock; // @[TensorGemm.scala 691:25]
  wire  wrpipe2_reset; // @[TensorGemm.scala 691:25]
  wire  wrpipe2_io_enq_valid; // @[TensorGemm.scala 691:25]
  wire [6:0] wrpipe2_io_enq_bits; // @[TensorGemm.scala 691:25]
  wire  wrpipe2_io_deq_valid; // @[TensorGemm.scala 691:25]
  wire [6:0] wrpipe2_io_deq_bits; // @[TensorGemm.scala 691:25]
  reg  delayed_valid; // @[Reg.scala 28:20]
  wire  _GEN_0 = m_io_valid; // @[Reg.scala 29:18 28:20 29:22]
  reg [6:0] delayed_acc_i; // @[Reg.scala 16:16]
  reg [6:0] delayed_inp_i; // @[Reg.scala 16:16]
  reg [5:0] delayed_wgt_i; // @[Reg.scala 16:16]
  reg [1:0] state; // @[TensorGemm.scala 566:22]
  reg [3:0] inflight; // @[TensorGemm.scala 567:25]
  reg [9:0] capture_dec_wgt_1; // @[TensorGemm.scala 569:24]
  reg [9:0] capture_dec_wgt_0; // @[TensorGemm.scala 569:24]
  reg [10:0] capture_dec_inp_1; // @[TensorGemm.scala 569:24]
  reg [10:0] capture_dec_inp_0; // @[TensorGemm.scala 569:24]
  reg [10:0] capture_dec_acc_1; // @[TensorGemm.scala 569:24]
  reg [10:0] capture_dec_acc_0; // @[TensorGemm.scala 569:24]
  reg  capture_dec_empty_0; // @[TensorGemm.scala 569:24]
  reg [13:0] capture_dec_lp_1; // @[TensorGemm.scala 569:24]
  reg [13:0] capture_dec_lp_0; // @[TensorGemm.scala 569:24]
  reg [13:0] capture_dec_uop_end; // @[TensorGemm.scala 569:24]
  reg [12:0] capture_dec_uop_begin; // @[TensorGemm.scala 569:24]
  reg  capture_dec_reset; // @[TensorGemm.scala 569:24]
  reg  capture_dec_push_next; // @[TensorGemm.scala 569:24]
  reg  capture_dec_push_prev; // @[TensorGemm.scala 569:24]
  reg  capture_dec_pop_next; // @[TensorGemm.scala 569:24]
  reg  capture_dec_pop_prev; // @[TensorGemm.scala 569:24]
  reg [2:0] capture_dec_op; // @[TensorGemm.scala 569:24]
  wire  _T = state == 2'h0; // @[TensorGemm.scala 572:14]
  wire  _T_5 = inflight == 4'h0; // @[TensorGemm.scala 579:42]
  wire  _T_6 = state == 2'h2 & inflight == 4'h0; // @[TensorGemm.scala 579:30]
  wire  _GEN_7 = state == 2'h1 & m_io_last ? 1'h0 : _T_6; // @[TensorGemm.scala 571:11 577:43]
  wire [34:0] lo = {capture_dec_uop_end,capture_dec_uop_begin,capture_dec_reset,capture_dec_push_next,
    capture_dec_push_prev,capture_dec_pop_next,capture_dec_pop_prev,capture_dec_op}; // @[TensorGemm.scala 585:41]
  wire [127:0] _T_8 = {capture_dec_wgt_1,capture_dec_wgt_0,capture_dec_inp_1,capture_dec_inp_0,capture_dec_acc_1,
    capture_dec_acc_0,capture_dec_empty_0,capture_dec_lp_1,capture_dec_lp_0,lo}; // @[TensorGemm.scala 585:41]
  wire [34:0] lo_1 = {io_dec_uop_end,io_dec_uop_begin,io_dec_reset,io_dec_push_next,io_dec_push_prev,io_dec_pop_next,
    io_dec_pop_prev,io_dec_op}; // @[TensorGemm.scala 585:59]
  wire [127:0] _T_9 = {io_dec_wgt_1,io_dec_wgt_0,io_dec_inp_1,io_dec_inp_0,io_dec_acc_1,io_dec_acc_0,io_dec_empty_0,
    io_dec_lp_1,io_dec_lp_0,lo_1}; // @[TensorGemm.scala 585:59]
  wire  _T_10 = _T_8 == _T_9; // @[TensorGemm.scala 585:48]
  wire  _T_13 = ~reset; // @[TensorGemm.scala 585:9]
  wire [10:0] _GEN_31 = {{4'd0}, delayed_acc_i}; // @[TensorGemm.scala 599:54]
  wire [10:0] uop_acc = io_uop_data_bits_u0 + _GEN_31; // @[TensorGemm.scala 599:54]
  wire [10:0] _GEN_32 = {{4'd0}, delayed_inp_i}; // @[TensorGemm.scala 600:41]
  wire [10:0] uop_inp = io_uop_data_bits_u1 + _GEN_32; // @[TensorGemm.scala 600:41]
  wire [9:0] _GEN_33 = {{4'd0}, delayed_wgt_i}; // @[TensorGemm.scala 601:54]
  wire [9:0] uop_wgt = io_uop_data_bits_u2 + _GEN_33; // @[TensorGemm.scala 601:54]
  reg  delayed_uop_valid; // @[TensorGemm.scala 618:34]
  reg  io_acc_rd_0_idx_valid_REG; // @[TensorGemm.scala 623:40]
  reg [6:0] io_acc_rd_0_idx_bits_REG; // @[TensorGemm.scala 624:39]
  wire  _T_39 = m_io_valid & wrpipeNs_io_deq_valid; // @[TensorGemm.scala 654:19]
  wire [3:0] _inflight_T_1 = inflight + 4'h1; // @[TensorGemm.scala 657:26]
  wire [3:0] _inflight_T_3 = inflight - 4'h1; // @[TensorGemm.scala 660:26]
  wire [3:0] _GEN_27 = wrpipeNs_io_deq_valid ? _inflight_T_3 : inflight; // @[TensorGemm.scala 658:37 660:14 567:25]
  reg  mvc_0_io_valid_reset_REG; // @[TensorGemm.scala 698:40]
  wire  _GEN_34 = ~_T_39; // @[TensorGemm.scala 656:11]
  TensorGemmIndexGenerator m ( // @[TensorGemm.scala 554:17]
    .clock(m_clock),
    .reset(m_reset),
    .io_start(m_io_start),
    .io_last(m_io_last),
    .io_dec_wgt_1(m_io_dec_wgt_1),
    .io_dec_wgt_0(m_io_dec_wgt_0),
    .io_dec_inp_1(m_io_dec_inp_1),
    .io_dec_inp_0(m_io_dec_inp_0),
    .io_dec_acc_1(m_io_dec_acc_1),
    .io_dec_acc_0(m_io_dec_acc_0),
    .io_dec_lp_1(m_io_dec_lp_1),
    .io_dec_lp_0(m_io_dec_lp_0),
    .io_dec_uop_end(m_io_dec_uop_end),
    .io_dec_uop_begin(m_io_dec_uop_begin),
    .io_acc_i(m_io_acc_i),
    .io_inp_i(m_io_inp_i),
    .io_wgt_i(m_io_wgt_i),
    .io_uop_idx(m_io_uop_idx),
    .io_valid(m_io_valid)
  );
  Pipe reset_pipe ( // @[TensorGemm.scala 603:26]
    .clock(reset_pipe_clock),
    .reset(reset_pipe_reset),
    .io_enq_valid(reset_pipe_io_enq_valid),
    .io_enq_bits(reset_pipe_io_enq_bits),
    .io_deq_valid(reset_pipe_io_deq_valid),
    .io_deq_bits(reset_pipe_io_deq_bits)
  );
  Pipe_1 acc_idx_pipe ( // @[TensorGemm.scala 610:28]
    .clock(acc_idx_pipe_clock),
    .reset(acc_idx_pipe_reset),
    .io_enq_valid(acc_idx_pipe_io_enq_valid),
    .io_enq_bits(acc_idx_pipe_io_enq_bits),
    .io_deq_valid(acc_idx_pipe_io_deq_valid),
    .io_deq_bits(acc_idx_pipe_io_deq_bits)
  );
  Pipe_2 wrpipe0 ( // @[TensorGemm.scala 637:23]
    .clock(wrpipe0_clock),
    .reset(wrpipe0_reset),
    .io_enq_valid(wrpipe0_io_enq_valid),
    .io_enq_bits(wrpipe0_io_enq_bits),
    .io_deq_valid(wrpipe0_io_deq_valid),
    .io_deq_bits(wrpipe0_io_deq_bits)
  );
  Pipe_1 wrpipeNs ( // @[TensorGemm.scala 641:24]
    .clock(wrpipeNs_clock),
    .reset(wrpipeNs_reset),
    .io_enq_valid(wrpipeNs_io_enq_valid),
    .io_enq_bits(wrpipeNs_io_enq_bits),
    .io_deq_valid(wrpipeNs_io_deq_valid),
    .io_deq_bits(wrpipeNs_io_deq_bits)
  );
  Pipe_1 wrpipe_0 ( // @[TensorGemm.scala 645:22]
    .clock(wrpipe_0_clock),
    .reset(wrpipe_0_reset),
    .io_enq_valid(wrpipe_0_io_enq_valid),
    .io_enq_bits(wrpipe_0_io_enq_bits),
    .io_deq_valid(wrpipe_0_io_deq_valid),
    .io_deq_bits(wrpipe_0_io_deq_bits)
  );
  MatrixVectorMultiplicationBypass mvc_0 ( // @[TensorGemm.scala 686:55]
    .clock(mvc_0_clock),
    .io_valid_reset(mvc_0_io_valid_reset),
    .io_inp_data_bits_0_0(mvc_0_io_inp_data_bits_0_0),
    .io_inp_data_bits_0_1(mvc_0_io_inp_data_bits_0_1),
    .io_inp_data_bits_0_2(mvc_0_io_inp_data_bits_0_2),
    .io_inp_data_bits_0_3(mvc_0_io_inp_data_bits_0_3),
    .io_inp_data_bits_0_4(mvc_0_io_inp_data_bits_0_4),
    .io_inp_data_bits_0_5(mvc_0_io_inp_data_bits_0_5),
    .io_inp_data_bits_0_6(mvc_0_io_inp_data_bits_0_6),
    .io_inp_data_bits_0_7(mvc_0_io_inp_data_bits_0_7),
    .io_inp_data_bits_0_8(mvc_0_io_inp_data_bits_0_8),
    .io_inp_data_bits_0_9(mvc_0_io_inp_data_bits_0_9),
    .io_inp_data_bits_0_10(mvc_0_io_inp_data_bits_0_10),
    .io_inp_data_bits_0_11(mvc_0_io_inp_data_bits_0_11),
    .io_inp_data_bits_0_12(mvc_0_io_inp_data_bits_0_12),
    .io_inp_data_bits_0_13(mvc_0_io_inp_data_bits_0_13),
    .io_inp_data_bits_0_14(mvc_0_io_inp_data_bits_0_14),
    .io_inp_data_bits_0_15(mvc_0_io_inp_data_bits_0_15),
    .io_wgt_data_bits_0_0(mvc_0_io_wgt_data_bits_0_0),
    .io_wgt_data_bits_0_1(mvc_0_io_wgt_data_bits_0_1),
    .io_wgt_data_bits_0_2(mvc_0_io_wgt_data_bits_0_2),
    .io_wgt_data_bits_0_3(mvc_0_io_wgt_data_bits_0_3),
    .io_wgt_data_bits_0_4(mvc_0_io_wgt_data_bits_0_4),
    .io_wgt_data_bits_0_5(mvc_0_io_wgt_data_bits_0_5),
    .io_wgt_data_bits_0_6(mvc_0_io_wgt_data_bits_0_6),
    .io_wgt_data_bits_0_7(mvc_0_io_wgt_data_bits_0_7),
    .io_wgt_data_bits_0_8(mvc_0_io_wgt_data_bits_0_8),
    .io_wgt_data_bits_0_9(mvc_0_io_wgt_data_bits_0_9),
    .io_wgt_data_bits_0_10(mvc_0_io_wgt_data_bits_0_10),
    .io_wgt_data_bits_0_11(mvc_0_io_wgt_data_bits_0_11),
    .io_wgt_data_bits_0_12(mvc_0_io_wgt_data_bits_0_12),
    .io_wgt_data_bits_0_13(mvc_0_io_wgt_data_bits_0_13),
    .io_wgt_data_bits_0_14(mvc_0_io_wgt_data_bits_0_14),
    .io_wgt_data_bits_0_15(mvc_0_io_wgt_data_bits_0_15),
    .io_wgt_data_bits_1_0(mvc_0_io_wgt_data_bits_1_0),
    .io_wgt_data_bits_1_1(mvc_0_io_wgt_data_bits_1_1),
    .io_wgt_data_bits_1_2(mvc_0_io_wgt_data_bits_1_2),
    .io_wgt_data_bits_1_3(mvc_0_io_wgt_data_bits_1_3),
    .io_wgt_data_bits_1_4(mvc_0_io_wgt_data_bits_1_4),
    .io_wgt_data_bits_1_5(mvc_0_io_wgt_data_bits_1_5),
    .io_wgt_data_bits_1_6(mvc_0_io_wgt_data_bits_1_6),
    .io_wgt_data_bits_1_7(mvc_0_io_wgt_data_bits_1_7),
    .io_wgt_data_bits_1_8(mvc_0_io_wgt_data_bits_1_8),
    .io_wgt_data_bits_1_9(mvc_0_io_wgt_data_bits_1_9),
    .io_wgt_data_bits_1_10(mvc_0_io_wgt_data_bits_1_10),
    .io_wgt_data_bits_1_11(mvc_0_io_wgt_data_bits_1_11),
    .io_wgt_data_bits_1_12(mvc_0_io_wgt_data_bits_1_12),
    .io_wgt_data_bits_1_13(mvc_0_io_wgt_data_bits_1_13),
    .io_wgt_data_bits_1_14(mvc_0_io_wgt_data_bits_1_14),
    .io_wgt_data_bits_1_15(mvc_0_io_wgt_data_bits_1_15),
    .io_wgt_data_bits_2_0(mvc_0_io_wgt_data_bits_2_0),
    .io_wgt_data_bits_2_1(mvc_0_io_wgt_data_bits_2_1),
    .io_wgt_data_bits_2_2(mvc_0_io_wgt_data_bits_2_2),
    .io_wgt_data_bits_2_3(mvc_0_io_wgt_data_bits_2_3),
    .io_wgt_data_bits_2_4(mvc_0_io_wgt_data_bits_2_4),
    .io_wgt_data_bits_2_5(mvc_0_io_wgt_data_bits_2_5),
    .io_wgt_data_bits_2_6(mvc_0_io_wgt_data_bits_2_6),
    .io_wgt_data_bits_2_7(mvc_0_io_wgt_data_bits_2_7),
    .io_wgt_data_bits_2_8(mvc_0_io_wgt_data_bits_2_8),
    .io_wgt_data_bits_2_9(mvc_0_io_wgt_data_bits_2_9),
    .io_wgt_data_bits_2_10(mvc_0_io_wgt_data_bits_2_10),
    .io_wgt_data_bits_2_11(mvc_0_io_wgt_data_bits_2_11),
    .io_wgt_data_bits_2_12(mvc_0_io_wgt_data_bits_2_12),
    .io_wgt_data_bits_2_13(mvc_0_io_wgt_data_bits_2_13),
    .io_wgt_data_bits_2_14(mvc_0_io_wgt_data_bits_2_14),
    .io_wgt_data_bits_2_15(mvc_0_io_wgt_data_bits_2_15),
    .io_wgt_data_bits_3_0(mvc_0_io_wgt_data_bits_3_0),
    .io_wgt_data_bits_3_1(mvc_0_io_wgt_data_bits_3_1),
    .io_wgt_data_bits_3_2(mvc_0_io_wgt_data_bits_3_2),
    .io_wgt_data_bits_3_3(mvc_0_io_wgt_data_bits_3_3),
    .io_wgt_data_bits_3_4(mvc_0_io_wgt_data_bits_3_4),
    .io_wgt_data_bits_3_5(mvc_0_io_wgt_data_bits_3_5),
    .io_wgt_data_bits_3_6(mvc_0_io_wgt_data_bits_3_6),
    .io_wgt_data_bits_3_7(mvc_0_io_wgt_data_bits_3_7),
    .io_wgt_data_bits_3_8(mvc_0_io_wgt_data_bits_3_8),
    .io_wgt_data_bits_3_9(mvc_0_io_wgt_data_bits_3_9),
    .io_wgt_data_bits_3_10(mvc_0_io_wgt_data_bits_3_10),
    .io_wgt_data_bits_3_11(mvc_0_io_wgt_data_bits_3_11),
    .io_wgt_data_bits_3_12(mvc_0_io_wgt_data_bits_3_12),
    .io_wgt_data_bits_3_13(mvc_0_io_wgt_data_bits_3_13),
    .io_wgt_data_bits_3_14(mvc_0_io_wgt_data_bits_3_14),
    .io_wgt_data_bits_3_15(mvc_0_io_wgt_data_bits_3_15),
    .io_wgt_data_bits_4_0(mvc_0_io_wgt_data_bits_4_0),
    .io_wgt_data_bits_4_1(mvc_0_io_wgt_data_bits_4_1),
    .io_wgt_data_bits_4_2(mvc_0_io_wgt_data_bits_4_2),
    .io_wgt_data_bits_4_3(mvc_0_io_wgt_data_bits_4_3),
    .io_wgt_data_bits_4_4(mvc_0_io_wgt_data_bits_4_4),
    .io_wgt_data_bits_4_5(mvc_0_io_wgt_data_bits_4_5),
    .io_wgt_data_bits_4_6(mvc_0_io_wgt_data_bits_4_6),
    .io_wgt_data_bits_4_7(mvc_0_io_wgt_data_bits_4_7),
    .io_wgt_data_bits_4_8(mvc_0_io_wgt_data_bits_4_8),
    .io_wgt_data_bits_4_9(mvc_0_io_wgt_data_bits_4_9),
    .io_wgt_data_bits_4_10(mvc_0_io_wgt_data_bits_4_10),
    .io_wgt_data_bits_4_11(mvc_0_io_wgt_data_bits_4_11),
    .io_wgt_data_bits_4_12(mvc_0_io_wgt_data_bits_4_12),
    .io_wgt_data_bits_4_13(mvc_0_io_wgt_data_bits_4_13),
    .io_wgt_data_bits_4_14(mvc_0_io_wgt_data_bits_4_14),
    .io_wgt_data_bits_4_15(mvc_0_io_wgt_data_bits_4_15),
    .io_wgt_data_bits_5_0(mvc_0_io_wgt_data_bits_5_0),
    .io_wgt_data_bits_5_1(mvc_0_io_wgt_data_bits_5_1),
    .io_wgt_data_bits_5_2(mvc_0_io_wgt_data_bits_5_2),
    .io_wgt_data_bits_5_3(mvc_0_io_wgt_data_bits_5_3),
    .io_wgt_data_bits_5_4(mvc_0_io_wgt_data_bits_5_4),
    .io_wgt_data_bits_5_5(mvc_0_io_wgt_data_bits_5_5),
    .io_wgt_data_bits_5_6(mvc_0_io_wgt_data_bits_5_6),
    .io_wgt_data_bits_5_7(mvc_0_io_wgt_data_bits_5_7),
    .io_wgt_data_bits_5_8(mvc_0_io_wgt_data_bits_5_8),
    .io_wgt_data_bits_5_9(mvc_0_io_wgt_data_bits_5_9),
    .io_wgt_data_bits_5_10(mvc_0_io_wgt_data_bits_5_10),
    .io_wgt_data_bits_5_11(mvc_0_io_wgt_data_bits_5_11),
    .io_wgt_data_bits_5_12(mvc_0_io_wgt_data_bits_5_12),
    .io_wgt_data_bits_5_13(mvc_0_io_wgt_data_bits_5_13),
    .io_wgt_data_bits_5_14(mvc_0_io_wgt_data_bits_5_14),
    .io_wgt_data_bits_5_15(mvc_0_io_wgt_data_bits_5_15),
    .io_wgt_data_bits_6_0(mvc_0_io_wgt_data_bits_6_0),
    .io_wgt_data_bits_6_1(mvc_0_io_wgt_data_bits_6_1),
    .io_wgt_data_bits_6_2(mvc_0_io_wgt_data_bits_6_2),
    .io_wgt_data_bits_6_3(mvc_0_io_wgt_data_bits_6_3),
    .io_wgt_data_bits_6_4(mvc_0_io_wgt_data_bits_6_4),
    .io_wgt_data_bits_6_5(mvc_0_io_wgt_data_bits_6_5),
    .io_wgt_data_bits_6_6(mvc_0_io_wgt_data_bits_6_6),
    .io_wgt_data_bits_6_7(mvc_0_io_wgt_data_bits_6_7),
    .io_wgt_data_bits_6_8(mvc_0_io_wgt_data_bits_6_8),
    .io_wgt_data_bits_6_9(mvc_0_io_wgt_data_bits_6_9),
    .io_wgt_data_bits_6_10(mvc_0_io_wgt_data_bits_6_10),
    .io_wgt_data_bits_6_11(mvc_0_io_wgt_data_bits_6_11),
    .io_wgt_data_bits_6_12(mvc_0_io_wgt_data_bits_6_12),
    .io_wgt_data_bits_6_13(mvc_0_io_wgt_data_bits_6_13),
    .io_wgt_data_bits_6_14(mvc_0_io_wgt_data_bits_6_14),
    .io_wgt_data_bits_6_15(mvc_0_io_wgt_data_bits_6_15),
    .io_wgt_data_bits_7_0(mvc_0_io_wgt_data_bits_7_0),
    .io_wgt_data_bits_7_1(mvc_0_io_wgt_data_bits_7_1),
    .io_wgt_data_bits_7_2(mvc_0_io_wgt_data_bits_7_2),
    .io_wgt_data_bits_7_3(mvc_0_io_wgt_data_bits_7_3),
    .io_wgt_data_bits_7_4(mvc_0_io_wgt_data_bits_7_4),
    .io_wgt_data_bits_7_5(mvc_0_io_wgt_data_bits_7_5),
    .io_wgt_data_bits_7_6(mvc_0_io_wgt_data_bits_7_6),
    .io_wgt_data_bits_7_7(mvc_0_io_wgt_data_bits_7_7),
    .io_wgt_data_bits_7_8(mvc_0_io_wgt_data_bits_7_8),
    .io_wgt_data_bits_7_9(mvc_0_io_wgt_data_bits_7_9),
    .io_wgt_data_bits_7_10(mvc_0_io_wgt_data_bits_7_10),
    .io_wgt_data_bits_7_11(mvc_0_io_wgt_data_bits_7_11),
    .io_wgt_data_bits_7_12(mvc_0_io_wgt_data_bits_7_12),
    .io_wgt_data_bits_7_13(mvc_0_io_wgt_data_bits_7_13),
    .io_wgt_data_bits_7_14(mvc_0_io_wgt_data_bits_7_14),
    .io_wgt_data_bits_7_15(mvc_0_io_wgt_data_bits_7_15),
    .io_wgt_data_bits_8_0(mvc_0_io_wgt_data_bits_8_0),
    .io_wgt_data_bits_8_1(mvc_0_io_wgt_data_bits_8_1),
    .io_wgt_data_bits_8_2(mvc_0_io_wgt_data_bits_8_2),
    .io_wgt_data_bits_8_3(mvc_0_io_wgt_data_bits_8_3),
    .io_wgt_data_bits_8_4(mvc_0_io_wgt_data_bits_8_4),
    .io_wgt_data_bits_8_5(mvc_0_io_wgt_data_bits_8_5),
    .io_wgt_data_bits_8_6(mvc_0_io_wgt_data_bits_8_6),
    .io_wgt_data_bits_8_7(mvc_0_io_wgt_data_bits_8_7),
    .io_wgt_data_bits_8_8(mvc_0_io_wgt_data_bits_8_8),
    .io_wgt_data_bits_8_9(mvc_0_io_wgt_data_bits_8_9),
    .io_wgt_data_bits_8_10(mvc_0_io_wgt_data_bits_8_10),
    .io_wgt_data_bits_8_11(mvc_0_io_wgt_data_bits_8_11),
    .io_wgt_data_bits_8_12(mvc_0_io_wgt_data_bits_8_12),
    .io_wgt_data_bits_8_13(mvc_0_io_wgt_data_bits_8_13),
    .io_wgt_data_bits_8_14(mvc_0_io_wgt_data_bits_8_14),
    .io_wgt_data_bits_8_15(mvc_0_io_wgt_data_bits_8_15),
    .io_wgt_data_bits_9_0(mvc_0_io_wgt_data_bits_9_0),
    .io_wgt_data_bits_9_1(mvc_0_io_wgt_data_bits_9_1),
    .io_wgt_data_bits_9_2(mvc_0_io_wgt_data_bits_9_2),
    .io_wgt_data_bits_9_3(mvc_0_io_wgt_data_bits_9_3),
    .io_wgt_data_bits_9_4(mvc_0_io_wgt_data_bits_9_4),
    .io_wgt_data_bits_9_5(mvc_0_io_wgt_data_bits_9_5),
    .io_wgt_data_bits_9_6(mvc_0_io_wgt_data_bits_9_6),
    .io_wgt_data_bits_9_7(mvc_0_io_wgt_data_bits_9_7),
    .io_wgt_data_bits_9_8(mvc_0_io_wgt_data_bits_9_8),
    .io_wgt_data_bits_9_9(mvc_0_io_wgt_data_bits_9_9),
    .io_wgt_data_bits_9_10(mvc_0_io_wgt_data_bits_9_10),
    .io_wgt_data_bits_9_11(mvc_0_io_wgt_data_bits_9_11),
    .io_wgt_data_bits_9_12(mvc_0_io_wgt_data_bits_9_12),
    .io_wgt_data_bits_9_13(mvc_0_io_wgt_data_bits_9_13),
    .io_wgt_data_bits_9_14(mvc_0_io_wgt_data_bits_9_14),
    .io_wgt_data_bits_9_15(mvc_0_io_wgt_data_bits_9_15),
    .io_wgt_data_bits_10_0(mvc_0_io_wgt_data_bits_10_0),
    .io_wgt_data_bits_10_1(mvc_0_io_wgt_data_bits_10_1),
    .io_wgt_data_bits_10_2(mvc_0_io_wgt_data_bits_10_2),
    .io_wgt_data_bits_10_3(mvc_0_io_wgt_data_bits_10_3),
    .io_wgt_data_bits_10_4(mvc_0_io_wgt_data_bits_10_4),
    .io_wgt_data_bits_10_5(mvc_0_io_wgt_data_bits_10_5),
    .io_wgt_data_bits_10_6(mvc_0_io_wgt_data_bits_10_6),
    .io_wgt_data_bits_10_7(mvc_0_io_wgt_data_bits_10_7),
    .io_wgt_data_bits_10_8(mvc_0_io_wgt_data_bits_10_8),
    .io_wgt_data_bits_10_9(mvc_0_io_wgt_data_bits_10_9),
    .io_wgt_data_bits_10_10(mvc_0_io_wgt_data_bits_10_10),
    .io_wgt_data_bits_10_11(mvc_0_io_wgt_data_bits_10_11),
    .io_wgt_data_bits_10_12(mvc_0_io_wgt_data_bits_10_12),
    .io_wgt_data_bits_10_13(mvc_0_io_wgt_data_bits_10_13),
    .io_wgt_data_bits_10_14(mvc_0_io_wgt_data_bits_10_14),
    .io_wgt_data_bits_10_15(mvc_0_io_wgt_data_bits_10_15),
    .io_wgt_data_bits_11_0(mvc_0_io_wgt_data_bits_11_0),
    .io_wgt_data_bits_11_1(mvc_0_io_wgt_data_bits_11_1),
    .io_wgt_data_bits_11_2(mvc_0_io_wgt_data_bits_11_2),
    .io_wgt_data_bits_11_3(mvc_0_io_wgt_data_bits_11_3),
    .io_wgt_data_bits_11_4(mvc_0_io_wgt_data_bits_11_4),
    .io_wgt_data_bits_11_5(mvc_0_io_wgt_data_bits_11_5),
    .io_wgt_data_bits_11_6(mvc_0_io_wgt_data_bits_11_6),
    .io_wgt_data_bits_11_7(mvc_0_io_wgt_data_bits_11_7),
    .io_wgt_data_bits_11_8(mvc_0_io_wgt_data_bits_11_8),
    .io_wgt_data_bits_11_9(mvc_0_io_wgt_data_bits_11_9),
    .io_wgt_data_bits_11_10(mvc_0_io_wgt_data_bits_11_10),
    .io_wgt_data_bits_11_11(mvc_0_io_wgt_data_bits_11_11),
    .io_wgt_data_bits_11_12(mvc_0_io_wgt_data_bits_11_12),
    .io_wgt_data_bits_11_13(mvc_0_io_wgt_data_bits_11_13),
    .io_wgt_data_bits_11_14(mvc_0_io_wgt_data_bits_11_14),
    .io_wgt_data_bits_11_15(mvc_0_io_wgt_data_bits_11_15),
    .io_wgt_data_bits_12_0(mvc_0_io_wgt_data_bits_12_0),
    .io_wgt_data_bits_12_1(mvc_0_io_wgt_data_bits_12_1),
    .io_wgt_data_bits_12_2(mvc_0_io_wgt_data_bits_12_2),
    .io_wgt_data_bits_12_3(mvc_0_io_wgt_data_bits_12_3),
    .io_wgt_data_bits_12_4(mvc_0_io_wgt_data_bits_12_4),
    .io_wgt_data_bits_12_5(mvc_0_io_wgt_data_bits_12_5),
    .io_wgt_data_bits_12_6(mvc_0_io_wgt_data_bits_12_6),
    .io_wgt_data_bits_12_7(mvc_0_io_wgt_data_bits_12_7),
    .io_wgt_data_bits_12_8(mvc_0_io_wgt_data_bits_12_8),
    .io_wgt_data_bits_12_9(mvc_0_io_wgt_data_bits_12_9),
    .io_wgt_data_bits_12_10(mvc_0_io_wgt_data_bits_12_10),
    .io_wgt_data_bits_12_11(mvc_0_io_wgt_data_bits_12_11),
    .io_wgt_data_bits_12_12(mvc_0_io_wgt_data_bits_12_12),
    .io_wgt_data_bits_12_13(mvc_0_io_wgt_data_bits_12_13),
    .io_wgt_data_bits_12_14(mvc_0_io_wgt_data_bits_12_14),
    .io_wgt_data_bits_12_15(mvc_0_io_wgt_data_bits_12_15),
    .io_wgt_data_bits_13_0(mvc_0_io_wgt_data_bits_13_0),
    .io_wgt_data_bits_13_1(mvc_0_io_wgt_data_bits_13_1),
    .io_wgt_data_bits_13_2(mvc_0_io_wgt_data_bits_13_2),
    .io_wgt_data_bits_13_3(mvc_0_io_wgt_data_bits_13_3),
    .io_wgt_data_bits_13_4(mvc_0_io_wgt_data_bits_13_4),
    .io_wgt_data_bits_13_5(mvc_0_io_wgt_data_bits_13_5),
    .io_wgt_data_bits_13_6(mvc_0_io_wgt_data_bits_13_6),
    .io_wgt_data_bits_13_7(mvc_0_io_wgt_data_bits_13_7),
    .io_wgt_data_bits_13_8(mvc_0_io_wgt_data_bits_13_8),
    .io_wgt_data_bits_13_9(mvc_0_io_wgt_data_bits_13_9),
    .io_wgt_data_bits_13_10(mvc_0_io_wgt_data_bits_13_10),
    .io_wgt_data_bits_13_11(mvc_0_io_wgt_data_bits_13_11),
    .io_wgt_data_bits_13_12(mvc_0_io_wgt_data_bits_13_12),
    .io_wgt_data_bits_13_13(mvc_0_io_wgt_data_bits_13_13),
    .io_wgt_data_bits_13_14(mvc_0_io_wgt_data_bits_13_14),
    .io_wgt_data_bits_13_15(mvc_0_io_wgt_data_bits_13_15),
    .io_wgt_data_bits_14_0(mvc_0_io_wgt_data_bits_14_0),
    .io_wgt_data_bits_14_1(mvc_0_io_wgt_data_bits_14_1),
    .io_wgt_data_bits_14_2(mvc_0_io_wgt_data_bits_14_2),
    .io_wgt_data_bits_14_3(mvc_0_io_wgt_data_bits_14_3),
    .io_wgt_data_bits_14_4(mvc_0_io_wgt_data_bits_14_4),
    .io_wgt_data_bits_14_5(mvc_0_io_wgt_data_bits_14_5),
    .io_wgt_data_bits_14_6(mvc_0_io_wgt_data_bits_14_6),
    .io_wgt_data_bits_14_7(mvc_0_io_wgt_data_bits_14_7),
    .io_wgt_data_bits_14_8(mvc_0_io_wgt_data_bits_14_8),
    .io_wgt_data_bits_14_9(mvc_0_io_wgt_data_bits_14_9),
    .io_wgt_data_bits_14_10(mvc_0_io_wgt_data_bits_14_10),
    .io_wgt_data_bits_14_11(mvc_0_io_wgt_data_bits_14_11),
    .io_wgt_data_bits_14_12(mvc_0_io_wgt_data_bits_14_12),
    .io_wgt_data_bits_14_13(mvc_0_io_wgt_data_bits_14_13),
    .io_wgt_data_bits_14_14(mvc_0_io_wgt_data_bits_14_14),
    .io_wgt_data_bits_14_15(mvc_0_io_wgt_data_bits_14_15),
    .io_wgt_data_bits_15_0(mvc_0_io_wgt_data_bits_15_0),
    .io_wgt_data_bits_15_1(mvc_0_io_wgt_data_bits_15_1),
    .io_wgt_data_bits_15_2(mvc_0_io_wgt_data_bits_15_2),
    .io_wgt_data_bits_15_3(mvc_0_io_wgt_data_bits_15_3),
    .io_wgt_data_bits_15_4(mvc_0_io_wgt_data_bits_15_4),
    .io_wgt_data_bits_15_5(mvc_0_io_wgt_data_bits_15_5),
    .io_wgt_data_bits_15_6(mvc_0_io_wgt_data_bits_15_6),
    .io_wgt_data_bits_15_7(mvc_0_io_wgt_data_bits_15_7),
    .io_wgt_data_bits_15_8(mvc_0_io_wgt_data_bits_15_8),
    .io_wgt_data_bits_15_9(mvc_0_io_wgt_data_bits_15_9),
    .io_wgt_data_bits_15_10(mvc_0_io_wgt_data_bits_15_10),
    .io_wgt_data_bits_15_11(mvc_0_io_wgt_data_bits_15_11),
    .io_wgt_data_bits_15_12(mvc_0_io_wgt_data_bits_15_12),
    .io_wgt_data_bits_15_13(mvc_0_io_wgt_data_bits_15_13),
    .io_wgt_data_bits_15_14(mvc_0_io_wgt_data_bits_15_14),
    .io_wgt_data_bits_15_15(mvc_0_io_wgt_data_bits_15_15),
    .io_wgt_data_bits_16_0(mvc_0_io_wgt_data_bits_16_0),
    .io_wgt_data_bits_16_1(mvc_0_io_wgt_data_bits_16_1),
    .io_wgt_data_bits_16_2(mvc_0_io_wgt_data_bits_16_2),
    .io_wgt_data_bits_16_3(mvc_0_io_wgt_data_bits_16_3),
    .io_wgt_data_bits_16_4(mvc_0_io_wgt_data_bits_16_4),
    .io_wgt_data_bits_16_5(mvc_0_io_wgt_data_bits_16_5),
    .io_wgt_data_bits_16_6(mvc_0_io_wgt_data_bits_16_6),
    .io_wgt_data_bits_16_7(mvc_0_io_wgt_data_bits_16_7),
    .io_wgt_data_bits_16_8(mvc_0_io_wgt_data_bits_16_8),
    .io_wgt_data_bits_16_9(mvc_0_io_wgt_data_bits_16_9),
    .io_wgt_data_bits_16_10(mvc_0_io_wgt_data_bits_16_10),
    .io_wgt_data_bits_16_11(mvc_0_io_wgt_data_bits_16_11),
    .io_wgt_data_bits_16_12(mvc_0_io_wgt_data_bits_16_12),
    .io_wgt_data_bits_16_13(mvc_0_io_wgt_data_bits_16_13),
    .io_wgt_data_bits_16_14(mvc_0_io_wgt_data_bits_16_14),
    .io_wgt_data_bits_16_15(mvc_0_io_wgt_data_bits_16_15),
    .io_wgt_data_bits_17_0(mvc_0_io_wgt_data_bits_17_0),
    .io_wgt_data_bits_17_1(mvc_0_io_wgt_data_bits_17_1),
    .io_wgt_data_bits_17_2(mvc_0_io_wgt_data_bits_17_2),
    .io_wgt_data_bits_17_3(mvc_0_io_wgt_data_bits_17_3),
    .io_wgt_data_bits_17_4(mvc_0_io_wgt_data_bits_17_4),
    .io_wgt_data_bits_17_5(mvc_0_io_wgt_data_bits_17_5),
    .io_wgt_data_bits_17_6(mvc_0_io_wgt_data_bits_17_6),
    .io_wgt_data_bits_17_7(mvc_0_io_wgt_data_bits_17_7),
    .io_wgt_data_bits_17_8(mvc_0_io_wgt_data_bits_17_8),
    .io_wgt_data_bits_17_9(mvc_0_io_wgt_data_bits_17_9),
    .io_wgt_data_bits_17_10(mvc_0_io_wgt_data_bits_17_10),
    .io_wgt_data_bits_17_11(mvc_0_io_wgt_data_bits_17_11),
    .io_wgt_data_bits_17_12(mvc_0_io_wgt_data_bits_17_12),
    .io_wgt_data_bits_17_13(mvc_0_io_wgt_data_bits_17_13),
    .io_wgt_data_bits_17_14(mvc_0_io_wgt_data_bits_17_14),
    .io_wgt_data_bits_17_15(mvc_0_io_wgt_data_bits_17_15),
    .io_wgt_data_bits_18_0(mvc_0_io_wgt_data_bits_18_0),
    .io_wgt_data_bits_18_1(mvc_0_io_wgt_data_bits_18_1),
    .io_wgt_data_bits_18_2(mvc_0_io_wgt_data_bits_18_2),
    .io_wgt_data_bits_18_3(mvc_0_io_wgt_data_bits_18_3),
    .io_wgt_data_bits_18_4(mvc_0_io_wgt_data_bits_18_4),
    .io_wgt_data_bits_18_5(mvc_0_io_wgt_data_bits_18_5),
    .io_wgt_data_bits_18_6(mvc_0_io_wgt_data_bits_18_6),
    .io_wgt_data_bits_18_7(mvc_0_io_wgt_data_bits_18_7),
    .io_wgt_data_bits_18_8(mvc_0_io_wgt_data_bits_18_8),
    .io_wgt_data_bits_18_9(mvc_0_io_wgt_data_bits_18_9),
    .io_wgt_data_bits_18_10(mvc_0_io_wgt_data_bits_18_10),
    .io_wgt_data_bits_18_11(mvc_0_io_wgt_data_bits_18_11),
    .io_wgt_data_bits_18_12(mvc_0_io_wgt_data_bits_18_12),
    .io_wgt_data_bits_18_13(mvc_0_io_wgt_data_bits_18_13),
    .io_wgt_data_bits_18_14(mvc_0_io_wgt_data_bits_18_14),
    .io_wgt_data_bits_18_15(mvc_0_io_wgt_data_bits_18_15),
    .io_wgt_data_bits_19_0(mvc_0_io_wgt_data_bits_19_0),
    .io_wgt_data_bits_19_1(mvc_0_io_wgt_data_bits_19_1),
    .io_wgt_data_bits_19_2(mvc_0_io_wgt_data_bits_19_2),
    .io_wgt_data_bits_19_3(mvc_0_io_wgt_data_bits_19_3),
    .io_wgt_data_bits_19_4(mvc_0_io_wgt_data_bits_19_4),
    .io_wgt_data_bits_19_5(mvc_0_io_wgt_data_bits_19_5),
    .io_wgt_data_bits_19_6(mvc_0_io_wgt_data_bits_19_6),
    .io_wgt_data_bits_19_7(mvc_0_io_wgt_data_bits_19_7),
    .io_wgt_data_bits_19_8(mvc_0_io_wgt_data_bits_19_8),
    .io_wgt_data_bits_19_9(mvc_0_io_wgt_data_bits_19_9),
    .io_wgt_data_bits_19_10(mvc_0_io_wgt_data_bits_19_10),
    .io_wgt_data_bits_19_11(mvc_0_io_wgt_data_bits_19_11),
    .io_wgt_data_bits_19_12(mvc_0_io_wgt_data_bits_19_12),
    .io_wgt_data_bits_19_13(mvc_0_io_wgt_data_bits_19_13),
    .io_wgt_data_bits_19_14(mvc_0_io_wgt_data_bits_19_14),
    .io_wgt_data_bits_19_15(mvc_0_io_wgt_data_bits_19_15),
    .io_wgt_data_bits_20_0(mvc_0_io_wgt_data_bits_20_0),
    .io_wgt_data_bits_20_1(mvc_0_io_wgt_data_bits_20_1),
    .io_wgt_data_bits_20_2(mvc_0_io_wgt_data_bits_20_2),
    .io_wgt_data_bits_20_3(mvc_0_io_wgt_data_bits_20_3),
    .io_wgt_data_bits_20_4(mvc_0_io_wgt_data_bits_20_4),
    .io_wgt_data_bits_20_5(mvc_0_io_wgt_data_bits_20_5),
    .io_wgt_data_bits_20_6(mvc_0_io_wgt_data_bits_20_6),
    .io_wgt_data_bits_20_7(mvc_0_io_wgt_data_bits_20_7),
    .io_wgt_data_bits_20_8(mvc_0_io_wgt_data_bits_20_8),
    .io_wgt_data_bits_20_9(mvc_0_io_wgt_data_bits_20_9),
    .io_wgt_data_bits_20_10(mvc_0_io_wgt_data_bits_20_10),
    .io_wgt_data_bits_20_11(mvc_0_io_wgt_data_bits_20_11),
    .io_wgt_data_bits_20_12(mvc_0_io_wgt_data_bits_20_12),
    .io_wgt_data_bits_20_13(mvc_0_io_wgt_data_bits_20_13),
    .io_wgt_data_bits_20_14(mvc_0_io_wgt_data_bits_20_14),
    .io_wgt_data_bits_20_15(mvc_0_io_wgt_data_bits_20_15),
    .io_wgt_data_bits_21_0(mvc_0_io_wgt_data_bits_21_0),
    .io_wgt_data_bits_21_1(mvc_0_io_wgt_data_bits_21_1),
    .io_wgt_data_bits_21_2(mvc_0_io_wgt_data_bits_21_2),
    .io_wgt_data_bits_21_3(mvc_0_io_wgt_data_bits_21_3),
    .io_wgt_data_bits_21_4(mvc_0_io_wgt_data_bits_21_4),
    .io_wgt_data_bits_21_5(mvc_0_io_wgt_data_bits_21_5),
    .io_wgt_data_bits_21_6(mvc_0_io_wgt_data_bits_21_6),
    .io_wgt_data_bits_21_7(mvc_0_io_wgt_data_bits_21_7),
    .io_wgt_data_bits_21_8(mvc_0_io_wgt_data_bits_21_8),
    .io_wgt_data_bits_21_9(mvc_0_io_wgt_data_bits_21_9),
    .io_wgt_data_bits_21_10(mvc_0_io_wgt_data_bits_21_10),
    .io_wgt_data_bits_21_11(mvc_0_io_wgt_data_bits_21_11),
    .io_wgt_data_bits_21_12(mvc_0_io_wgt_data_bits_21_12),
    .io_wgt_data_bits_21_13(mvc_0_io_wgt_data_bits_21_13),
    .io_wgt_data_bits_21_14(mvc_0_io_wgt_data_bits_21_14),
    .io_wgt_data_bits_21_15(mvc_0_io_wgt_data_bits_21_15),
    .io_wgt_data_bits_22_0(mvc_0_io_wgt_data_bits_22_0),
    .io_wgt_data_bits_22_1(mvc_0_io_wgt_data_bits_22_1),
    .io_wgt_data_bits_22_2(mvc_0_io_wgt_data_bits_22_2),
    .io_wgt_data_bits_22_3(mvc_0_io_wgt_data_bits_22_3),
    .io_wgt_data_bits_22_4(mvc_0_io_wgt_data_bits_22_4),
    .io_wgt_data_bits_22_5(mvc_0_io_wgt_data_bits_22_5),
    .io_wgt_data_bits_22_6(mvc_0_io_wgt_data_bits_22_6),
    .io_wgt_data_bits_22_7(mvc_0_io_wgt_data_bits_22_7),
    .io_wgt_data_bits_22_8(mvc_0_io_wgt_data_bits_22_8),
    .io_wgt_data_bits_22_9(mvc_0_io_wgt_data_bits_22_9),
    .io_wgt_data_bits_22_10(mvc_0_io_wgt_data_bits_22_10),
    .io_wgt_data_bits_22_11(mvc_0_io_wgt_data_bits_22_11),
    .io_wgt_data_bits_22_12(mvc_0_io_wgt_data_bits_22_12),
    .io_wgt_data_bits_22_13(mvc_0_io_wgt_data_bits_22_13),
    .io_wgt_data_bits_22_14(mvc_0_io_wgt_data_bits_22_14),
    .io_wgt_data_bits_22_15(mvc_0_io_wgt_data_bits_22_15),
    .io_wgt_data_bits_23_0(mvc_0_io_wgt_data_bits_23_0),
    .io_wgt_data_bits_23_1(mvc_0_io_wgt_data_bits_23_1),
    .io_wgt_data_bits_23_2(mvc_0_io_wgt_data_bits_23_2),
    .io_wgt_data_bits_23_3(mvc_0_io_wgt_data_bits_23_3),
    .io_wgt_data_bits_23_4(mvc_0_io_wgt_data_bits_23_4),
    .io_wgt_data_bits_23_5(mvc_0_io_wgt_data_bits_23_5),
    .io_wgt_data_bits_23_6(mvc_0_io_wgt_data_bits_23_6),
    .io_wgt_data_bits_23_7(mvc_0_io_wgt_data_bits_23_7),
    .io_wgt_data_bits_23_8(mvc_0_io_wgt_data_bits_23_8),
    .io_wgt_data_bits_23_9(mvc_0_io_wgt_data_bits_23_9),
    .io_wgt_data_bits_23_10(mvc_0_io_wgt_data_bits_23_10),
    .io_wgt_data_bits_23_11(mvc_0_io_wgt_data_bits_23_11),
    .io_wgt_data_bits_23_12(mvc_0_io_wgt_data_bits_23_12),
    .io_wgt_data_bits_23_13(mvc_0_io_wgt_data_bits_23_13),
    .io_wgt_data_bits_23_14(mvc_0_io_wgt_data_bits_23_14),
    .io_wgt_data_bits_23_15(mvc_0_io_wgt_data_bits_23_15),
    .io_wgt_data_bits_24_0(mvc_0_io_wgt_data_bits_24_0),
    .io_wgt_data_bits_24_1(mvc_0_io_wgt_data_bits_24_1),
    .io_wgt_data_bits_24_2(mvc_0_io_wgt_data_bits_24_2),
    .io_wgt_data_bits_24_3(mvc_0_io_wgt_data_bits_24_3),
    .io_wgt_data_bits_24_4(mvc_0_io_wgt_data_bits_24_4),
    .io_wgt_data_bits_24_5(mvc_0_io_wgt_data_bits_24_5),
    .io_wgt_data_bits_24_6(mvc_0_io_wgt_data_bits_24_6),
    .io_wgt_data_bits_24_7(mvc_0_io_wgt_data_bits_24_7),
    .io_wgt_data_bits_24_8(mvc_0_io_wgt_data_bits_24_8),
    .io_wgt_data_bits_24_9(mvc_0_io_wgt_data_bits_24_9),
    .io_wgt_data_bits_24_10(mvc_0_io_wgt_data_bits_24_10),
    .io_wgt_data_bits_24_11(mvc_0_io_wgt_data_bits_24_11),
    .io_wgt_data_bits_24_12(mvc_0_io_wgt_data_bits_24_12),
    .io_wgt_data_bits_24_13(mvc_0_io_wgt_data_bits_24_13),
    .io_wgt_data_bits_24_14(mvc_0_io_wgt_data_bits_24_14),
    .io_wgt_data_bits_24_15(mvc_0_io_wgt_data_bits_24_15),
    .io_wgt_data_bits_25_0(mvc_0_io_wgt_data_bits_25_0),
    .io_wgt_data_bits_25_1(mvc_0_io_wgt_data_bits_25_1),
    .io_wgt_data_bits_25_2(mvc_0_io_wgt_data_bits_25_2),
    .io_wgt_data_bits_25_3(mvc_0_io_wgt_data_bits_25_3),
    .io_wgt_data_bits_25_4(mvc_0_io_wgt_data_bits_25_4),
    .io_wgt_data_bits_25_5(mvc_0_io_wgt_data_bits_25_5),
    .io_wgt_data_bits_25_6(mvc_0_io_wgt_data_bits_25_6),
    .io_wgt_data_bits_25_7(mvc_0_io_wgt_data_bits_25_7),
    .io_wgt_data_bits_25_8(mvc_0_io_wgt_data_bits_25_8),
    .io_wgt_data_bits_25_9(mvc_0_io_wgt_data_bits_25_9),
    .io_wgt_data_bits_25_10(mvc_0_io_wgt_data_bits_25_10),
    .io_wgt_data_bits_25_11(mvc_0_io_wgt_data_bits_25_11),
    .io_wgt_data_bits_25_12(mvc_0_io_wgt_data_bits_25_12),
    .io_wgt_data_bits_25_13(mvc_0_io_wgt_data_bits_25_13),
    .io_wgt_data_bits_25_14(mvc_0_io_wgt_data_bits_25_14),
    .io_wgt_data_bits_25_15(mvc_0_io_wgt_data_bits_25_15),
    .io_wgt_data_bits_26_0(mvc_0_io_wgt_data_bits_26_0),
    .io_wgt_data_bits_26_1(mvc_0_io_wgt_data_bits_26_1),
    .io_wgt_data_bits_26_2(mvc_0_io_wgt_data_bits_26_2),
    .io_wgt_data_bits_26_3(mvc_0_io_wgt_data_bits_26_3),
    .io_wgt_data_bits_26_4(mvc_0_io_wgt_data_bits_26_4),
    .io_wgt_data_bits_26_5(mvc_0_io_wgt_data_bits_26_5),
    .io_wgt_data_bits_26_6(mvc_0_io_wgt_data_bits_26_6),
    .io_wgt_data_bits_26_7(mvc_0_io_wgt_data_bits_26_7),
    .io_wgt_data_bits_26_8(mvc_0_io_wgt_data_bits_26_8),
    .io_wgt_data_bits_26_9(mvc_0_io_wgt_data_bits_26_9),
    .io_wgt_data_bits_26_10(mvc_0_io_wgt_data_bits_26_10),
    .io_wgt_data_bits_26_11(mvc_0_io_wgt_data_bits_26_11),
    .io_wgt_data_bits_26_12(mvc_0_io_wgt_data_bits_26_12),
    .io_wgt_data_bits_26_13(mvc_0_io_wgt_data_bits_26_13),
    .io_wgt_data_bits_26_14(mvc_0_io_wgt_data_bits_26_14),
    .io_wgt_data_bits_26_15(mvc_0_io_wgt_data_bits_26_15),
    .io_wgt_data_bits_27_0(mvc_0_io_wgt_data_bits_27_0),
    .io_wgt_data_bits_27_1(mvc_0_io_wgt_data_bits_27_1),
    .io_wgt_data_bits_27_2(mvc_0_io_wgt_data_bits_27_2),
    .io_wgt_data_bits_27_3(mvc_0_io_wgt_data_bits_27_3),
    .io_wgt_data_bits_27_4(mvc_0_io_wgt_data_bits_27_4),
    .io_wgt_data_bits_27_5(mvc_0_io_wgt_data_bits_27_5),
    .io_wgt_data_bits_27_6(mvc_0_io_wgt_data_bits_27_6),
    .io_wgt_data_bits_27_7(mvc_0_io_wgt_data_bits_27_7),
    .io_wgt_data_bits_27_8(mvc_0_io_wgt_data_bits_27_8),
    .io_wgt_data_bits_27_9(mvc_0_io_wgt_data_bits_27_9),
    .io_wgt_data_bits_27_10(mvc_0_io_wgt_data_bits_27_10),
    .io_wgt_data_bits_27_11(mvc_0_io_wgt_data_bits_27_11),
    .io_wgt_data_bits_27_12(mvc_0_io_wgt_data_bits_27_12),
    .io_wgt_data_bits_27_13(mvc_0_io_wgt_data_bits_27_13),
    .io_wgt_data_bits_27_14(mvc_0_io_wgt_data_bits_27_14),
    .io_wgt_data_bits_27_15(mvc_0_io_wgt_data_bits_27_15),
    .io_wgt_data_bits_28_0(mvc_0_io_wgt_data_bits_28_0),
    .io_wgt_data_bits_28_1(mvc_0_io_wgt_data_bits_28_1),
    .io_wgt_data_bits_28_2(mvc_0_io_wgt_data_bits_28_2),
    .io_wgt_data_bits_28_3(mvc_0_io_wgt_data_bits_28_3),
    .io_wgt_data_bits_28_4(mvc_0_io_wgt_data_bits_28_4),
    .io_wgt_data_bits_28_5(mvc_0_io_wgt_data_bits_28_5),
    .io_wgt_data_bits_28_6(mvc_0_io_wgt_data_bits_28_6),
    .io_wgt_data_bits_28_7(mvc_0_io_wgt_data_bits_28_7),
    .io_wgt_data_bits_28_8(mvc_0_io_wgt_data_bits_28_8),
    .io_wgt_data_bits_28_9(mvc_0_io_wgt_data_bits_28_9),
    .io_wgt_data_bits_28_10(mvc_0_io_wgt_data_bits_28_10),
    .io_wgt_data_bits_28_11(mvc_0_io_wgt_data_bits_28_11),
    .io_wgt_data_bits_28_12(mvc_0_io_wgt_data_bits_28_12),
    .io_wgt_data_bits_28_13(mvc_0_io_wgt_data_bits_28_13),
    .io_wgt_data_bits_28_14(mvc_0_io_wgt_data_bits_28_14),
    .io_wgt_data_bits_28_15(mvc_0_io_wgt_data_bits_28_15),
    .io_wgt_data_bits_29_0(mvc_0_io_wgt_data_bits_29_0),
    .io_wgt_data_bits_29_1(mvc_0_io_wgt_data_bits_29_1),
    .io_wgt_data_bits_29_2(mvc_0_io_wgt_data_bits_29_2),
    .io_wgt_data_bits_29_3(mvc_0_io_wgt_data_bits_29_3),
    .io_wgt_data_bits_29_4(mvc_0_io_wgt_data_bits_29_4),
    .io_wgt_data_bits_29_5(mvc_0_io_wgt_data_bits_29_5),
    .io_wgt_data_bits_29_6(mvc_0_io_wgt_data_bits_29_6),
    .io_wgt_data_bits_29_7(mvc_0_io_wgt_data_bits_29_7),
    .io_wgt_data_bits_29_8(mvc_0_io_wgt_data_bits_29_8),
    .io_wgt_data_bits_29_9(mvc_0_io_wgt_data_bits_29_9),
    .io_wgt_data_bits_29_10(mvc_0_io_wgt_data_bits_29_10),
    .io_wgt_data_bits_29_11(mvc_0_io_wgt_data_bits_29_11),
    .io_wgt_data_bits_29_12(mvc_0_io_wgt_data_bits_29_12),
    .io_wgt_data_bits_29_13(mvc_0_io_wgt_data_bits_29_13),
    .io_wgt_data_bits_29_14(mvc_0_io_wgt_data_bits_29_14),
    .io_wgt_data_bits_29_15(mvc_0_io_wgt_data_bits_29_15),
    .io_wgt_data_bits_30_0(mvc_0_io_wgt_data_bits_30_0),
    .io_wgt_data_bits_30_1(mvc_0_io_wgt_data_bits_30_1),
    .io_wgt_data_bits_30_2(mvc_0_io_wgt_data_bits_30_2),
    .io_wgt_data_bits_30_3(mvc_0_io_wgt_data_bits_30_3),
    .io_wgt_data_bits_30_4(mvc_0_io_wgt_data_bits_30_4),
    .io_wgt_data_bits_30_5(mvc_0_io_wgt_data_bits_30_5),
    .io_wgt_data_bits_30_6(mvc_0_io_wgt_data_bits_30_6),
    .io_wgt_data_bits_30_7(mvc_0_io_wgt_data_bits_30_7),
    .io_wgt_data_bits_30_8(mvc_0_io_wgt_data_bits_30_8),
    .io_wgt_data_bits_30_9(mvc_0_io_wgt_data_bits_30_9),
    .io_wgt_data_bits_30_10(mvc_0_io_wgt_data_bits_30_10),
    .io_wgt_data_bits_30_11(mvc_0_io_wgt_data_bits_30_11),
    .io_wgt_data_bits_30_12(mvc_0_io_wgt_data_bits_30_12),
    .io_wgt_data_bits_30_13(mvc_0_io_wgt_data_bits_30_13),
    .io_wgt_data_bits_30_14(mvc_0_io_wgt_data_bits_30_14),
    .io_wgt_data_bits_30_15(mvc_0_io_wgt_data_bits_30_15),
    .io_wgt_data_bits_31_0(mvc_0_io_wgt_data_bits_31_0),
    .io_wgt_data_bits_31_1(mvc_0_io_wgt_data_bits_31_1),
    .io_wgt_data_bits_31_2(mvc_0_io_wgt_data_bits_31_2),
    .io_wgt_data_bits_31_3(mvc_0_io_wgt_data_bits_31_3),
    .io_wgt_data_bits_31_4(mvc_0_io_wgt_data_bits_31_4),
    .io_wgt_data_bits_31_5(mvc_0_io_wgt_data_bits_31_5),
    .io_wgt_data_bits_31_6(mvc_0_io_wgt_data_bits_31_6),
    .io_wgt_data_bits_31_7(mvc_0_io_wgt_data_bits_31_7),
    .io_wgt_data_bits_31_8(mvc_0_io_wgt_data_bits_31_8),
    .io_wgt_data_bits_31_9(mvc_0_io_wgt_data_bits_31_9),
    .io_wgt_data_bits_31_10(mvc_0_io_wgt_data_bits_31_10),
    .io_wgt_data_bits_31_11(mvc_0_io_wgt_data_bits_31_11),
    .io_wgt_data_bits_31_12(mvc_0_io_wgt_data_bits_31_12),
    .io_wgt_data_bits_31_13(mvc_0_io_wgt_data_bits_31_13),
    .io_wgt_data_bits_31_14(mvc_0_io_wgt_data_bits_31_14),
    .io_wgt_data_bits_31_15(mvc_0_io_wgt_data_bits_31_15),
    .io_acc_i_data_valid(mvc_0_io_acc_i_data_valid),
    .io_acc_i_data_bits_0_0(mvc_0_io_acc_i_data_bits_0_0),
    .io_acc_i_data_bits_0_1(mvc_0_io_acc_i_data_bits_0_1),
    .io_acc_i_data_bits_0_2(mvc_0_io_acc_i_data_bits_0_2),
    .io_acc_i_data_bits_0_3(mvc_0_io_acc_i_data_bits_0_3),
    .io_acc_i_data_bits_0_4(mvc_0_io_acc_i_data_bits_0_4),
    .io_acc_i_data_bits_0_5(mvc_0_io_acc_i_data_bits_0_5),
    .io_acc_i_data_bits_0_6(mvc_0_io_acc_i_data_bits_0_6),
    .io_acc_i_data_bits_0_7(mvc_0_io_acc_i_data_bits_0_7),
    .io_acc_i_data_bits_0_8(mvc_0_io_acc_i_data_bits_0_8),
    .io_acc_i_data_bits_0_9(mvc_0_io_acc_i_data_bits_0_9),
    .io_acc_i_data_bits_0_10(mvc_0_io_acc_i_data_bits_0_10),
    .io_acc_i_data_bits_0_11(mvc_0_io_acc_i_data_bits_0_11),
    .io_acc_i_data_bits_0_12(mvc_0_io_acc_i_data_bits_0_12),
    .io_acc_i_data_bits_0_13(mvc_0_io_acc_i_data_bits_0_13),
    .io_acc_i_data_bits_0_14(mvc_0_io_acc_i_data_bits_0_14),
    .io_acc_i_data_bits_0_15(mvc_0_io_acc_i_data_bits_0_15),
    .io_acc_i_data_bits_0_16(mvc_0_io_acc_i_data_bits_0_16),
    .io_acc_i_data_bits_0_17(mvc_0_io_acc_i_data_bits_0_17),
    .io_acc_i_data_bits_0_18(mvc_0_io_acc_i_data_bits_0_18),
    .io_acc_i_data_bits_0_19(mvc_0_io_acc_i_data_bits_0_19),
    .io_acc_i_data_bits_0_20(mvc_0_io_acc_i_data_bits_0_20),
    .io_acc_i_data_bits_0_21(mvc_0_io_acc_i_data_bits_0_21),
    .io_acc_i_data_bits_0_22(mvc_0_io_acc_i_data_bits_0_22),
    .io_acc_i_data_bits_0_23(mvc_0_io_acc_i_data_bits_0_23),
    .io_acc_i_data_bits_0_24(mvc_0_io_acc_i_data_bits_0_24),
    .io_acc_i_data_bits_0_25(mvc_0_io_acc_i_data_bits_0_25),
    .io_acc_i_data_bits_0_26(mvc_0_io_acc_i_data_bits_0_26),
    .io_acc_i_data_bits_0_27(mvc_0_io_acc_i_data_bits_0_27),
    .io_acc_i_data_bits_0_28(mvc_0_io_acc_i_data_bits_0_28),
    .io_acc_i_data_bits_0_29(mvc_0_io_acc_i_data_bits_0_29),
    .io_acc_i_data_bits_0_30(mvc_0_io_acc_i_data_bits_0_30),
    .io_acc_i_data_bits_0_31(mvc_0_io_acc_i_data_bits_0_31),
    .io_acc_o_data_valid(mvc_0_io_acc_o_data_valid),
    .io_acc_o_data_bits_0_0(mvc_0_io_acc_o_data_bits_0_0),
    .io_acc_o_data_bits_0_1(mvc_0_io_acc_o_data_bits_0_1),
    .io_acc_o_data_bits_0_2(mvc_0_io_acc_o_data_bits_0_2),
    .io_acc_o_data_bits_0_3(mvc_0_io_acc_o_data_bits_0_3),
    .io_acc_o_data_bits_0_4(mvc_0_io_acc_o_data_bits_0_4),
    .io_acc_o_data_bits_0_5(mvc_0_io_acc_o_data_bits_0_5),
    .io_acc_o_data_bits_0_6(mvc_0_io_acc_o_data_bits_0_6),
    .io_acc_o_data_bits_0_7(mvc_0_io_acc_o_data_bits_0_7),
    .io_acc_o_data_bits_0_8(mvc_0_io_acc_o_data_bits_0_8),
    .io_acc_o_data_bits_0_9(mvc_0_io_acc_o_data_bits_0_9),
    .io_acc_o_data_bits_0_10(mvc_0_io_acc_o_data_bits_0_10),
    .io_acc_o_data_bits_0_11(mvc_0_io_acc_o_data_bits_0_11),
    .io_acc_o_data_bits_0_12(mvc_0_io_acc_o_data_bits_0_12),
    .io_acc_o_data_bits_0_13(mvc_0_io_acc_o_data_bits_0_13),
    .io_acc_o_data_bits_0_14(mvc_0_io_acc_o_data_bits_0_14),
    .io_acc_o_data_bits_0_15(mvc_0_io_acc_o_data_bits_0_15),
    .io_acc_o_data_bits_0_16(mvc_0_io_acc_o_data_bits_0_16),
    .io_acc_o_data_bits_0_17(mvc_0_io_acc_o_data_bits_0_17),
    .io_acc_o_data_bits_0_18(mvc_0_io_acc_o_data_bits_0_18),
    .io_acc_o_data_bits_0_19(mvc_0_io_acc_o_data_bits_0_19),
    .io_acc_o_data_bits_0_20(mvc_0_io_acc_o_data_bits_0_20),
    .io_acc_o_data_bits_0_21(mvc_0_io_acc_o_data_bits_0_21),
    .io_acc_o_data_bits_0_22(mvc_0_io_acc_o_data_bits_0_22),
    .io_acc_o_data_bits_0_23(mvc_0_io_acc_o_data_bits_0_23),
    .io_acc_o_data_bits_0_24(mvc_0_io_acc_o_data_bits_0_24),
    .io_acc_o_data_bits_0_25(mvc_0_io_acc_o_data_bits_0_25),
    .io_acc_o_data_bits_0_26(mvc_0_io_acc_o_data_bits_0_26),
    .io_acc_o_data_bits_0_27(mvc_0_io_acc_o_data_bits_0_27),
    .io_acc_o_data_bits_0_28(mvc_0_io_acc_o_data_bits_0_28),
    .io_acc_o_data_bits_0_29(mvc_0_io_acc_o_data_bits_0_29),
    .io_acc_o_data_bits_0_30(mvc_0_io_acc_o_data_bits_0_30),
    .io_acc_o_data_bits_0_31(mvc_0_io_acc_o_data_bits_0_31),
    .io_out_data_valid(mvc_0_io_out_data_valid),
    .io_out_data_bits_0_0(mvc_0_io_out_data_bits_0_0),
    .io_out_data_bits_0_1(mvc_0_io_out_data_bits_0_1),
    .io_out_data_bits_0_2(mvc_0_io_out_data_bits_0_2),
    .io_out_data_bits_0_3(mvc_0_io_out_data_bits_0_3),
    .io_out_data_bits_0_4(mvc_0_io_out_data_bits_0_4),
    .io_out_data_bits_0_5(mvc_0_io_out_data_bits_0_5),
    .io_out_data_bits_0_6(mvc_0_io_out_data_bits_0_6),
    .io_out_data_bits_0_7(mvc_0_io_out_data_bits_0_7),
    .io_out_data_bits_0_8(mvc_0_io_out_data_bits_0_8),
    .io_out_data_bits_0_9(mvc_0_io_out_data_bits_0_9),
    .io_out_data_bits_0_10(mvc_0_io_out_data_bits_0_10),
    .io_out_data_bits_0_11(mvc_0_io_out_data_bits_0_11),
    .io_out_data_bits_0_12(mvc_0_io_out_data_bits_0_12),
    .io_out_data_bits_0_13(mvc_0_io_out_data_bits_0_13),
    .io_out_data_bits_0_14(mvc_0_io_out_data_bits_0_14),
    .io_out_data_bits_0_15(mvc_0_io_out_data_bits_0_15),
    .io_out_data_bits_0_16(mvc_0_io_out_data_bits_0_16),
    .io_out_data_bits_0_17(mvc_0_io_out_data_bits_0_17),
    .io_out_data_bits_0_18(mvc_0_io_out_data_bits_0_18),
    .io_out_data_bits_0_19(mvc_0_io_out_data_bits_0_19),
    .io_out_data_bits_0_20(mvc_0_io_out_data_bits_0_20),
    .io_out_data_bits_0_21(mvc_0_io_out_data_bits_0_21),
    .io_out_data_bits_0_22(mvc_0_io_out_data_bits_0_22),
    .io_out_data_bits_0_23(mvc_0_io_out_data_bits_0_23),
    .io_out_data_bits_0_24(mvc_0_io_out_data_bits_0_24),
    .io_out_data_bits_0_25(mvc_0_io_out_data_bits_0_25),
    .io_out_data_bits_0_26(mvc_0_io_out_data_bits_0_26),
    .io_out_data_bits_0_27(mvc_0_io_out_data_bits_0_27),
    .io_out_data_bits_0_28(mvc_0_io_out_data_bits_0_28),
    .io_out_data_bits_0_29(mvc_0_io_out_data_bits_0_29),
    .io_out_data_bits_0_30(mvc_0_io_out_data_bits_0_30),
    .io_out_data_bits_0_31(mvc_0_io_out_data_bits_0_31),
    .io_bypass_cond(mvc_0_io_bypass_cond)
  );
  Pipe_1 wrpipe2 ( // @[TensorGemm.scala 691:25]
    .clock(wrpipe2_clock),
    .reset(wrpipe2_reset),
    .io_enq_valid(wrpipe2_io_enq_valid),
    .io_enq_bits(wrpipe2_io_enq_bits),
    .io_deq_valid(wrpipe2_io_deq_valid),
    .io_deq_bits(wrpipe2_io_deq_bits)
  );
  assign io_done = state == 2'h0 & io_start ? 1'h0 : _GEN_7; // @[TensorGemm.scala 571:11 572:37]
  assign io_uop_idx_valid = m_io_valid; // @[TensorGemm.scala 592:20]
  assign io_uop_idx_bits = m_io_uop_idx; // @[TensorGemm.scala 591:19]
  assign io_inp_rd_0_idx_valid = delayed_valid; // @[TensorGemm.scala 616:26]
  assign io_inp_rd_0_idx_bits = uop_inp[6:0]; // @[TensorGemm.scala 617:25]
  assign io_wgt_rd_0_idx_valid = delayed_valid; // @[TensorGemm.scala 627:30]
  assign io_wgt_rd_0_idx_bits = uop_wgt[5:0]; // @[TensorGemm.scala 628:29]
  assign io_acc_rd_0_idx_valid = io_acc_rd_0_idx_valid_REG; // @[TensorGemm.scala 623:30]
  assign io_acc_rd_0_idx_bits = io_acc_rd_0_idx_bits_REG; // @[TensorGemm.scala 624:29]
  assign io_acc_wr_0_valid = wrpipe_0_io_deq_valid; // @[TensorGemm.scala 723:27]
  assign io_acc_wr_0_bits_idx = wrpipe_0_io_deq_bits; // @[TensorGemm.scala 724:30]
  assign io_acc_wr_0_bits_data_0_0 = mvc_0_io_acc_o_data_bits_0_0; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_1 = mvc_0_io_acc_o_data_bits_0_1; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_2 = mvc_0_io_acc_o_data_bits_0_2; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_3 = mvc_0_io_acc_o_data_bits_0_3; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_4 = mvc_0_io_acc_o_data_bits_0_4; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_5 = mvc_0_io_acc_o_data_bits_0_5; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_6 = mvc_0_io_acc_o_data_bits_0_6; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_7 = mvc_0_io_acc_o_data_bits_0_7; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_8 = mvc_0_io_acc_o_data_bits_0_8; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_9 = mvc_0_io_acc_o_data_bits_0_9; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_10 = mvc_0_io_acc_o_data_bits_0_10; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_11 = mvc_0_io_acc_o_data_bits_0_11; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_12 = mvc_0_io_acc_o_data_bits_0_12; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_13 = mvc_0_io_acc_o_data_bits_0_13; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_14 = mvc_0_io_acc_o_data_bits_0_14; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_15 = mvc_0_io_acc_o_data_bits_0_15; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_16 = mvc_0_io_acc_o_data_bits_0_16; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_17 = mvc_0_io_acc_o_data_bits_0_17; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_18 = mvc_0_io_acc_o_data_bits_0_18; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_19 = mvc_0_io_acc_o_data_bits_0_19; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_20 = mvc_0_io_acc_o_data_bits_0_20; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_21 = mvc_0_io_acc_o_data_bits_0_21; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_22 = mvc_0_io_acc_o_data_bits_0_22; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_23 = mvc_0_io_acc_o_data_bits_0_23; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_24 = mvc_0_io_acc_o_data_bits_0_24; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_25 = mvc_0_io_acc_o_data_bits_0_25; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_26 = mvc_0_io_acc_o_data_bits_0_26; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_27 = mvc_0_io_acc_o_data_bits_0_27; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_28 = mvc_0_io_acc_o_data_bits_0_28; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_29 = mvc_0_io_acc_o_data_bits_0_29; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_30 = mvc_0_io_acc_o_data_bits_0_30; // @[TensorGemm.scala 718:62]
  assign io_acc_wr_0_bits_data_0_31 = mvc_0_io_acc_o_data_bits_0_31; // @[TensorGemm.scala 718:62]
  assign io_out_wr_0_valid = wrpipeNs_io_deq_valid & mvc_0_io_out_data_valid; // @[TensorGemm.scala 742:47]
  assign io_out_wr_0_bits_idx = wrpipeNs_io_deq_bits; // @[TensorGemm.scala 743:25]
  assign io_out_wr_0_bits_data_0_0 = mvc_0_io_out_data_bits_0_0; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_1 = mvc_0_io_out_data_bits_0_1; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_2 = mvc_0_io_out_data_bits_0_2; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_3 = mvc_0_io_out_data_bits_0_3; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_4 = mvc_0_io_out_data_bits_0_4; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_5 = mvc_0_io_out_data_bits_0_5; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_6 = mvc_0_io_out_data_bits_0_6; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_7 = mvc_0_io_out_data_bits_0_7; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_8 = mvc_0_io_out_data_bits_0_8; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_9 = mvc_0_io_out_data_bits_0_9; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_10 = mvc_0_io_out_data_bits_0_10; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_11 = mvc_0_io_out_data_bits_0_11; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_12 = mvc_0_io_out_data_bits_0_12; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_13 = mvc_0_io_out_data_bits_0_13; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_14 = mvc_0_io_out_data_bits_0_14; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_15 = mvc_0_io_out_data_bits_0_15; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_16 = mvc_0_io_out_data_bits_0_16; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_17 = mvc_0_io_out_data_bits_0_17; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_18 = mvc_0_io_out_data_bits_0_18; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_19 = mvc_0_io_out_data_bits_0_19; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_20 = mvc_0_io_out_data_bits_0_20; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_21 = mvc_0_io_out_data_bits_0_21; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_22 = mvc_0_io_out_data_bits_0_22; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_23 = mvc_0_io_out_data_bits_0_23; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_24 = mvc_0_io_out_data_bits_0_24; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_25 = mvc_0_io_out_data_bits_0_25; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_26 = mvc_0_io_out_data_bits_0_26; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_27 = mvc_0_io_out_data_bits_0_27; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_28 = mvc_0_io_out_data_bits_0_28; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_29 = mvc_0_io_out_data_bits_0_29; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_30 = mvc_0_io_out_data_bits_0_30; // @[TensorGemm.scala 733:21 737:63]
  assign io_out_wr_0_bits_data_0_31 = mvc_0_io_out_data_bits_0_31; // @[TensorGemm.scala 733:21 737:63]
  assign m_clock = clock;
  assign m_reset = reset;
  assign m_io_start = io_start; // @[TensorGemm.scala 588:14]
  assign m_io_dec_wgt_1 = io_dec_wgt_1; // @[TensorGemm.scala 590:12]
  assign m_io_dec_wgt_0 = io_dec_wgt_0; // @[TensorGemm.scala 590:12]
  assign m_io_dec_inp_1 = io_dec_inp_1; // @[TensorGemm.scala 590:12]
  assign m_io_dec_inp_0 = io_dec_inp_0; // @[TensorGemm.scala 590:12]
  assign m_io_dec_acc_1 = io_dec_acc_1; // @[TensorGemm.scala 590:12]
  assign m_io_dec_acc_0 = io_dec_acc_0; // @[TensorGemm.scala 590:12]
  assign m_io_dec_lp_1 = io_dec_lp_1; // @[TensorGemm.scala 590:12]
  assign m_io_dec_lp_0 = io_dec_lp_0; // @[TensorGemm.scala 590:12]
  assign m_io_dec_uop_end = io_dec_uop_end; // @[TensorGemm.scala 590:12]
  assign m_io_dec_uop_begin = io_dec_uop_begin; // @[TensorGemm.scala 590:12]
  assign reset_pipe_clock = clock;
  assign reset_pipe_reset = reset;
  assign reset_pipe_io_enq_valid = m_io_valid; // @[TensorGemm.scala 607:27]
  assign reset_pipe_io_enq_bits = capture_dec_reset; // @[TensorGemm.scala 608:26]
  assign acc_idx_pipe_clock = clock;
  assign acc_idx_pipe_reset = reset;
  assign acc_idx_pipe_io_enq_valid = delayed_valid; // @[TensorGemm.scala 612:29]
  assign acc_idx_pipe_io_enq_bits = uop_acc[6:0]; // @[TensorGemm.scala 613:28]
  assign wrpipe0_clock = clock;
  assign wrpipe0_reset = reset;
  assign wrpipe0_io_enq_valid = delayed_valid; // @[TensorGemm.scala 638:24]
  assign wrpipe0_io_enq_bits = uop_acc[6:0]; // @[TensorGemm.scala 639:23]
  assign wrpipeNs_clock = clock;
  assign wrpipeNs_reset = reset;
  assign wrpipeNs_io_enq_valid = wrpipe0_io_deq_valid; // @[TensorGemm.scala 642:19]
  assign wrpipeNs_io_enq_bits = wrpipe0_io_deq_bits; // @[TensorGemm.scala 642:19]
  assign wrpipe_0_clock = clock;
  assign wrpipe_0_reset = reset;
  assign wrpipe_0_io_enq_valid = wrpipe0_io_deq_valid; // @[TensorGemm.scala 646:17]
  assign wrpipe_0_io_enq_bits = wrpipe0_io_deq_bits; // @[TensorGemm.scala 646:17]
  assign mvc_0_clock = clock;
  assign mvc_0_io_valid_reset = mvc_0_io_valid_reset_REG; // @[TensorGemm.scala 698:30]
  assign mvc_0_io_inp_data_bits_0_0 = io_inp_rd_0_data_bits_0_0; // @[TensorGemm.scala 700:27]
  assign mvc_0_io_inp_data_bits_0_1 = io_inp_rd_0_data_bits_0_1; // @[TensorGemm.scala 700:27]
  assign mvc_0_io_inp_data_bits_0_2 = io_inp_rd_0_data_bits_0_2; // @[TensorGemm.scala 700:27]
  assign mvc_0_io_inp_data_bits_0_3 = io_inp_rd_0_data_bits_0_3; // @[TensorGemm.scala 700:27]
  assign mvc_0_io_inp_data_bits_0_4 = io_inp_rd_0_data_bits_0_4; // @[TensorGemm.scala 700:27]
  assign mvc_0_io_inp_data_bits_0_5 = io_inp_rd_0_data_bits_0_5; // @[TensorGemm.scala 700:27]
  assign mvc_0_io_inp_data_bits_0_6 = io_inp_rd_0_data_bits_0_6; // @[TensorGemm.scala 700:27]
  assign mvc_0_io_inp_data_bits_0_7 = io_inp_rd_0_data_bits_0_7; // @[TensorGemm.scala 700:27]
  assign mvc_0_io_inp_data_bits_0_8 = io_inp_rd_0_data_bits_0_8; // @[TensorGemm.scala 700:27]
  assign mvc_0_io_inp_data_bits_0_9 = io_inp_rd_0_data_bits_0_9; // @[TensorGemm.scala 700:27]
  assign mvc_0_io_inp_data_bits_0_10 = io_inp_rd_0_data_bits_0_10; // @[TensorGemm.scala 700:27]
  assign mvc_0_io_inp_data_bits_0_11 = io_inp_rd_0_data_bits_0_11; // @[TensorGemm.scala 700:27]
  assign mvc_0_io_inp_data_bits_0_12 = io_inp_rd_0_data_bits_0_12; // @[TensorGemm.scala 700:27]
  assign mvc_0_io_inp_data_bits_0_13 = io_inp_rd_0_data_bits_0_13; // @[TensorGemm.scala 700:27]
  assign mvc_0_io_inp_data_bits_0_14 = io_inp_rd_0_data_bits_0_14; // @[TensorGemm.scala 700:27]
  assign mvc_0_io_inp_data_bits_0_15 = io_inp_rd_0_data_bits_0_15; // @[TensorGemm.scala 700:27]
  assign mvc_0_io_wgt_data_bits_0_0 = io_wgt_rd_0_data_bits_0_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_0_1 = io_wgt_rd_0_data_bits_0_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_0_2 = io_wgt_rd_0_data_bits_0_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_0_3 = io_wgt_rd_0_data_bits_0_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_0_4 = io_wgt_rd_0_data_bits_0_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_0_5 = io_wgt_rd_0_data_bits_0_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_0_6 = io_wgt_rd_0_data_bits_0_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_0_7 = io_wgt_rd_0_data_bits_0_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_0_8 = io_wgt_rd_0_data_bits_0_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_0_9 = io_wgt_rd_0_data_bits_0_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_0_10 = io_wgt_rd_0_data_bits_0_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_0_11 = io_wgt_rd_0_data_bits_0_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_0_12 = io_wgt_rd_0_data_bits_0_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_0_13 = io_wgt_rd_0_data_bits_0_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_0_14 = io_wgt_rd_0_data_bits_0_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_0_15 = io_wgt_rd_0_data_bits_0_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_1_0 = io_wgt_rd_0_data_bits_1_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_1_1 = io_wgt_rd_0_data_bits_1_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_1_2 = io_wgt_rd_0_data_bits_1_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_1_3 = io_wgt_rd_0_data_bits_1_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_1_4 = io_wgt_rd_0_data_bits_1_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_1_5 = io_wgt_rd_0_data_bits_1_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_1_6 = io_wgt_rd_0_data_bits_1_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_1_7 = io_wgt_rd_0_data_bits_1_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_1_8 = io_wgt_rd_0_data_bits_1_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_1_9 = io_wgt_rd_0_data_bits_1_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_1_10 = io_wgt_rd_0_data_bits_1_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_1_11 = io_wgt_rd_0_data_bits_1_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_1_12 = io_wgt_rd_0_data_bits_1_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_1_13 = io_wgt_rd_0_data_bits_1_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_1_14 = io_wgt_rd_0_data_bits_1_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_1_15 = io_wgt_rd_0_data_bits_1_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_2_0 = io_wgt_rd_0_data_bits_2_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_2_1 = io_wgt_rd_0_data_bits_2_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_2_2 = io_wgt_rd_0_data_bits_2_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_2_3 = io_wgt_rd_0_data_bits_2_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_2_4 = io_wgt_rd_0_data_bits_2_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_2_5 = io_wgt_rd_0_data_bits_2_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_2_6 = io_wgt_rd_0_data_bits_2_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_2_7 = io_wgt_rd_0_data_bits_2_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_2_8 = io_wgt_rd_0_data_bits_2_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_2_9 = io_wgt_rd_0_data_bits_2_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_2_10 = io_wgt_rd_0_data_bits_2_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_2_11 = io_wgt_rd_0_data_bits_2_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_2_12 = io_wgt_rd_0_data_bits_2_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_2_13 = io_wgt_rd_0_data_bits_2_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_2_14 = io_wgt_rd_0_data_bits_2_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_2_15 = io_wgt_rd_0_data_bits_2_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_3_0 = io_wgt_rd_0_data_bits_3_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_3_1 = io_wgt_rd_0_data_bits_3_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_3_2 = io_wgt_rd_0_data_bits_3_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_3_3 = io_wgt_rd_0_data_bits_3_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_3_4 = io_wgt_rd_0_data_bits_3_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_3_5 = io_wgt_rd_0_data_bits_3_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_3_6 = io_wgt_rd_0_data_bits_3_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_3_7 = io_wgt_rd_0_data_bits_3_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_3_8 = io_wgt_rd_0_data_bits_3_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_3_9 = io_wgt_rd_0_data_bits_3_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_3_10 = io_wgt_rd_0_data_bits_3_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_3_11 = io_wgt_rd_0_data_bits_3_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_3_12 = io_wgt_rd_0_data_bits_3_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_3_13 = io_wgt_rd_0_data_bits_3_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_3_14 = io_wgt_rd_0_data_bits_3_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_3_15 = io_wgt_rd_0_data_bits_3_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_4_0 = io_wgt_rd_0_data_bits_4_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_4_1 = io_wgt_rd_0_data_bits_4_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_4_2 = io_wgt_rd_0_data_bits_4_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_4_3 = io_wgt_rd_0_data_bits_4_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_4_4 = io_wgt_rd_0_data_bits_4_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_4_5 = io_wgt_rd_0_data_bits_4_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_4_6 = io_wgt_rd_0_data_bits_4_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_4_7 = io_wgt_rd_0_data_bits_4_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_4_8 = io_wgt_rd_0_data_bits_4_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_4_9 = io_wgt_rd_0_data_bits_4_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_4_10 = io_wgt_rd_0_data_bits_4_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_4_11 = io_wgt_rd_0_data_bits_4_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_4_12 = io_wgt_rd_0_data_bits_4_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_4_13 = io_wgt_rd_0_data_bits_4_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_4_14 = io_wgt_rd_0_data_bits_4_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_4_15 = io_wgt_rd_0_data_bits_4_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_5_0 = io_wgt_rd_0_data_bits_5_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_5_1 = io_wgt_rd_0_data_bits_5_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_5_2 = io_wgt_rd_0_data_bits_5_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_5_3 = io_wgt_rd_0_data_bits_5_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_5_4 = io_wgt_rd_0_data_bits_5_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_5_5 = io_wgt_rd_0_data_bits_5_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_5_6 = io_wgt_rd_0_data_bits_5_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_5_7 = io_wgt_rd_0_data_bits_5_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_5_8 = io_wgt_rd_0_data_bits_5_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_5_9 = io_wgt_rd_0_data_bits_5_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_5_10 = io_wgt_rd_0_data_bits_5_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_5_11 = io_wgt_rd_0_data_bits_5_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_5_12 = io_wgt_rd_0_data_bits_5_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_5_13 = io_wgt_rd_0_data_bits_5_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_5_14 = io_wgt_rd_0_data_bits_5_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_5_15 = io_wgt_rd_0_data_bits_5_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_6_0 = io_wgt_rd_0_data_bits_6_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_6_1 = io_wgt_rd_0_data_bits_6_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_6_2 = io_wgt_rd_0_data_bits_6_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_6_3 = io_wgt_rd_0_data_bits_6_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_6_4 = io_wgt_rd_0_data_bits_6_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_6_5 = io_wgt_rd_0_data_bits_6_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_6_6 = io_wgt_rd_0_data_bits_6_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_6_7 = io_wgt_rd_0_data_bits_6_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_6_8 = io_wgt_rd_0_data_bits_6_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_6_9 = io_wgt_rd_0_data_bits_6_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_6_10 = io_wgt_rd_0_data_bits_6_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_6_11 = io_wgt_rd_0_data_bits_6_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_6_12 = io_wgt_rd_0_data_bits_6_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_6_13 = io_wgt_rd_0_data_bits_6_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_6_14 = io_wgt_rd_0_data_bits_6_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_6_15 = io_wgt_rd_0_data_bits_6_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_7_0 = io_wgt_rd_0_data_bits_7_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_7_1 = io_wgt_rd_0_data_bits_7_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_7_2 = io_wgt_rd_0_data_bits_7_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_7_3 = io_wgt_rd_0_data_bits_7_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_7_4 = io_wgt_rd_0_data_bits_7_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_7_5 = io_wgt_rd_0_data_bits_7_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_7_6 = io_wgt_rd_0_data_bits_7_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_7_7 = io_wgt_rd_0_data_bits_7_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_7_8 = io_wgt_rd_0_data_bits_7_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_7_9 = io_wgt_rd_0_data_bits_7_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_7_10 = io_wgt_rd_0_data_bits_7_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_7_11 = io_wgt_rd_0_data_bits_7_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_7_12 = io_wgt_rd_0_data_bits_7_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_7_13 = io_wgt_rd_0_data_bits_7_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_7_14 = io_wgt_rd_0_data_bits_7_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_7_15 = io_wgt_rd_0_data_bits_7_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_8_0 = io_wgt_rd_0_data_bits_8_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_8_1 = io_wgt_rd_0_data_bits_8_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_8_2 = io_wgt_rd_0_data_bits_8_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_8_3 = io_wgt_rd_0_data_bits_8_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_8_4 = io_wgt_rd_0_data_bits_8_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_8_5 = io_wgt_rd_0_data_bits_8_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_8_6 = io_wgt_rd_0_data_bits_8_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_8_7 = io_wgt_rd_0_data_bits_8_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_8_8 = io_wgt_rd_0_data_bits_8_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_8_9 = io_wgt_rd_0_data_bits_8_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_8_10 = io_wgt_rd_0_data_bits_8_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_8_11 = io_wgt_rd_0_data_bits_8_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_8_12 = io_wgt_rd_0_data_bits_8_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_8_13 = io_wgt_rd_0_data_bits_8_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_8_14 = io_wgt_rd_0_data_bits_8_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_8_15 = io_wgt_rd_0_data_bits_8_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_9_0 = io_wgt_rd_0_data_bits_9_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_9_1 = io_wgt_rd_0_data_bits_9_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_9_2 = io_wgt_rd_0_data_bits_9_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_9_3 = io_wgt_rd_0_data_bits_9_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_9_4 = io_wgt_rd_0_data_bits_9_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_9_5 = io_wgt_rd_0_data_bits_9_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_9_6 = io_wgt_rd_0_data_bits_9_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_9_7 = io_wgt_rd_0_data_bits_9_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_9_8 = io_wgt_rd_0_data_bits_9_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_9_9 = io_wgt_rd_0_data_bits_9_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_9_10 = io_wgt_rd_0_data_bits_9_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_9_11 = io_wgt_rd_0_data_bits_9_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_9_12 = io_wgt_rd_0_data_bits_9_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_9_13 = io_wgt_rd_0_data_bits_9_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_9_14 = io_wgt_rd_0_data_bits_9_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_9_15 = io_wgt_rd_0_data_bits_9_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_10_0 = io_wgt_rd_0_data_bits_10_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_10_1 = io_wgt_rd_0_data_bits_10_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_10_2 = io_wgt_rd_0_data_bits_10_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_10_3 = io_wgt_rd_0_data_bits_10_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_10_4 = io_wgt_rd_0_data_bits_10_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_10_5 = io_wgt_rd_0_data_bits_10_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_10_6 = io_wgt_rd_0_data_bits_10_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_10_7 = io_wgt_rd_0_data_bits_10_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_10_8 = io_wgt_rd_0_data_bits_10_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_10_9 = io_wgt_rd_0_data_bits_10_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_10_10 = io_wgt_rd_0_data_bits_10_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_10_11 = io_wgt_rd_0_data_bits_10_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_10_12 = io_wgt_rd_0_data_bits_10_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_10_13 = io_wgt_rd_0_data_bits_10_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_10_14 = io_wgt_rd_0_data_bits_10_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_10_15 = io_wgt_rd_0_data_bits_10_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_11_0 = io_wgt_rd_0_data_bits_11_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_11_1 = io_wgt_rd_0_data_bits_11_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_11_2 = io_wgt_rd_0_data_bits_11_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_11_3 = io_wgt_rd_0_data_bits_11_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_11_4 = io_wgt_rd_0_data_bits_11_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_11_5 = io_wgt_rd_0_data_bits_11_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_11_6 = io_wgt_rd_0_data_bits_11_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_11_7 = io_wgt_rd_0_data_bits_11_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_11_8 = io_wgt_rd_0_data_bits_11_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_11_9 = io_wgt_rd_0_data_bits_11_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_11_10 = io_wgt_rd_0_data_bits_11_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_11_11 = io_wgt_rd_0_data_bits_11_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_11_12 = io_wgt_rd_0_data_bits_11_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_11_13 = io_wgt_rd_0_data_bits_11_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_11_14 = io_wgt_rd_0_data_bits_11_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_11_15 = io_wgt_rd_0_data_bits_11_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_12_0 = io_wgt_rd_0_data_bits_12_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_12_1 = io_wgt_rd_0_data_bits_12_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_12_2 = io_wgt_rd_0_data_bits_12_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_12_3 = io_wgt_rd_0_data_bits_12_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_12_4 = io_wgt_rd_0_data_bits_12_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_12_5 = io_wgt_rd_0_data_bits_12_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_12_6 = io_wgt_rd_0_data_bits_12_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_12_7 = io_wgt_rd_0_data_bits_12_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_12_8 = io_wgt_rd_0_data_bits_12_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_12_9 = io_wgt_rd_0_data_bits_12_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_12_10 = io_wgt_rd_0_data_bits_12_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_12_11 = io_wgt_rd_0_data_bits_12_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_12_12 = io_wgt_rd_0_data_bits_12_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_12_13 = io_wgt_rd_0_data_bits_12_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_12_14 = io_wgt_rd_0_data_bits_12_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_12_15 = io_wgt_rd_0_data_bits_12_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_13_0 = io_wgt_rd_0_data_bits_13_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_13_1 = io_wgt_rd_0_data_bits_13_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_13_2 = io_wgt_rd_0_data_bits_13_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_13_3 = io_wgt_rd_0_data_bits_13_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_13_4 = io_wgt_rd_0_data_bits_13_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_13_5 = io_wgt_rd_0_data_bits_13_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_13_6 = io_wgt_rd_0_data_bits_13_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_13_7 = io_wgt_rd_0_data_bits_13_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_13_8 = io_wgt_rd_0_data_bits_13_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_13_9 = io_wgt_rd_0_data_bits_13_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_13_10 = io_wgt_rd_0_data_bits_13_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_13_11 = io_wgt_rd_0_data_bits_13_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_13_12 = io_wgt_rd_0_data_bits_13_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_13_13 = io_wgt_rd_0_data_bits_13_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_13_14 = io_wgt_rd_0_data_bits_13_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_13_15 = io_wgt_rd_0_data_bits_13_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_14_0 = io_wgt_rd_0_data_bits_14_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_14_1 = io_wgt_rd_0_data_bits_14_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_14_2 = io_wgt_rd_0_data_bits_14_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_14_3 = io_wgt_rd_0_data_bits_14_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_14_4 = io_wgt_rd_0_data_bits_14_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_14_5 = io_wgt_rd_0_data_bits_14_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_14_6 = io_wgt_rd_0_data_bits_14_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_14_7 = io_wgt_rd_0_data_bits_14_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_14_8 = io_wgt_rd_0_data_bits_14_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_14_9 = io_wgt_rd_0_data_bits_14_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_14_10 = io_wgt_rd_0_data_bits_14_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_14_11 = io_wgt_rd_0_data_bits_14_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_14_12 = io_wgt_rd_0_data_bits_14_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_14_13 = io_wgt_rd_0_data_bits_14_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_14_14 = io_wgt_rd_0_data_bits_14_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_14_15 = io_wgt_rd_0_data_bits_14_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_15_0 = io_wgt_rd_0_data_bits_15_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_15_1 = io_wgt_rd_0_data_bits_15_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_15_2 = io_wgt_rd_0_data_bits_15_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_15_3 = io_wgt_rd_0_data_bits_15_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_15_4 = io_wgt_rd_0_data_bits_15_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_15_5 = io_wgt_rd_0_data_bits_15_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_15_6 = io_wgt_rd_0_data_bits_15_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_15_7 = io_wgt_rd_0_data_bits_15_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_15_8 = io_wgt_rd_0_data_bits_15_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_15_9 = io_wgt_rd_0_data_bits_15_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_15_10 = io_wgt_rd_0_data_bits_15_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_15_11 = io_wgt_rd_0_data_bits_15_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_15_12 = io_wgt_rd_0_data_bits_15_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_15_13 = io_wgt_rd_0_data_bits_15_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_15_14 = io_wgt_rd_0_data_bits_15_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_15_15 = io_wgt_rd_0_data_bits_15_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_16_0 = io_wgt_rd_0_data_bits_16_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_16_1 = io_wgt_rd_0_data_bits_16_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_16_2 = io_wgt_rd_0_data_bits_16_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_16_3 = io_wgt_rd_0_data_bits_16_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_16_4 = io_wgt_rd_0_data_bits_16_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_16_5 = io_wgt_rd_0_data_bits_16_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_16_6 = io_wgt_rd_0_data_bits_16_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_16_7 = io_wgt_rd_0_data_bits_16_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_16_8 = io_wgt_rd_0_data_bits_16_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_16_9 = io_wgt_rd_0_data_bits_16_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_16_10 = io_wgt_rd_0_data_bits_16_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_16_11 = io_wgt_rd_0_data_bits_16_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_16_12 = io_wgt_rd_0_data_bits_16_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_16_13 = io_wgt_rd_0_data_bits_16_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_16_14 = io_wgt_rd_0_data_bits_16_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_16_15 = io_wgt_rd_0_data_bits_16_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_17_0 = io_wgt_rd_0_data_bits_17_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_17_1 = io_wgt_rd_0_data_bits_17_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_17_2 = io_wgt_rd_0_data_bits_17_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_17_3 = io_wgt_rd_0_data_bits_17_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_17_4 = io_wgt_rd_0_data_bits_17_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_17_5 = io_wgt_rd_0_data_bits_17_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_17_6 = io_wgt_rd_0_data_bits_17_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_17_7 = io_wgt_rd_0_data_bits_17_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_17_8 = io_wgt_rd_0_data_bits_17_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_17_9 = io_wgt_rd_0_data_bits_17_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_17_10 = io_wgt_rd_0_data_bits_17_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_17_11 = io_wgt_rd_0_data_bits_17_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_17_12 = io_wgt_rd_0_data_bits_17_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_17_13 = io_wgt_rd_0_data_bits_17_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_17_14 = io_wgt_rd_0_data_bits_17_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_17_15 = io_wgt_rd_0_data_bits_17_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_18_0 = io_wgt_rd_0_data_bits_18_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_18_1 = io_wgt_rd_0_data_bits_18_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_18_2 = io_wgt_rd_0_data_bits_18_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_18_3 = io_wgt_rd_0_data_bits_18_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_18_4 = io_wgt_rd_0_data_bits_18_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_18_5 = io_wgt_rd_0_data_bits_18_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_18_6 = io_wgt_rd_0_data_bits_18_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_18_7 = io_wgt_rd_0_data_bits_18_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_18_8 = io_wgt_rd_0_data_bits_18_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_18_9 = io_wgt_rd_0_data_bits_18_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_18_10 = io_wgt_rd_0_data_bits_18_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_18_11 = io_wgt_rd_0_data_bits_18_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_18_12 = io_wgt_rd_0_data_bits_18_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_18_13 = io_wgt_rd_0_data_bits_18_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_18_14 = io_wgt_rd_0_data_bits_18_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_18_15 = io_wgt_rd_0_data_bits_18_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_19_0 = io_wgt_rd_0_data_bits_19_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_19_1 = io_wgt_rd_0_data_bits_19_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_19_2 = io_wgt_rd_0_data_bits_19_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_19_3 = io_wgt_rd_0_data_bits_19_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_19_4 = io_wgt_rd_0_data_bits_19_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_19_5 = io_wgt_rd_0_data_bits_19_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_19_6 = io_wgt_rd_0_data_bits_19_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_19_7 = io_wgt_rd_0_data_bits_19_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_19_8 = io_wgt_rd_0_data_bits_19_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_19_9 = io_wgt_rd_0_data_bits_19_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_19_10 = io_wgt_rd_0_data_bits_19_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_19_11 = io_wgt_rd_0_data_bits_19_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_19_12 = io_wgt_rd_0_data_bits_19_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_19_13 = io_wgt_rd_0_data_bits_19_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_19_14 = io_wgt_rd_0_data_bits_19_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_19_15 = io_wgt_rd_0_data_bits_19_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_20_0 = io_wgt_rd_0_data_bits_20_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_20_1 = io_wgt_rd_0_data_bits_20_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_20_2 = io_wgt_rd_0_data_bits_20_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_20_3 = io_wgt_rd_0_data_bits_20_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_20_4 = io_wgt_rd_0_data_bits_20_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_20_5 = io_wgt_rd_0_data_bits_20_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_20_6 = io_wgt_rd_0_data_bits_20_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_20_7 = io_wgt_rd_0_data_bits_20_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_20_8 = io_wgt_rd_0_data_bits_20_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_20_9 = io_wgt_rd_0_data_bits_20_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_20_10 = io_wgt_rd_0_data_bits_20_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_20_11 = io_wgt_rd_0_data_bits_20_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_20_12 = io_wgt_rd_0_data_bits_20_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_20_13 = io_wgt_rd_0_data_bits_20_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_20_14 = io_wgt_rd_0_data_bits_20_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_20_15 = io_wgt_rd_0_data_bits_20_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_21_0 = io_wgt_rd_0_data_bits_21_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_21_1 = io_wgt_rd_0_data_bits_21_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_21_2 = io_wgt_rd_0_data_bits_21_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_21_3 = io_wgt_rd_0_data_bits_21_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_21_4 = io_wgt_rd_0_data_bits_21_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_21_5 = io_wgt_rd_0_data_bits_21_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_21_6 = io_wgt_rd_0_data_bits_21_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_21_7 = io_wgt_rd_0_data_bits_21_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_21_8 = io_wgt_rd_0_data_bits_21_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_21_9 = io_wgt_rd_0_data_bits_21_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_21_10 = io_wgt_rd_0_data_bits_21_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_21_11 = io_wgt_rd_0_data_bits_21_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_21_12 = io_wgt_rd_0_data_bits_21_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_21_13 = io_wgt_rd_0_data_bits_21_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_21_14 = io_wgt_rd_0_data_bits_21_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_21_15 = io_wgt_rd_0_data_bits_21_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_22_0 = io_wgt_rd_0_data_bits_22_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_22_1 = io_wgt_rd_0_data_bits_22_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_22_2 = io_wgt_rd_0_data_bits_22_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_22_3 = io_wgt_rd_0_data_bits_22_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_22_4 = io_wgt_rd_0_data_bits_22_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_22_5 = io_wgt_rd_0_data_bits_22_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_22_6 = io_wgt_rd_0_data_bits_22_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_22_7 = io_wgt_rd_0_data_bits_22_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_22_8 = io_wgt_rd_0_data_bits_22_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_22_9 = io_wgt_rd_0_data_bits_22_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_22_10 = io_wgt_rd_0_data_bits_22_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_22_11 = io_wgt_rd_0_data_bits_22_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_22_12 = io_wgt_rd_0_data_bits_22_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_22_13 = io_wgt_rd_0_data_bits_22_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_22_14 = io_wgt_rd_0_data_bits_22_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_22_15 = io_wgt_rd_0_data_bits_22_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_23_0 = io_wgt_rd_0_data_bits_23_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_23_1 = io_wgt_rd_0_data_bits_23_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_23_2 = io_wgt_rd_0_data_bits_23_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_23_3 = io_wgt_rd_0_data_bits_23_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_23_4 = io_wgt_rd_0_data_bits_23_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_23_5 = io_wgt_rd_0_data_bits_23_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_23_6 = io_wgt_rd_0_data_bits_23_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_23_7 = io_wgt_rd_0_data_bits_23_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_23_8 = io_wgt_rd_0_data_bits_23_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_23_9 = io_wgt_rd_0_data_bits_23_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_23_10 = io_wgt_rd_0_data_bits_23_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_23_11 = io_wgt_rd_0_data_bits_23_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_23_12 = io_wgt_rd_0_data_bits_23_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_23_13 = io_wgt_rd_0_data_bits_23_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_23_14 = io_wgt_rd_0_data_bits_23_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_23_15 = io_wgt_rd_0_data_bits_23_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_24_0 = io_wgt_rd_0_data_bits_24_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_24_1 = io_wgt_rd_0_data_bits_24_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_24_2 = io_wgt_rd_0_data_bits_24_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_24_3 = io_wgt_rd_0_data_bits_24_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_24_4 = io_wgt_rd_0_data_bits_24_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_24_5 = io_wgt_rd_0_data_bits_24_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_24_6 = io_wgt_rd_0_data_bits_24_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_24_7 = io_wgt_rd_0_data_bits_24_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_24_8 = io_wgt_rd_0_data_bits_24_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_24_9 = io_wgt_rd_0_data_bits_24_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_24_10 = io_wgt_rd_0_data_bits_24_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_24_11 = io_wgt_rd_0_data_bits_24_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_24_12 = io_wgt_rd_0_data_bits_24_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_24_13 = io_wgt_rd_0_data_bits_24_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_24_14 = io_wgt_rd_0_data_bits_24_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_24_15 = io_wgt_rd_0_data_bits_24_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_25_0 = io_wgt_rd_0_data_bits_25_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_25_1 = io_wgt_rd_0_data_bits_25_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_25_2 = io_wgt_rd_0_data_bits_25_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_25_3 = io_wgt_rd_0_data_bits_25_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_25_4 = io_wgt_rd_0_data_bits_25_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_25_5 = io_wgt_rd_0_data_bits_25_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_25_6 = io_wgt_rd_0_data_bits_25_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_25_7 = io_wgt_rd_0_data_bits_25_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_25_8 = io_wgt_rd_0_data_bits_25_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_25_9 = io_wgt_rd_0_data_bits_25_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_25_10 = io_wgt_rd_0_data_bits_25_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_25_11 = io_wgt_rd_0_data_bits_25_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_25_12 = io_wgt_rd_0_data_bits_25_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_25_13 = io_wgt_rd_0_data_bits_25_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_25_14 = io_wgt_rd_0_data_bits_25_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_25_15 = io_wgt_rd_0_data_bits_25_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_26_0 = io_wgt_rd_0_data_bits_26_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_26_1 = io_wgt_rd_0_data_bits_26_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_26_2 = io_wgt_rd_0_data_bits_26_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_26_3 = io_wgt_rd_0_data_bits_26_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_26_4 = io_wgt_rd_0_data_bits_26_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_26_5 = io_wgt_rd_0_data_bits_26_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_26_6 = io_wgt_rd_0_data_bits_26_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_26_7 = io_wgt_rd_0_data_bits_26_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_26_8 = io_wgt_rd_0_data_bits_26_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_26_9 = io_wgt_rd_0_data_bits_26_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_26_10 = io_wgt_rd_0_data_bits_26_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_26_11 = io_wgt_rd_0_data_bits_26_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_26_12 = io_wgt_rd_0_data_bits_26_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_26_13 = io_wgt_rd_0_data_bits_26_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_26_14 = io_wgt_rd_0_data_bits_26_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_26_15 = io_wgt_rd_0_data_bits_26_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_27_0 = io_wgt_rd_0_data_bits_27_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_27_1 = io_wgt_rd_0_data_bits_27_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_27_2 = io_wgt_rd_0_data_bits_27_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_27_3 = io_wgt_rd_0_data_bits_27_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_27_4 = io_wgt_rd_0_data_bits_27_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_27_5 = io_wgt_rd_0_data_bits_27_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_27_6 = io_wgt_rd_0_data_bits_27_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_27_7 = io_wgt_rd_0_data_bits_27_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_27_8 = io_wgt_rd_0_data_bits_27_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_27_9 = io_wgt_rd_0_data_bits_27_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_27_10 = io_wgt_rd_0_data_bits_27_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_27_11 = io_wgt_rd_0_data_bits_27_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_27_12 = io_wgt_rd_0_data_bits_27_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_27_13 = io_wgt_rd_0_data_bits_27_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_27_14 = io_wgt_rd_0_data_bits_27_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_27_15 = io_wgt_rd_0_data_bits_27_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_28_0 = io_wgt_rd_0_data_bits_28_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_28_1 = io_wgt_rd_0_data_bits_28_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_28_2 = io_wgt_rd_0_data_bits_28_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_28_3 = io_wgt_rd_0_data_bits_28_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_28_4 = io_wgt_rd_0_data_bits_28_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_28_5 = io_wgt_rd_0_data_bits_28_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_28_6 = io_wgt_rd_0_data_bits_28_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_28_7 = io_wgt_rd_0_data_bits_28_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_28_8 = io_wgt_rd_0_data_bits_28_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_28_9 = io_wgt_rd_0_data_bits_28_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_28_10 = io_wgt_rd_0_data_bits_28_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_28_11 = io_wgt_rd_0_data_bits_28_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_28_12 = io_wgt_rd_0_data_bits_28_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_28_13 = io_wgt_rd_0_data_bits_28_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_28_14 = io_wgt_rd_0_data_bits_28_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_28_15 = io_wgt_rd_0_data_bits_28_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_29_0 = io_wgt_rd_0_data_bits_29_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_29_1 = io_wgt_rd_0_data_bits_29_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_29_2 = io_wgt_rd_0_data_bits_29_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_29_3 = io_wgt_rd_0_data_bits_29_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_29_4 = io_wgt_rd_0_data_bits_29_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_29_5 = io_wgt_rd_0_data_bits_29_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_29_6 = io_wgt_rd_0_data_bits_29_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_29_7 = io_wgt_rd_0_data_bits_29_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_29_8 = io_wgt_rd_0_data_bits_29_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_29_9 = io_wgt_rd_0_data_bits_29_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_29_10 = io_wgt_rd_0_data_bits_29_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_29_11 = io_wgt_rd_0_data_bits_29_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_29_12 = io_wgt_rd_0_data_bits_29_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_29_13 = io_wgt_rd_0_data_bits_29_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_29_14 = io_wgt_rd_0_data_bits_29_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_29_15 = io_wgt_rd_0_data_bits_29_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_30_0 = io_wgt_rd_0_data_bits_30_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_30_1 = io_wgt_rd_0_data_bits_30_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_30_2 = io_wgt_rd_0_data_bits_30_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_30_3 = io_wgt_rd_0_data_bits_30_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_30_4 = io_wgt_rd_0_data_bits_30_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_30_5 = io_wgt_rd_0_data_bits_30_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_30_6 = io_wgt_rd_0_data_bits_30_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_30_7 = io_wgt_rd_0_data_bits_30_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_30_8 = io_wgt_rd_0_data_bits_30_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_30_9 = io_wgt_rd_0_data_bits_30_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_30_10 = io_wgt_rd_0_data_bits_30_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_30_11 = io_wgt_rd_0_data_bits_30_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_30_12 = io_wgt_rd_0_data_bits_30_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_30_13 = io_wgt_rd_0_data_bits_30_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_30_14 = io_wgt_rd_0_data_bits_30_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_30_15 = io_wgt_rd_0_data_bits_30_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_31_0 = io_wgt_rd_0_data_bits_31_0; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_31_1 = io_wgt_rd_0_data_bits_31_1; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_31_2 = io_wgt_rd_0_data_bits_31_2; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_31_3 = io_wgt_rd_0_data_bits_31_3; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_31_4 = io_wgt_rd_0_data_bits_31_4; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_31_5 = io_wgt_rd_0_data_bits_31_5; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_31_6 = io_wgt_rd_0_data_bits_31_6; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_31_7 = io_wgt_rd_0_data_bits_31_7; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_31_8 = io_wgt_rd_0_data_bits_31_8; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_31_9 = io_wgt_rd_0_data_bits_31_9; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_31_10 = io_wgt_rd_0_data_bits_31_10; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_31_11 = io_wgt_rd_0_data_bits_31_11; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_31_12 = io_wgt_rd_0_data_bits_31_12; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_31_13 = io_wgt_rd_0_data_bits_31_13; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_31_14 = io_wgt_rd_0_data_bits_31_14; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_wgt_data_bits_31_15 = io_wgt_rd_0_data_bits_31_15; // @[TensorGemm.scala 702:27]
  assign mvc_0_io_acc_i_data_valid = io_acc_rd_0_data_valid; // @[TensorGemm.scala 703:35]
  assign mvc_0_io_acc_i_data_bits_0_0 = io_acc_rd_0_data_bits_0_0; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_1 = io_acc_rd_0_data_bits_0_1; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_2 = io_acc_rd_0_data_bits_0_2; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_3 = io_acc_rd_0_data_bits_0_3; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_4 = io_acc_rd_0_data_bits_0_4; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_5 = io_acc_rd_0_data_bits_0_5; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_6 = io_acc_rd_0_data_bits_0_6; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_7 = io_acc_rd_0_data_bits_0_7; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_8 = io_acc_rd_0_data_bits_0_8; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_9 = io_acc_rd_0_data_bits_0_9; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_10 = io_acc_rd_0_data_bits_0_10; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_11 = io_acc_rd_0_data_bits_0_11; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_12 = io_acc_rd_0_data_bits_0_12; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_13 = io_acc_rd_0_data_bits_0_13; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_14 = io_acc_rd_0_data_bits_0_14; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_15 = io_acc_rd_0_data_bits_0_15; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_16 = io_acc_rd_0_data_bits_0_16; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_17 = io_acc_rd_0_data_bits_0_17; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_18 = io_acc_rd_0_data_bits_0_18; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_19 = io_acc_rd_0_data_bits_0_19; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_20 = io_acc_rd_0_data_bits_0_20; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_21 = io_acc_rd_0_data_bits_0_21; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_22 = io_acc_rd_0_data_bits_0_22; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_23 = io_acc_rd_0_data_bits_0_23; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_24 = io_acc_rd_0_data_bits_0_24; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_25 = io_acc_rd_0_data_bits_0_25; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_26 = io_acc_rd_0_data_bits_0_26; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_27 = io_acc_rd_0_data_bits_0_27; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_28 = io_acc_rd_0_data_bits_0_28; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_29 = io_acc_rd_0_data_bits_0_29; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_30 = io_acc_rd_0_data_bits_0_30; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_acc_i_data_bits_0_31 = io_acc_rd_0_data_bits_0_31; // @[TensorGemm.scala 709:68]
  assign mvc_0_io_bypass_cond = wrpipe_0_io_deq_bits == wrpipe2_io_deq_bits & wrpipe_0_io_deq_valid &
    wrpipe2_io_deq_valid; // @[TensorGemm.scala 695:85]
  assign wrpipe2_clock = clock;
  assign wrpipe2_reset = reset;
  assign wrpipe2_io_enq_valid = wrpipe_0_io_deq_valid; // @[TensorGemm.scala 692:20]
  assign wrpipe2_io_enq_bits = wrpipe_0_io_deq_bits; // @[TensorGemm.scala 692:20]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      delayed_valid <= 1'h0; // @[Reg.scala 28:20]
    end else begin
      delayed_valid <= _GEN_0;
    end
    delayed_acc_i <= m_io_acc_i; // @[Reg.scala 16:16 17:{18,22}]
    delayed_inp_i <= m_io_inp_i; // @[Reg.scala 16:16 17:{18,22}]
    delayed_wgt_i <= m_io_wgt_i; // @[Reg.scala 16:16 17:{18,22}]
    if (reset) begin // @[TensorGemm.scala 566:22]
      state <= 2'h0; // @[TensorGemm.scala 566:22]
    end else if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      state <= 2'h1; // @[TensorGemm.scala 573:11]
    end else if (state == 2'h1 & m_io_last) begin // @[TensorGemm.scala 577:43]
      state <= 2'h2; // @[TensorGemm.scala 578:11]
    end else if (state == 2'h2 & inflight == 4'h0) begin // @[TensorGemm.scala 579:51]
      state <= 2'h0; // @[TensorGemm.scala 580:11]
    end
    if (reset) begin // @[TensorGemm.scala 567:25]
      inflight <= 4'h0; // @[TensorGemm.scala 567:25]
    end else if (_T) begin // @[TensorGemm.scala 662:25]
      inflight <= 4'h0; // @[TensorGemm.scala 664:14]
    end else if (!(m_io_valid & wrpipeNs_io_deq_valid)) begin // @[TensorGemm.scala 654:45]
      if (m_io_valid) begin // @[TensorGemm.scala 655:26]
        inflight <= _inflight_T_1; // @[TensorGemm.scala 657:14]
      end else begin
        inflight <= _GEN_27;
      end
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_wgt_1 <= io_dec_wgt_1; // @[TensorGemm.scala 574:17]
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_wgt_0 <= io_dec_wgt_0; // @[TensorGemm.scala 574:17]
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_inp_1 <= io_dec_inp_1; // @[TensorGemm.scala 574:17]
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_inp_0 <= io_dec_inp_0; // @[TensorGemm.scala 574:17]
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_acc_1 <= io_dec_acc_1; // @[TensorGemm.scala 574:17]
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_acc_0 <= io_dec_acc_0; // @[TensorGemm.scala 574:17]
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_empty_0 <= io_dec_empty_0; // @[TensorGemm.scala 574:17]
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_lp_1 <= io_dec_lp_1; // @[TensorGemm.scala 574:17]
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_lp_0 <= io_dec_lp_0; // @[TensorGemm.scala 574:17]
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_uop_end <= io_dec_uop_end; // @[TensorGemm.scala 574:17]
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_uop_begin <= io_dec_uop_begin; // @[TensorGemm.scala 574:17]
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_reset <= io_dec_reset; // @[TensorGemm.scala 574:17]
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_push_next <= io_dec_push_next; // @[TensorGemm.scala 574:17]
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_push_prev <= io_dec_push_prev; // @[TensorGemm.scala 574:17]
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_pop_next <= io_dec_pop_next; // @[TensorGemm.scala 574:17]
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_pop_prev <= io_dec_pop_prev; // @[TensorGemm.scala 574:17]
    end
    if (state == 2'h0 & io_start) begin // @[TensorGemm.scala 572:37]
      capture_dec_op <= io_dec_op; // @[TensorGemm.scala 574:17]
    end
    if (reset) begin // @[TensorGemm.scala 618:34]
      delayed_uop_valid <= 1'h0; // @[TensorGemm.scala 618:34]
    end else begin
      delayed_uop_valid <= delayed_valid; // @[TensorGemm.scala 618:34]
    end
    if (reset) begin // @[TensorGemm.scala 623:40]
      io_acc_rd_0_idx_valid_REG <= 1'h0; // @[TensorGemm.scala 623:40]
    end else begin
      io_acc_rd_0_idx_valid_REG <= acc_idx_pipe_io_deq_valid; // @[TensorGemm.scala 623:40]
    end
    io_acc_rd_0_idx_bits_REG <= acc_idx_pipe_io_deq_bits; // @[TensorGemm.scala 624:39]
    if (reset) begin // @[TensorGemm.scala 698:40]
      mvc_0_io_valid_reset_REG <= 1'h0; // @[TensorGemm.scala 698:40]
    end else begin
      mvc_0_io_valid_reset_REG <= reset_pipe_io_deq_bits & reset_pipe_io_deq_valid; // @[TensorGemm.scala 698:40]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(state != 2'h1 | _T_8 == _T_9)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorGemm.scala:585 assert(state =/= sRun  || capture_dec.asUInt === io.dec.asUInt)\n"
            ); // @[TensorGemm.scala 585:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & ~(state != 2'h2 | _T_10)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorGemm.scala:586 assert(state =/= sWait || capture_dec.asUInt === io.dec.asUInt)\n"
            ); // @[TensorGemm.scala 586:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & ~(io_uop_data_valid == delayed_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorGemm.scala:596 assert(delayedUopData.valid === delayed_valid)\n"); // @[TensorGemm.scala 596:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & ~(io_inp_rd_0_data_valid == delayed_uop_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorGemm.scala:621 assert(io.inp.rd(0).data.valid === delayed_uop_valid)\n"); // @[TensorGemm.scala 621:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & ~(io_wgt_rd_0_data_valid == delayed_uop_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorGemm.scala:630 assert(io.wgt.rd(idx).data.valid === ShiftRegister(delayed_uop_valid, scratchpadReadLatency))\n"
            ); // @[TensorGemm.scala 630:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & ~(io_acc_rd_0_data_valid == wrpipe_0_io_deq_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorGemm.scala:651 assert(io.acc.rd(idx).data.valid === wrpipe(idx).io.deq.valid)\n"
            ); // @[TensorGemm.scala 651:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_39 & m_io_valid & _T_13 & ~(inflight != 4'hf)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorGemm.scala:656 assert(inflight =/= ((1<<inflightBits)-1).U)\n"); // @[TensorGemm.scala 656:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_34 & ~m_io_valid & wrpipeNs_io_deq_valid & _T_13 & ~(inflight != 4'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TensorGemm.scala:659 assert(inflight =/= 0.U)\n"); // @[TensorGemm.scala 659:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & _T_13 & ~_T_5) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TensorGemm.scala:663 assert(inflight === 0.U)\n"); // @[TensorGemm.scala 663:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13 & ~(mvc_0_io_acc_o_data_valid == (wrpipe_0_io_deq_valid | mvc_0_io_valid_reset))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorGemm.scala:704 assert(mvc(idx1).io.acc_o.data.valid === (wrpipe(idx1).io.deq.valid | mvc(idx1).io.valid_reset))\n"
            ); // @[TensorGemm.scala 704:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  delayed_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  delayed_acc_i = _RAND_1[6:0];
  _RAND_2 = {1{`RANDOM}};
  delayed_inp_i = _RAND_2[6:0];
  _RAND_3 = {1{`RANDOM}};
  delayed_wgt_i = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  inflight = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  capture_dec_wgt_1 = _RAND_6[9:0];
  _RAND_7 = {1{`RANDOM}};
  capture_dec_wgt_0 = _RAND_7[9:0];
  _RAND_8 = {1{`RANDOM}};
  capture_dec_inp_1 = _RAND_8[10:0];
  _RAND_9 = {1{`RANDOM}};
  capture_dec_inp_0 = _RAND_9[10:0];
  _RAND_10 = {1{`RANDOM}};
  capture_dec_acc_1 = _RAND_10[10:0];
  _RAND_11 = {1{`RANDOM}};
  capture_dec_acc_0 = _RAND_11[10:0];
  _RAND_12 = {1{`RANDOM}};
  capture_dec_empty_0 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  capture_dec_lp_1 = _RAND_13[13:0];
  _RAND_14 = {1{`RANDOM}};
  capture_dec_lp_0 = _RAND_14[13:0];
  _RAND_15 = {1{`RANDOM}};
  capture_dec_uop_end = _RAND_15[13:0];
  _RAND_16 = {1{`RANDOM}};
  capture_dec_uop_begin = _RAND_16[12:0];
  _RAND_17 = {1{`RANDOM}};
  capture_dec_reset = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  capture_dec_push_next = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  capture_dec_push_prev = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  capture_dec_pop_next = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  capture_dec_pop_prev = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  capture_dec_op = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  delayed_uop_valid = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  io_acc_rd_0_idx_valid_REG = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  io_acc_rd_0_idx_bits_REG = _RAND_25[6:0];
  _RAND_26 = {1{`RANDOM}};
  mvc_0_io_valid_reset_REG = _RAND_26[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(state != 2'h1 | _T_8 == _T_9); // @[TensorGemm.scala 585:9]
    end
    //
    if (_T_13) begin
      assert(state != 2'h2 | _T_10); // @[TensorGemm.scala 586:9]
    end
    //
    if (_T_13) begin
      assert(io_uop_data_valid == delayed_valid); // @[TensorGemm.scala 596:9]
    end
    //
    if (_T_13) begin
      assert(io_inp_rd_0_data_valid == delayed_uop_valid); // @[TensorGemm.scala 621:9]
    end
    //
    if (_T_13) begin
      assert(io_wgt_rd_0_data_valid == delayed_uop_valid); // @[TensorGemm.scala 630:11]
    end
    //
    if (_T_13) begin
      assert(io_acc_rd_0_data_valid == wrpipe_0_io_deq_valid); // @[TensorGemm.scala 651:11]
    end
    //
    if (~_T_39 & m_io_valid & _T_13) begin
      assert(inflight != 4'hf); // @[TensorGemm.scala 656:11]
    end
    //
    if (_GEN_34 & ~m_io_valid & wrpipeNs_io_deq_valid & _T_13) begin
      assert(inflight != 4'h0); // @[TensorGemm.scala 659:11]
    end
    //
    if (_T & _T_13) begin
      assert(_T_5); // @[TensorGemm.scala 663:11]
    end
    //
    if (_T_13) begin
      assert(mvc_0_io_acc_o_data_valid == (wrpipe_0_io_deq_valid | mvc_0_io_valid_reset)); // @[TensorGemm.scala 704:11]
    end
  end
endmodule
module TensorAluIndexGenerator(
  input         clock,
  input         reset,
  input         io_start,
  output        io_last,
  input         io_dec_alu_use_imm,
  input  [10:0] io_dec_src_1,
  input  [10:0] io_dec_src_0,
  input  [10:0] io_dec_dst_1,
  input  [10:0] io_dec_dst_0,
  input  [13:0] io_dec_lp_1,
  input  [13:0] io_dec_lp_0,
  input  [13:0] io_dec_uop_end,
  input  [12:0] io_dec_uop_begin,
  output        io_valid,
  output        io_src_valid,
  output [6:0]  io_dst_idx,
  output [6:0]  io_src_idx,
  output [6:0]  io_uop_idx
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
`endif // RANDOMIZE_REG_INIT
  reg  running; // @[TensorAlu.scala 119:24]
  reg  stutter; // @[TensorAlu.scala 120:24]
  wire  advance = io_dec_alu_use_imm | stutter; // @[TensorAlu.scala 122:36]
  wire  _T = ~running; // @[TensorAlu.scala 124:8]
  wire  _T_2 = ~advance; // @[TensorAlu.scala 126:26]
  wire  _GEN_0 = io_last ? 1'h0 : running; // @[TensorAlu.scala 129:20 130:15 119:24]
  wire  _GEN_1 = running & advance ? _GEN_0 : running; // @[TensorAlu.scala 119:24 128:35]
  wire  _GEN_2 = running & advance ? 1'h0 : stutter; // @[TensorAlu.scala 128:35 132:13 120:24]
  wire  _GEN_3 = running & ~advance | _GEN_2; // @[TensorAlu.scala 126:36 127:13]
  wire  _GEN_4 = running & ~advance ? running : _GEN_1; // @[TensorAlu.scala 119:24 126:36]
  wire  _GEN_5 = ~running & io_start | _GEN_4; // @[TensorAlu.scala 124:30 125:13]
  reg [13:0] cnt_i; // @[TensorAlu.scala 135:18]
  reg [6:0] dst_i; // @[TensorAlu.scala 136:18]
  reg [6:0] src_i; // @[TensorAlu.scala 137:18]
  reg [13:0] cnt_o; // @[TensorAlu.scala 139:18]
  reg [6:0] dst_o; // @[TensorAlu.scala 140:18]
  reg [6:0] src_o; // @[TensorAlu.scala 141:18]
  reg [13:0] uop_idx; // @[TensorAlu.scala 143:20]
  wire [13:0] _T_7 = io_dec_uop_end - 14'h1; // @[TensorAlu.scala 158:38]
  wire [13:0] _uop_idx_T_1 = uop_idx + 14'h1; // @[TensorAlu.scala 159:26]
  wire [13:0] _T_10 = io_dec_lp_1 - 14'h1; // @[TensorAlu.scala 162:35]
  wire [13:0] _cnt_i_T_1 = cnt_i + 14'h1; // @[TensorAlu.scala 163:24]
  wire [10:0] _GEN_45 = {{4'd0}, dst_i}; // @[TensorAlu.scala 164:24]
  wire [10:0] _dst_i_T_1 = _GEN_45 + io_dec_dst_1; // @[TensorAlu.scala 164:24]
  wire [10:0] _GEN_46 = {{4'd0}, src_i}; // @[TensorAlu.scala 165:24]
  wire [10:0] _src_i_T_1 = _GEN_46 + io_dec_src_1; // @[TensorAlu.scala 165:24]
  wire [13:0] _T_13 = io_dec_lp_0 - 14'h1; // @[TensorAlu.scala 167:37]
  wire [10:0] _GEN_47 = {{4'd0}, dst_o}; // @[TensorAlu.scala 168:31]
  wire [10:0] dst_tmp = _GEN_47 + io_dec_dst_0; // @[TensorAlu.scala 168:31]
  wire [10:0] _GEN_48 = {{4'd0}, src_o}; // @[TensorAlu.scala 169:31]
  wire [10:0] src_tmp = _GEN_48 + io_dec_src_0; // @[TensorAlu.scala 169:31]
  wire [13:0] _cnt_o_T_1 = cnt_o + 14'h1; // @[TensorAlu.scala 170:26]
  wire [13:0] _GEN_7 = cnt_o != _T_13 ? _cnt_o_T_1 : cnt_o; // @[TensorAlu.scala 167:44 170:17 139:18]
  wire [10:0] _GEN_8 = cnt_o != _T_13 ? dst_tmp : {{4'd0}, dst_o}; // @[TensorAlu.scala 167:44 171:17 140:18]
  wire [10:0] _GEN_9 = cnt_o != _T_13 ? src_tmp : {{4'd0}, src_o}; // @[TensorAlu.scala 167:44 172:17 141:18]
  wire [13:0] _GEN_10 = cnt_o != _T_13 ? 14'h0 : cnt_i; // @[TensorAlu.scala 167:44 173:17 135:18]
  wire [10:0] _GEN_11 = cnt_o != _T_13 ? dst_tmp : {{4'd0}, dst_i}; // @[TensorAlu.scala 167:44 174:17 136:18]
  wire [10:0] _GEN_12 = cnt_o != _T_13 ? src_tmp : {{4'd0}, src_i}; // @[TensorAlu.scala 167:44 175:17 137:18]
  wire  _GEN_13 = cnt_o != _T_13 ? 1'h0 : 1'h1; // @[TensorAlu.scala 117:11 167:44 177:19]
  wire [10:0] _GEN_15 = cnt_i != _T_10 ? _dst_i_T_1 : _GEN_11; // @[TensorAlu.scala 162:42 164:15]
  wire [10:0] _GEN_16 = cnt_i != _T_10 ? _src_i_T_1 : _GEN_12; // @[TensorAlu.scala 162:42 165:15]
  wire [10:0] _GEN_18 = cnt_i != _T_10 ? {{4'd0}, dst_o} : _GEN_8; // @[TensorAlu.scala 140:18 162:42]
  wire [10:0] _GEN_19 = cnt_i != _T_10 ? {{4'd0}, src_o} : _GEN_9; // @[TensorAlu.scala 141:18 162:42]
  wire  _GEN_20 = cnt_i != _T_10 ? 1'h0 : _GEN_13; // @[TensorAlu.scala 117:11 162:42]
  wire [10:0] _GEN_23 = uop_idx != _T_7 ? {{4'd0}, dst_i} : _GEN_15; // @[TensorAlu.scala 136:18 158:45]
  wire [10:0] _GEN_24 = uop_idx != _T_7 ? {{4'd0}, src_i} : _GEN_16; // @[TensorAlu.scala 137:18 158:45]
  wire [10:0] _GEN_26 = uop_idx != _T_7 ? {{4'd0}, dst_o} : _GEN_18; // @[TensorAlu.scala 140:18 158:45]
  wire [10:0] _GEN_27 = uop_idx != _T_7 ? {{4'd0}, src_o} : _GEN_19; // @[TensorAlu.scala 141:18 158:45]
  wire  _GEN_28 = uop_idx != _T_7 ? 1'h0 : _GEN_20; // @[TensorAlu.scala 117:11 158:45]
  wire [10:0] _GEN_31 = advance ? _GEN_23 : {{4'd0}, dst_i}; // @[TensorAlu.scala 136:18 157:25]
  wire [10:0] _GEN_32 = advance ? _GEN_24 : {{4'd0}, src_i}; // @[TensorAlu.scala 137:18 157:25]
  wire [10:0] _GEN_34 = advance ? _GEN_26 : {{4'd0}, dst_o}; // @[TensorAlu.scala 140:18 157:25]
  wire [10:0] _GEN_35 = advance ? _GEN_27 : {{4'd0}, src_o}; // @[TensorAlu.scala 141:18 157:25]
  wire  _GEN_36 = advance & _GEN_28; // @[TensorAlu.scala 117:11 157:25]
  wire [10:0] _GEN_38 = _T ? 11'h0 : _GEN_31; // @[TensorAlu.scala 153:18 154:25]
  wire [10:0] _GEN_39 = _T ? 11'h0 : _GEN_32; // @[TensorAlu.scala 153:18 154:39]
  wire [10:0] _GEN_41 = _T ? 11'h0 : _GEN_34; // @[TensorAlu.scala 153:18 155:25]
  wire [10:0] _GEN_42 = _T ? 11'h0 : _GEN_35; // @[TensorAlu.scala 153:18 155:39]
  assign io_last = _T ? 1'h0 : _GEN_36; // @[TensorAlu.scala 117:11 153:18]
  assign io_valid = running & advance; // @[TensorAlu.scala 145:23]
  assign io_src_valid = running & _T_2; // @[TensorAlu.scala 146:27]
  assign io_dst_idx = dst_i; // @[TensorAlu.scala 147:14]
  assign io_src_idx = src_i; // @[TensorAlu.scala 148:14]
  assign io_uop_idx = uop_idx[6:0]; // @[TensorAlu.scala 149:14]
  always @(posedge clock) begin
    if (reset) begin // @[TensorAlu.scala 119:24]
      running <= 1'h0; // @[TensorAlu.scala 119:24]
    end else begin
      running <= _GEN_5;
    end
    if (reset) begin // @[TensorAlu.scala 120:24]
      stutter <= 1'h0; // @[TensorAlu.scala 120:24]
    end else if (!(~running & io_start)) begin // @[TensorAlu.scala 124:30]
      stutter <= _GEN_3;
    end
    if (_T) begin // @[TensorAlu.scala 153:18]
      cnt_i <= 14'h0; // @[TensorAlu.scala 154:11]
    end else if (advance) begin // @[TensorAlu.scala 157:25]
      if (!(uop_idx != _T_7)) begin // @[TensorAlu.scala 158:45]
        if (cnt_i != _T_10) begin // @[TensorAlu.scala 162:42]
          cnt_i <= _cnt_i_T_1; // @[TensorAlu.scala 163:15]
        end else begin
          cnt_i <= _GEN_10;
        end
      end
    end
    dst_i <= _GEN_38[6:0];
    src_i <= _GEN_39[6:0];
    if (_T) begin // @[TensorAlu.scala 153:18]
      cnt_o <= 14'h0; // @[TensorAlu.scala 155:11]
    end else if (advance) begin // @[TensorAlu.scala 157:25]
      if (!(uop_idx != _T_7)) begin // @[TensorAlu.scala 158:45]
        if (!(cnt_i != _T_10)) begin // @[TensorAlu.scala 162:42]
          cnt_o <= _GEN_7;
        end
      end
    end
    dst_o <= _GEN_41[6:0];
    src_o <= _GEN_42[6:0];
    if (_T) begin // @[TensorAlu.scala 153:18]
      uop_idx <= {{1'd0}, io_dec_uop_begin}; // @[TensorAlu.scala 156:13]
    end else if (advance) begin // @[TensorAlu.scala 157:25]
      if (uop_idx != _T_7) begin // @[TensorAlu.scala 158:45]
        uop_idx <= _uop_idx_T_1; // @[TensorAlu.scala 159:15]
      end else begin
        uop_idx <= {{1'd0}, io_dec_uop_begin}; // @[TensorAlu.scala 161:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  running = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  stutter = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  cnt_i = _RAND_2[13:0];
  _RAND_3 = {1{`RANDOM}};
  dst_i = _RAND_3[6:0];
  _RAND_4 = {1{`RANDOM}};
  src_i = _RAND_4[6:0];
  _RAND_5 = {1{`RANDOM}};
  cnt_o = _RAND_5[13:0];
  _RAND_6 = {1{`RANDOM}};
  dst_o = _RAND_6[6:0];
  _RAND_7 = {1{`RANDOM}};
  src_o = _RAND_7[6:0];
  _RAND_8 = {1{`RANDOM}};
  uop_idx = _RAND_8[13:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Alu(
  input  [2:0]  io_opcode,
  input  [31:0] io_a,
  input  [31:0] io_b,
  output [31:0] io_y
);
  wire [31:0] ub = io_b; // @[TensorAlu.scala 37:17]
  wire [4:0] _m_T_1 = ~ub[4:0]; // @[TensorAlu.scala 39:11]
  wire [4:0] m = _m_T_1 + 5'h1; // @[TensorAlu.scala 39:29]
  wire [31:0] fop_0 = $signed(io_a) < $signed(io_b) ? $signed(io_a) : $signed(io_b); // @[TensorAlu.scala 43:20]
  wire [31:0] fop_1 = $signed(io_a) < $signed(io_b) ? $signed(io_b) : $signed(io_a); // @[TensorAlu.scala 43:50]
  wire [31:0] fop_2 = $signed(io_a) + $signed(io_b); // @[TensorAlu.scala 44:10]
  wire [31:0] fop_3 = $signed(io_a) >>> ub[4:0]; // @[TensorAlu.scala 44:23]
  wire [62:0] _GEN_1 = {{31{io_a[31]}},io_a}; // @[TensorAlu.scala 44:34]
  wire [62:0] fop_4 = $signed(_GEN_1) << m; // @[TensorAlu.scala 44:34]
  wire [31:0] _io_y_T_1 = 3'h0 == io_opcode ? $signed(fop_0) : $signed(io_a); // @[Mux.scala 81:58]
  wire [31:0] _io_y_T_3 = 3'h1 == io_opcode ? $signed(fop_1) : $signed(_io_y_T_1); // @[Mux.scala 81:58]
  wire [31:0] _io_y_T_5 = 3'h2 == io_opcode ? $signed(fop_2) : $signed(_io_y_T_3); // @[Mux.scala 81:58]
  wire [31:0] _io_y_T_7 = 3'h3 == io_opcode ? $signed(fop_3) : $signed(_io_y_T_5); // @[Mux.scala 81:58]
  wire [62:0] _io_y_T_9 = 3'h4 == io_opcode ? $signed(fop_4) : $signed({{31{_io_y_T_7[31]}},_io_y_T_7}); // @[Mux.scala 81:58]
  assign io_y = _io_y_T_9[31:0]; // @[TensorAlu.scala 47:8]
endmodule
module AluReg(
  input         clock,
  input  [2:0]  io_opcode,
  input         io_a_valid,
  input  [31:0] io_a_bits,
  input         io_b_valid,
  input  [31:0] io_b_bits,
  output        io_y_valid,
  output [31:0] io_y_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] alu_io_opcode; // @[TensorAlu.scala 58:19]
  wire [31:0] alu_io_a; // @[TensorAlu.scala 58:19]
  wire [31:0] alu_io_b; // @[TensorAlu.scala 58:19]
  wire [31:0] alu_io_y; // @[TensorAlu.scala 58:19]
  reg [31:0] rA; // @[Reg.scala 16:16]
  reg [31:0] rB; // @[Reg.scala 16:16]
  reg  valid; // @[TensorAlu.scala 61:22]
  Alu alu ( // @[TensorAlu.scala 58:19]
    .io_opcode(alu_io_opcode),
    .io_a(alu_io_a),
    .io_b(alu_io_b),
    .io_y(alu_io_y)
  );
  assign io_y_valid = valid; // @[TensorAlu.scala 70:14]
  assign io_y_bits = alu_io_y; // @[TensorAlu.scala 71:25]
  assign alu_io_opcode = io_opcode; // @[TensorAlu.scala 63:17]
  assign alu_io_a = rA; // @[TensorAlu.scala 66:18]
  assign alu_io_b = rB; // @[TensorAlu.scala 67:18]
  always @(posedge clock) begin
    if (io_a_valid) begin // @[Reg.scala 17:18]
      rA <= io_a_bits; // @[Reg.scala 17:22]
    end
    if (io_b_valid) begin // @[Reg.scala 17:18]
      rB <= io_b_bits; // @[Reg.scala 17:22]
    end
    valid <= io_b_valid; // @[TensorAlu.scala 61:22]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rA = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  rB = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  valid = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module AluVector(
  input         clock,
  input  [2:0]  io_opcode,
  input         io_acc_a_data_valid,
  input  [31:0] io_acc_a_data_bits_0_0,
  input  [31:0] io_acc_a_data_bits_0_1,
  input  [31:0] io_acc_a_data_bits_0_2,
  input  [31:0] io_acc_a_data_bits_0_3,
  input  [31:0] io_acc_a_data_bits_0_4,
  input  [31:0] io_acc_a_data_bits_0_5,
  input  [31:0] io_acc_a_data_bits_0_6,
  input  [31:0] io_acc_a_data_bits_0_7,
  input  [31:0] io_acc_a_data_bits_0_8,
  input  [31:0] io_acc_a_data_bits_0_9,
  input  [31:0] io_acc_a_data_bits_0_10,
  input  [31:0] io_acc_a_data_bits_0_11,
  input  [31:0] io_acc_a_data_bits_0_12,
  input  [31:0] io_acc_a_data_bits_0_13,
  input  [31:0] io_acc_a_data_bits_0_14,
  input  [31:0] io_acc_a_data_bits_0_15,
  input  [31:0] io_acc_a_data_bits_0_16,
  input  [31:0] io_acc_a_data_bits_0_17,
  input  [31:0] io_acc_a_data_bits_0_18,
  input  [31:0] io_acc_a_data_bits_0_19,
  input  [31:0] io_acc_a_data_bits_0_20,
  input  [31:0] io_acc_a_data_bits_0_21,
  input  [31:0] io_acc_a_data_bits_0_22,
  input  [31:0] io_acc_a_data_bits_0_23,
  input  [31:0] io_acc_a_data_bits_0_24,
  input  [31:0] io_acc_a_data_bits_0_25,
  input  [31:0] io_acc_a_data_bits_0_26,
  input  [31:0] io_acc_a_data_bits_0_27,
  input  [31:0] io_acc_a_data_bits_0_28,
  input  [31:0] io_acc_a_data_bits_0_29,
  input  [31:0] io_acc_a_data_bits_0_30,
  input  [31:0] io_acc_a_data_bits_0_31,
  input         io_acc_b_data_valid,
  input  [31:0] io_acc_b_data_bits_0_0,
  input  [31:0] io_acc_b_data_bits_0_1,
  input  [31:0] io_acc_b_data_bits_0_2,
  input  [31:0] io_acc_b_data_bits_0_3,
  input  [31:0] io_acc_b_data_bits_0_4,
  input  [31:0] io_acc_b_data_bits_0_5,
  input  [31:0] io_acc_b_data_bits_0_6,
  input  [31:0] io_acc_b_data_bits_0_7,
  input  [31:0] io_acc_b_data_bits_0_8,
  input  [31:0] io_acc_b_data_bits_0_9,
  input  [31:0] io_acc_b_data_bits_0_10,
  input  [31:0] io_acc_b_data_bits_0_11,
  input  [31:0] io_acc_b_data_bits_0_12,
  input  [31:0] io_acc_b_data_bits_0_13,
  input  [31:0] io_acc_b_data_bits_0_14,
  input  [31:0] io_acc_b_data_bits_0_15,
  input  [31:0] io_acc_b_data_bits_0_16,
  input  [31:0] io_acc_b_data_bits_0_17,
  input  [31:0] io_acc_b_data_bits_0_18,
  input  [31:0] io_acc_b_data_bits_0_19,
  input  [31:0] io_acc_b_data_bits_0_20,
  input  [31:0] io_acc_b_data_bits_0_21,
  input  [31:0] io_acc_b_data_bits_0_22,
  input  [31:0] io_acc_b_data_bits_0_23,
  input  [31:0] io_acc_b_data_bits_0_24,
  input  [31:0] io_acc_b_data_bits_0_25,
  input  [31:0] io_acc_b_data_bits_0_26,
  input  [31:0] io_acc_b_data_bits_0_27,
  input  [31:0] io_acc_b_data_bits_0_28,
  input  [31:0] io_acc_b_data_bits_0_29,
  input  [31:0] io_acc_b_data_bits_0_30,
  input  [31:0] io_acc_b_data_bits_0_31,
  output        io_acc_y_data_valid,
  output [31:0] io_acc_y_data_bits_0_0,
  output [31:0] io_acc_y_data_bits_0_1,
  output [31:0] io_acc_y_data_bits_0_2,
  output [31:0] io_acc_y_data_bits_0_3,
  output [31:0] io_acc_y_data_bits_0_4,
  output [31:0] io_acc_y_data_bits_0_5,
  output [31:0] io_acc_y_data_bits_0_6,
  output [31:0] io_acc_y_data_bits_0_7,
  output [31:0] io_acc_y_data_bits_0_8,
  output [31:0] io_acc_y_data_bits_0_9,
  output [31:0] io_acc_y_data_bits_0_10,
  output [31:0] io_acc_y_data_bits_0_11,
  output [31:0] io_acc_y_data_bits_0_12,
  output [31:0] io_acc_y_data_bits_0_13,
  output [31:0] io_acc_y_data_bits_0_14,
  output [31:0] io_acc_y_data_bits_0_15,
  output [31:0] io_acc_y_data_bits_0_16,
  output [31:0] io_acc_y_data_bits_0_17,
  output [31:0] io_acc_y_data_bits_0_18,
  output [31:0] io_acc_y_data_bits_0_19,
  output [31:0] io_acc_y_data_bits_0_20,
  output [31:0] io_acc_y_data_bits_0_21,
  output [31:0] io_acc_y_data_bits_0_22,
  output [31:0] io_acc_y_data_bits_0_23,
  output [31:0] io_acc_y_data_bits_0_24,
  output [31:0] io_acc_y_data_bits_0_25,
  output [31:0] io_acc_y_data_bits_0_26,
  output [31:0] io_acc_y_data_bits_0_27,
  output [31:0] io_acc_y_data_bits_0_28,
  output [31:0] io_acc_y_data_bits_0_29,
  output [31:0] io_acc_y_data_bits_0_30,
  output [31:0] io_acc_y_data_bits_0_31,
  output        io_out_data_valid,
  output [7:0]  io_out_data_bits_0_0,
  output [7:0]  io_out_data_bits_0_1,
  output [7:0]  io_out_data_bits_0_2,
  output [7:0]  io_out_data_bits_0_3,
  output [7:0]  io_out_data_bits_0_4,
  output [7:0]  io_out_data_bits_0_5,
  output [7:0]  io_out_data_bits_0_6,
  output [7:0]  io_out_data_bits_0_7,
  output [7:0]  io_out_data_bits_0_8,
  output [7:0]  io_out_data_bits_0_9,
  output [7:0]  io_out_data_bits_0_10,
  output [7:0]  io_out_data_bits_0_11,
  output [7:0]  io_out_data_bits_0_12,
  output [7:0]  io_out_data_bits_0_13,
  output [7:0]  io_out_data_bits_0_14,
  output [7:0]  io_out_data_bits_0_15,
  output [7:0]  io_out_data_bits_0_16,
  output [7:0]  io_out_data_bits_0_17,
  output [7:0]  io_out_data_bits_0_18,
  output [7:0]  io_out_data_bits_0_19,
  output [7:0]  io_out_data_bits_0_20,
  output [7:0]  io_out_data_bits_0_21,
  output [7:0]  io_out_data_bits_0_22,
  output [7:0]  io_out_data_bits_0_23,
  output [7:0]  io_out_data_bits_0_24,
  output [7:0]  io_out_data_bits_0_25,
  output [7:0]  io_out_data_bits_0_26,
  output [7:0]  io_out_data_bits_0_27,
  output [7:0]  io_out_data_bits_0_28,
  output [7:0]  io_out_data_bits_0_29,
  output [7:0]  io_out_data_bits_0_30,
  output [7:0]  io_out_data_bits_0_31
);
  wire  f_0_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_0_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_0_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_0_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_0_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_0_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_0_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_0_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_1_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_1_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_1_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_1_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_1_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_1_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_1_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_1_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_2_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_2_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_2_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_2_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_2_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_2_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_2_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_2_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_3_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_3_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_3_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_3_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_3_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_3_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_3_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_3_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_4_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_4_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_4_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_4_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_4_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_4_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_4_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_4_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_5_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_5_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_5_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_5_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_5_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_5_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_5_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_5_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_6_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_6_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_6_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_6_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_6_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_6_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_6_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_6_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_7_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_7_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_7_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_7_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_7_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_7_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_7_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_7_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_8_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_8_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_8_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_8_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_8_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_8_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_8_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_8_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_9_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_9_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_9_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_9_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_9_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_9_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_9_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_9_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_10_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_10_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_10_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_10_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_10_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_10_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_10_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_10_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_11_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_11_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_11_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_11_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_11_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_11_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_11_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_11_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_12_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_12_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_12_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_12_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_12_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_12_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_12_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_12_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_13_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_13_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_13_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_13_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_13_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_13_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_13_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_13_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_14_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_14_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_14_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_14_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_14_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_14_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_14_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_14_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_15_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_15_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_15_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_15_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_15_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_15_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_15_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_15_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_16_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_16_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_16_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_16_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_16_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_16_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_16_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_16_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_17_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_17_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_17_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_17_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_17_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_17_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_17_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_17_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_18_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_18_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_18_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_18_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_18_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_18_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_18_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_18_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_19_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_19_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_19_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_19_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_19_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_19_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_19_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_19_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_20_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_20_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_20_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_20_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_20_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_20_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_20_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_20_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_21_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_21_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_21_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_21_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_21_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_21_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_21_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_21_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_22_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_22_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_22_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_22_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_22_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_22_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_22_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_22_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_23_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_23_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_23_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_23_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_23_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_23_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_23_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_23_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_24_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_24_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_24_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_24_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_24_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_24_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_24_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_24_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_25_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_25_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_25_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_25_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_25_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_25_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_25_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_25_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_26_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_26_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_26_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_26_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_26_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_26_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_26_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_26_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_27_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_27_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_27_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_27_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_27_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_27_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_27_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_27_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_28_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_28_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_28_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_28_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_28_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_28_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_28_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_28_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_29_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_29_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_29_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_29_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_29_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_29_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_29_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_29_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_30_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_30_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_30_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_30_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_30_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_30_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_30_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_30_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  f_31_clock; // @[TensorAlu.scala 84:36]
  wire [2:0] f_31_io_opcode; // @[TensorAlu.scala 84:36]
  wire  f_31_io_a_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_31_io_a_bits; // @[TensorAlu.scala 84:36]
  wire  f_31_io_b_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_31_io_b_bits; // @[TensorAlu.scala 84:36]
  wire  f_31_io_y_valid; // @[TensorAlu.scala 84:36]
  wire [31:0] f_31_io_y_bits; // @[TensorAlu.scala 84:36]
  wire  valid_1 = f_1_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_0 = f_0_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_3 = f_3_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_2 = f_2_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_5 = f_5_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_4 = f_4_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_7 = f_7_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_6 = f_6_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire [7:0] io_acc_y_data_valid_lo_lo = {valid_7,valid_6,valid_5,valid_4,valid_3,valid_2,valid_1,valid_0}; // @[TensorAlu.scala 96:32]
  wire  valid_9 = f_9_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_8 = f_8_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_11 = f_11_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_10 = f_10_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_13 = f_13_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_12 = f_12_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_15 = f_15_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_14 = f_14_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire [15:0] io_acc_y_data_valid_lo = {valid_15,valid_14,valid_13,valid_12,valid_11,valid_10,valid_9,valid_8,
    io_acc_y_data_valid_lo_lo}; // @[TensorAlu.scala 96:32]
  wire  valid_17 = f_17_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_16 = f_16_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_19 = f_19_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_18 = f_18_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_21 = f_21_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_20 = f_20_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_23 = f_23_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_22 = f_22_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire [7:0] io_acc_y_data_valid_hi_lo = {valid_23,valid_22,valid_21,valid_20,valid_19,valid_18,valid_17,valid_16}; // @[TensorAlu.scala 96:32]
  wire  valid_25 = f_25_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_24 = f_24_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_27 = f_27_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_26 = f_26_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_29 = f_29_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_28 = f_28_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_31 = f_31_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire  valid_30 = f_30_io_y_valid; // @[TensorAlu.scala 85:19 92:14]
  wire [31:0] _io_acc_y_data_valid_T = {valid_31,valid_30,valid_29,valid_28,valid_27,valid_26,valid_25,valid_24,
    io_acc_y_data_valid_hi_lo,io_acc_y_data_valid_lo}; // @[TensorAlu.scala 96:32]
  AluReg f_0 ( // @[TensorAlu.scala 84:36]
    .clock(f_0_clock),
    .io_opcode(f_0_io_opcode),
    .io_a_valid(f_0_io_a_valid),
    .io_a_bits(f_0_io_a_bits),
    .io_b_valid(f_0_io_b_valid),
    .io_b_bits(f_0_io_b_bits),
    .io_y_valid(f_0_io_y_valid),
    .io_y_bits(f_0_io_y_bits)
  );
  AluReg f_1 ( // @[TensorAlu.scala 84:36]
    .clock(f_1_clock),
    .io_opcode(f_1_io_opcode),
    .io_a_valid(f_1_io_a_valid),
    .io_a_bits(f_1_io_a_bits),
    .io_b_valid(f_1_io_b_valid),
    .io_b_bits(f_1_io_b_bits),
    .io_y_valid(f_1_io_y_valid),
    .io_y_bits(f_1_io_y_bits)
  );
  AluReg f_2 ( // @[TensorAlu.scala 84:36]
    .clock(f_2_clock),
    .io_opcode(f_2_io_opcode),
    .io_a_valid(f_2_io_a_valid),
    .io_a_bits(f_2_io_a_bits),
    .io_b_valid(f_2_io_b_valid),
    .io_b_bits(f_2_io_b_bits),
    .io_y_valid(f_2_io_y_valid),
    .io_y_bits(f_2_io_y_bits)
  );
  AluReg f_3 ( // @[TensorAlu.scala 84:36]
    .clock(f_3_clock),
    .io_opcode(f_3_io_opcode),
    .io_a_valid(f_3_io_a_valid),
    .io_a_bits(f_3_io_a_bits),
    .io_b_valid(f_3_io_b_valid),
    .io_b_bits(f_3_io_b_bits),
    .io_y_valid(f_3_io_y_valid),
    .io_y_bits(f_3_io_y_bits)
  );
  AluReg f_4 ( // @[TensorAlu.scala 84:36]
    .clock(f_4_clock),
    .io_opcode(f_4_io_opcode),
    .io_a_valid(f_4_io_a_valid),
    .io_a_bits(f_4_io_a_bits),
    .io_b_valid(f_4_io_b_valid),
    .io_b_bits(f_4_io_b_bits),
    .io_y_valid(f_4_io_y_valid),
    .io_y_bits(f_4_io_y_bits)
  );
  AluReg f_5 ( // @[TensorAlu.scala 84:36]
    .clock(f_5_clock),
    .io_opcode(f_5_io_opcode),
    .io_a_valid(f_5_io_a_valid),
    .io_a_bits(f_5_io_a_bits),
    .io_b_valid(f_5_io_b_valid),
    .io_b_bits(f_5_io_b_bits),
    .io_y_valid(f_5_io_y_valid),
    .io_y_bits(f_5_io_y_bits)
  );
  AluReg f_6 ( // @[TensorAlu.scala 84:36]
    .clock(f_6_clock),
    .io_opcode(f_6_io_opcode),
    .io_a_valid(f_6_io_a_valid),
    .io_a_bits(f_6_io_a_bits),
    .io_b_valid(f_6_io_b_valid),
    .io_b_bits(f_6_io_b_bits),
    .io_y_valid(f_6_io_y_valid),
    .io_y_bits(f_6_io_y_bits)
  );
  AluReg f_7 ( // @[TensorAlu.scala 84:36]
    .clock(f_7_clock),
    .io_opcode(f_7_io_opcode),
    .io_a_valid(f_7_io_a_valid),
    .io_a_bits(f_7_io_a_bits),
    .io_b_valid(f_7_io_b_valid),
    .io_b_bits(f_7_io_b_bits),
    .io_y_valid(f_7_io_y_valid),
    .io_y_bits(f_7_io_y_bits)
  );
  AluReg f_8 ( // @[TensorAlu.scala 84:36]
    .clock(f_8_clock),
    .io_opcode(f_8_io_opcode),
    .io_a_valid(f_8_io_a_valid),
    .io_a_bits(f_8_io_a_bits),
    .io_b_valid(f_8_io_b_valid),
    .io_b_bits(f_8_io_b_bits),
    .io_y_valid(f_8_io_y_valid),
    .io_y_bits(f_8_io_y_bits)
  );
  AluReg f_9 ( // @[TensorAlu.scala 84:36]
    .clock(f_9_clock),
    .io_opcode(f_9_io_opcode),
    .io_a_valid(f_9_io_a_valid),
    .io_a_bits(f_9_io_a_bits),
    .io_b_valid(f_9_io_b_valid),
    .io_b_bits(f_9_io_b_bits),
    .io_y_valid(f_9_io_y_valid),
    .io_y_bits(f_9_io_y_bits)
  );
  AluReg f_10 ( // @[TensorAlu.scala 84:36]
    .clock(f_10_clock),
    .io_opcode(f_10_io_opcode),
    .io_a_valid(f_10_io_a_valid),
    .io_a_bits(f_10_io_a_bits),
    .io_b_valid(f_10_io_b_valid),
    .io_b_bits(f_10_io_b_bits),
    .io_y_valid(f_10_io_y_valid),
    .io_y_bits(f_10_io_y_bits)
  );
  AluReg f_11 ( // @[TensorAlu.scala 84:36]
    .clock(f_11_clock),
    .io_opcode(f_11_io_opcode),
    .io_a_valid(f_11_io_a_valid),
    .io_a_bits(f_11_io_a_bits),
    .io_b_valid(f_11_io_b_valid),
    .io_b_bits(f_11_io_b_bits),
    .io_y_valid(f_11_io_y_valid),
    .io_y_bits(f_11_io_y_bits)
  );
  AluReg f_12 ( // @[TensorAlu.scala 84:36]
    .clock(f_12_clock),
    .io_opcode(f_12_io_opcode),
    .io_a_valid(f_12_io_a_valid),
    .io_a_bits(f_12_io_a_bits),
    .io_b_valid(f_12_io_b_valid),
    .io_b_bits(f_12_io_b_bits),
    .io_y_valid(f_12_io_y_valid),
    .io_y_bits(f_12_io_y_bits)
  );
  AluReg f_13 ( // @[TensorAlu.scala 84:36]
    .clock(f_13_clock),
    .io_opcode(f_13_io_opcode),
    .io_a_valid(f_13_io_a_valid),
    .io_a_bits(f_13_io_a_bits),
    .io_b_valid(f_13_io_b_valid),
    .io_b_bits(f_13_io_b_bits),
    .io_y_valid(f_13_io_y_valid),
    .io_y_bits(f_13_io_y_bits)
  );
  AluReg f_14 ( // @[TensorAlu.scala 84:36]
    .clock(f_14_clock),
    .io_opcode(f_14_io_opcode),
    .io_a_valid(f_14_io_a_valid),
    .io_a_bits(f_14_io_a_bits),
    .io_b_valid(f_14_io_b_valid),
    .io_b_bits(f_14_io_b_bits),
    .io_y_valid(f_14_io_y_valid),
    .io_y_bits(f_14_io_y_bits)
  );
  AluReg f_15 ( // @[TensorAlu.scala 84:36]
    .clock(f_15_clock),
    .io_opcode(f_15_io_opcode),
    .io_a_valid(f_15_io_a_valid),
    .io_a_bits(f_15_io_a_bits),
    .io_b_valid(f_15_io_b_valid),
    .io_b_bits(f_15_io_b_bits),
    .io_y_valid(f_15_io_y_valid),
    .io_y_bits(f_15_io_y_bits)
  );
  AluReg f_16 ( // @[TensorAlu.scala 84:36]
    .clock(f_16_clock),
    .io_opcode(f_16_io_opcode),
    .io_a_valid(f_16_io_a_valid),
    .io_a_bits(f_16_io_a_bits),
    .io_b_valid(f_16_io_b_valid),
    .io_b_bits(f_16_io_b_bits),
    .io_y_valid(f_16_io_y_valid),
    .io_y_bits(f_16_io_y_bits)
  );
  AluReg f_17 ( // @[TensorAlu.scala 84:36]
    .clock(f_17_clock),
    .io_opcode(f_17_io_opcode),
    .io_a_valid(f_17_io_a_valid),
    .io_a_bits(f_17_io_a_bits),
    .io_b_valid(f_17_io_b_valid),
    .io_b_bits(f_17_io_b_bits),
    .io_y_valid(f_17_io_y_valid),
    .io_y_bits(f_17_io_y_bits)
  );
  AluReg f_18 ( // @[TensorAlu.scala 84:36]
    .clock(f_18_clock),
    .io_opcode(f_18_io_opcode),
    .io_a_valid(f_18_io_a_valid),
    .io_a_bits(f_18_io_a_bits),
    .io_b_valid(f_18_io_b_valid),
    .io_b_bits(f_18_io_b_bits),
    .io_y_valid(f_18_io_y_valid),
    .io_y_bits(f_18_io_y_bits)
  );
  AluReg f_19 ( // @[TensorAlu.scala 84:36]
    .clock(f_19_clock),
    .io_opcode(f_19_io_opcode),
    .io_a_valid(f_19_io_a_valid),
    .io_a_bits(f_19_io_a_bits),
    .io_b_valid(f_19_io_b_valid),
    .io_b_bits(f_19_io_b_bits),
    .io_y_valid(f_19_io_y_valid),
    .io_y_bits(f_19_io_y_bits)
  );
  AluReg f_20 ( // @[TensorAlu.scala 84:36]
    .clock(f_20_clock),
    .io_opcode(f_20_io_opcode),
    .io_a_valid(f_20_io_a_valid),
    .io_a_bits(f_20_io_a_bits),
    .io_b_valid(f_20_io_b_valid),
    .io_b_bits(f_20_io_b_bits),
    .io_y_valid(f_20_io_y_valid),
    .io_y_bits(f_20_io_y_bits)
  );
  AluReg f_21 ( // @[TensorAlu.scala 84:36]
    .clock(f_21_clock),
    .io_opcode(f_21_io_opcode),
    .io_a_valid(f_21_io_a_valid),
    .io_a_bits(f_21_io_a_bits),
    .io_b_valid(f_21_io_b_valid),
    .io_b_bits(f_21_io_b_bits),
    .io_y_valid(f_21_io_y_valid),
    .io_y_bits(f_21_io_y_bits)
  );
  AluReg f_22 ( // @[TensorAlu.scala 84:36]
    .clock(f_22_clock),
    .io_opcode(f_22_io_opcode),
    .io_a_valid(f_22_io_a_valid),
    .io_a_bits(f_22_io_a_bits),
    .io_b_valid(f_22_io_b_valid),
    .io_b_bits(f_22_io_b_bits),
    .io_y_valid(f_22_io_y_valid),
    .io_y_bits(f_22_io_y_bits)
  );
  AluReg f_23 ( // @[TensorAlu.scala 84:36]
    .clock(f_23_clock),
    .io_opcode(f_23_io_opcode),
    .io_a_valid(f_23_io_a_valid),
    .io_a_bits(f_23_io_a_bits),
    .io_b_valid(f_23_io_b_valid),
    .io_b_bits(f_23_io_b_bits),
    .io_y_valid(f_23_io_y_valid),
    .io_y_bits(f_23_io_y_bits)
  );
  AluReg f_24 ( // @[TensorAlu.scala 84:36]
    .clock(f_24_clock),
    .io_opcode(f_24_io_opcode),
    .io_a_valid(f_24_io_a_valid),
    .io_a_bits(f_24_io_a_bits),
    .io_b_valid(f_24_io_b_valid),
    .io_b_bits(f_24_io_b_bits),
    .io_y_valid(f_24_io_y_valid),
    .io_y_bits(f_24_io_y_bits)
  );
  AluReg f_25 ( // @[TensorAlu.scala 84:36]
    .clock(f_25_clock),
    .io_opcode(f_25_io_opcode),
    .io_a_valid(f_25_io_a_valid),
    .io_a_bits(f_25_io_a_bits),
    .io_b_valid(f_25_io_b_valid),
    .io_b_bits(f_25_io_b_bits),
    .io_y_valid(f_25_io_y_valid),
    .io_y_bits(f_25_io_y_bits)
  );
  AluReg f_26 ( // @[TensorAlu.scala 84:36]
    .clock(f_26_clock),
    .io_opcode(f_26_io_opcode),
    .io_a_valid(f_26_io_a_valid),
    .io_a_bits(f_26_io_a_bits),
    .io_b_valid(f_26_io_b_valid),
    .io_b_bits(f_26_io_b_bits),
    .io_y_valid(f_26_io_y_valid),
    .io_y_bits(f_26_io_y_bits)
  );
  AluReg f_27 ( // @[TensorAlu.scala 84:36]
    .clock(f_27_clock),
    .io_opcode(f_27_io_opcode),
    .io_a_valid(f_27_io_a_valid),
    .io_a_bits(f_27_io_a_bits),
    .io_b_valid(f_27_io_b_valid),
    .io_b_bits(f_27_io_b_bits),
    .io_y_valid(f_27_io_y_valid),
    .io_y_bits(f_27_io_y_bits)
  );
  AluReg f_28 ( // @[TensorAlu.scala 84:36]
    .clock(f_28_clock),
    .io_opcode(f_28_io_opcode),
    .io_a_valid(f_28_io_a_valid),
    .io_a_bits(f_28_io_a_bits),
    .io_b_valid(f_28_io_b_valid),
    .io_b_bits(f_28_io_b_bits),
    .io_y_valid(f_28_io_y_valid),
    .io_y_bits(f_28_io_y_bits)
  );
  AluReg f_29 ( // @[TensorAlu.scala 84:36]
    .clock(f_29_clock),
    .io_opcode(f_29_io_opcode),
    .io_a_valid(f_29_io_a_valid),
    .io_a_bits(f_29_io_a_bits),
    .io_b_valid(f_29_io_b_valid),
    .io_b_bits(f_29_io_b_bits),
    .io_y_valid(f_29_io_y_valid),
    .io_y_bits(f_29_io_y_bits)
  );
  AluReg f_30 ( // @[TensorAlu.scala 84:36]
    .clock(f_30_clock),
    .io_opcode(f_30_io_opcode),
    .io_a_valid(f_30_io_a_valid),
    .io_a_bits(f_30_io_a_bits),
    .io_b_valid(f_30_io_b_valid),
    .io_b_bits(f_30_io_b_bits),
    .io_y_valid(f_30_io_y_valid),
    .io_y_bits(f_30_io_y_bits)
  );
  AluReg f_31 ( // @[TensorAlu.scala 84:36]
    .clock(f_31_clock),
    .io_opcode(f_31_io_opcode),
    .io_a_valid(f_31_io_a_valid),
    .io_a_bits(f_31_io_a_bits),
    .io_b_valid(f_31_io_b_valid),
    .io_b_bits(f_31_io_b_bits),
    .io_y_valid(f_31_io_y_valid),
    .io_y_bits(f_31_io_y_bits)
  );
  assign io_acc_y_data_valid = &_io_acc_y_data_valid_T; // @[TensorAlu.scala 96:39]
  assign io_acc_y_data_bits_0_0 = f_0_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_1 = f_1_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_2 = f_2_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_3 = f_3_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_4 = f_4_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_5 = f_5_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_6 = f_6_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_7 = f_7_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_8 = f_8_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_9 = f_9_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_10 = f_10_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_11 = f_11_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_12 = f_12_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_13 = f_13_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_14 = f_14_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_15 = f_15_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_16 = f_16_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_17 = f_17_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_18 = f_18_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_19 = f_19_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_20 = f_20_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_21 = f_21_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_22 = f_22_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_23 = f_23_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_24 = f_24_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_25 = f_25_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_26 = f_26_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_27 = f_27_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_28 = f_28_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_29 = f_29_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_30 = f_30_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_acc_y_data_bits_0_31 = f_31_io_y_bits; // @[TensorAlu.scala 93:30]
  assign io_out_data_valid = &_io_acc_y_data_valid_T; // @[TensorAlu.scala 97:37]
  assign io_out_data_bits_0_0 = f_0_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_1 = f_1_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_2 = f_2_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_3 = f_3_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_4 = f_4_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_5 = f_5_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_6 = f_6_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_7 = f_7_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_8 = f_8_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_9 = f_9_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_10 = f_10_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_11 = f_11_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_12 = f_12_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_13 = f_13_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_14 = f_14_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_15 = f_15_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_16 = f_16_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_17 = f_17_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_18 = f_18_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_19 = f_19_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_20 = f_20_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_21 = f_21_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_22 = f_22_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_23 = f_23_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_24 = f_24_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_25 = f_25_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_26 = f_26_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_27 = f_27_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_28 = f_28_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_29 = f_29_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_30 = f_30_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign io_out_data_bits_0_31 = f_31_io_y_bits[7:0]; // @[TensorAlu.scala 94:28]
  assign f_0_clock = clock;
  assign f_0_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_0_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_0_io_a_bits = io_acc_a_data_bits_0_0; // @[TensorAlu.scala 89:20]
  assign f_0_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_0_io_b_bits = io_acc_b_data_bits_0_0; // @[TensorAlu.scala 91:20]
  assign f_1_clock = clock;
  assign f_1_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_1_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_1_io_a_bits = io_acc_a_data_bits_0_1; // @[TensorAlu.scala 89:20]
  assign f_1_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_1_io_b_bits = io_acc_b_data_bits_0_1; // @[TensorAlu.scala 91:20]
  assign f_2_clock = clock;
  assign f_2_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_2_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_2_io_a_bits = io_acc_a_data_bits_0_2; // @[TensorAlu.scala 89:20]
  assign f_2_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_2_io_b_bits = io_acc_b_data_bits_0_2; // @[TensorAlu.scala 91:20]
  assign f_3_clock = clock;
  assign f_3_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_3_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_3_io_a_bits = io_acc_a_data_bits_0_3; // @[TensorAlu.scala 89:20]
  assign f_3_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_3_io_b_bits = io_acc_b_data_bits_0_3; // @[TensorAlu.scala 91:20]
  assign f_4_clock = clock;
  assign f_4_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_4_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_4_io_a_bits = io_acc_a_data_bits_0_4; // @[TensorAlu.scala 89:20]
  assign f_4_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_4_io_b_bits = io_acc_b_data_bits_0_4; // @[TensorAlu.scala 91:20]
  assign f_5_clock = clock;
  assign f_5_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_5_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_5_io_a_bits = io_acc_a_data_bits_0_5; // @[TensorAlu.scala 89:20]
  assign f_5_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_5_io_b_bits = io_acc_b_data_bits_0_5; // @[TensorAlu.scala 91:20]
  assign f_6_clock = clock;
  assign f_6_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_6_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_6_io_a_bits = io_acc_a_data_bits_0_6; // @[TensorAlu.scala 89:20]
  assign f_6_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_6_io_b_bits = io_acc_b_data_bits_0_6; // @[TensorAlu.scala 91:20]
  assign f_7_clock = clock;
  assign f_7_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_7_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_7_io_a_bits = io_acc_a_data_bits_0_7; // @[TensorAlu.scala 89:20]
  assign f_7_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_7_io_b_bits = io_acc_b_data_bits_0_7; // @[TensorAlu.scala 91:20]
  assign f_8_clock = clock;
  assign f_8_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_8_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_8_io_a_bits = io_acc_a_data_bits_0_8; // @[TensorAlu.scala 89:20]
  assign f_8_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_8_io_b_bits = io_acc_b_data_bits_0_8; // @[TensorAlu.scala 91:20]
  assign f_9_clock = clock;
  assign f_9_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_9_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_9_io_a_bits = io_acc_a_data_bits_0_9; // @[TensorAlu.scala 89:20]
  assign f_9_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_9_io_b_bits = io_acc_b_data_bits_0_9; // @[TensorAlu.scala 91:20]
  assign f_10_clock = clock;
  assign f_10_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_10_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_10_io_a_bits = io_acc_a_data_bits_0_10; // @[TensorAlu.scala 89:20]
  assign f_10_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_10_io_b_bits = io_acc_b_data_bits_0_10; // @[TensorAlu.scala 91:20]
  assign f_11_clock = clock;
  assign f_11_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_11_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_11_io_a_bits = io_acc_a_data_bits_0_11; // @[TensorAlu.scala 89:20]
  assign f_11_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_11_io_b_bits = io_acc_b_data_bits_0_11; // @[TensorAlu.scala 91:20]
  assign f_12_clock = clock;
  assign f_12_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_12_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_12_io_a_bits = io_acc_a_data_bits_0_12; // @[TensorAlu.scala 89:20]
  assign f_12_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_12_io_b_bits = io_acc_b_data_bits_0_12; // @[TensorAlu.scala 91:20]
  assign f_13_clock = clock;
  assign f_13_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_13_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_13_io_a_bits = io_acc_a_data_bits_0_13; // @[TensorAlu.scala 89:20]
  assign f_13_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_13_io_b_bits = io_acc_b_data_bits_0_13; // @[TensorAlu.scala 91:20]
  assign f_14_clock = clock;
  assign f_14_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_14_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_14_io_a_bits = io_acc_a_data_bits_0_14; // @[TensorAlu.scala 89:20]
  assign f_14_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_14_io_b_bits = io_acc_b_data_bits_0_14; // @[TensorAlu.scala 91:20]
  assign f_15_clock = clock;
  assign f_15_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_15_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_15_io_a_bits = io_acc_a_data_bits_0_15; // @[TensorAlu.scala 89:20]
  assign f_15_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_15_io_b_bits = io_acc_b_data_bits_0_15; // @[TensorAlu.scala 91:20]
  assign f_16_clock = clock;
  assign f_16_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_16_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_16_io_a_bits = io_acc_a_data_bits_0_16; // @[TensorAlu.scala 89:20]
  assign f_16_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_16_io_b_bits = io_acc_b_data_bits_0_16; // @[TensorAlu.scala 91:20]
  assign f_17_clock = clock;
  assign f_17_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_17_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_17_io_a_bits = io_acc_a_data_bits_0_17; // @[TensorAlu.scala 89:20]
  assign f_17_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_17_io_b_bits = io_acc_b_data_bits_0_17; // @[TensorAlu.scala 91:20]
  assign f_18_clock = clock;
  assign f_18_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_18_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_18_io_a_bits = io_acc_a_data_bits_0_18; // @[TensorAlu.scala 89:20]
  assign f_18_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_18_io_b_bits = io_acc_b_data_bits_0_18; // @[TensorAlu.scala 91:20]
  assign f_19_clock = clock;
  assign f_19_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_19_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_19_io_a_bits = io_acc_a_data_bits_0_19; // @[TensorAlu.scala 89:20]
  assign f_19_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_19_io_b_bits = io_acc_b_data_bits_0_19; // @[TensorAlu.scala 91:20]
  assign f_20_clock = clock;
  assign f_20_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_20_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_20_io_a_bits = io_acc_a_data_bits_0_20; // @[TensorAlu.scala 89:20]
  assign f_20_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_20_io_b_bits = io_acc_b_data_bits_0_20; // @[TensorAlu.scala 91:20]
  assign f_21_clock = clock;
  assign f_21_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_21_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_21_io_a_bits = io_acc_a_data_bits_0_21; // @[TensorAlu.scala 89:20]
  assign f_21_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_21_io_b_bits = io_acc_b_data_bits_0_21; // @[TensorAlu.scala 91:20]
  assign f_22_clock = clock;
  assign f_22_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_22_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_22_io_a_bits = io_acc_a_data_bits_0_22; // @[TensorAlu.scala 89:20]
  assign f_22_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_22_io_b_bits = io_acc_b_data_bits_0_22; // @[TensorAlu.scala 91:20]
  assign f_23_clock = clock;
  assign f_23_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_23_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_23_io_a_bits = io_acc_a_data_bits_0_23; // @[TensorAlu.scala 89:20]
  assign f_23_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_23_io_b_bits = io_acc_b_data_bits_0_23; // @[TensorAlu.scala 91:20]
  assign f_24_clock = clock;
  assign f_24_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_24_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_24_io_a_bits = io_acc_a_data_bits_0_24; // @[TensorAlu.scala 89:20]
  assign f_24_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_24_io_b_bits = io_acc_b_data_bits_0_24; // @[TensorAlu.scala 91:20]
  assign f_25_clock = clock;
  assign f_25_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_25_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_25_io_a_bits = io_acc_a_data_bits_0_25; // @[TensorAlu.scala 89:20]
  assign f_25_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_25_io_b_bits = io_acc_b_data_bits_0_25; // @[TensorAlu.scala 91:20]
  assign f_26_clock = clock;
  assign f_26_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_26_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_26_io_a_bits = io_acc_a_data_bits_0_26; // @[TensorAlu.scala 89:20]
  assign f_26_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_26_io_b_bits = io_acc_b_data_bits_0_26; // @[TensorAlu.scala 91:20]
  assign f_27_clock = clock;
  assign f_27_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_27_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_27_io_a_bits = io_acc_a_data_bits_0_27; // @[TensorAlu.scala 89:20]
  assign f_27_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_27_io_b_bits = io_acc_b_data_bits_0_27; // @[TensorAlu.scala 91:20]
  assign f_28_clock = clock;
  assign f_28_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_28_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_28_io_a_bits = io_acc_a_data_bits_0_28; // @[TensorAlu.scala 89:20]
  assign f_28_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_28_io_b_bits = io_acc_b_data_bits_0_28; // @[TensorAlu.scala 91:20]
  assign f_29_clock = clock;
  assign f_29_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_29_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_29_io_a_bits = io_acc_a_data_bits_0_29; // @[TensorAlu.scala 89:20]
  assign f_29_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_29_io_b_bits = io_acc_b_data_bits_0_29; // @[TensorAlu.scala 91:20]
  assign f_30_clock = clock;
  assign f_30_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_30_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_30_io_a_bits = io_acc_a_data_bits_0_30; // @[TensorAlu.scala 89:20]
  assign f_30_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_30_io_b_bits = io_acc_b_data_bits_0_30; // @[TensorAlu.scala 91:20]
  assign f_31_clock = clock;
  assign f_31_io_opcode = io_opcode; // @[TensorAlu.scala 87:20]
  assign f_31_io_a_valid = io_acc_a_data_valid; // @[TensorAlu.scala 88:21]
  assign f_31_io_a_bits = io_acc_a_data_bits_0_31; // @[TensorAlu.scala 89:20]
  assign f_31_io_b_valid = io_acc_b_data_valid; // @[TensorAlu.scala 90:21]
  assign f_31_io_b_bits = io_acc_b_data_bits_0_31; // @[TensorAlu.scala 91:20]
endmodule
module TensorAlu(
  input         clock,
  input         reset,
  input         io_start,
  output        io_done,
  input  [15:0] io_dec_alu_imm,
  input         io_dec_alu_use_imm,
  input  [2:0]  io_dec_alu_op,
  input  [10:0] io_dec_src_1,
  input  [10:0] io_dec_src_0,
  input  [10:0] io_dec_dst_1,
  input  [10:0] io_dec_dst_0,
  input  [13:0] io_dec_lp_1,
  input  [13:0] io_dec_lp_0,
  input  [13:0] io_dec_uop_end,
  input  [12:0] io_dec_uop_begin,
  output        io_uop_idx_valid,
  output [6:0]  io_uop_idx_bits,
  input  [9:0]  io_uop_data_bits_u2,
  input  [10:0] io_uop_data_bits_u1,
  input  [10:0] io_uop_data_bits_u0,
  output        io_acc_rd_0_idx_valid,
  output [6:0]  io_acc_rd_0_idx_bits,
  input         io_acc_rd_0_data_valid,
  input  [31:0] io_acc_rd_0_data_bits_0_0,
  input  [31:0] io_acc_rd_0_data_bits_0_1,
  input  [31:0] io_acc_rd_0_data_bits_0_2,
  input  [31:0] io_acc_rd_0_data_bits_0_3,
  input  [31:0] io_acc_rd_0_data_bits_0_4,
  input  [31:0] io_acc_rd_0_data_bits_0_5,
  input  [31:0] io_acc_rd_0_data_bits_0_6,
  input  [31:0] io_acc_rd_0_data_bits_0_7,
  input  [31:0] io_acc_rd_0_data_bits_0_8,
  input  [31:0] io_acc_rd_0_data_bits_0_9,
  input  [31:0] io_acc_rd_0_data_bits_0_10,
  input  [31:0] io_acc_rd_0_data_bits_0_11,
  input  [31:0] io_acc_rd_0_data_bits_0_12,
  input  [31:0] io_acc_rd_0_data_bits_0_13,
  input  [31:0] io_acc_rd_0_data_bits_0_14,
  input  [31:0] io_acc_rd_0_data_bits_0_15,
  input  [31:0] io_acc_rd_0_data_bits_0_16,
  input  [31:0] io_acc_rd_0_data_bits_0_17,
  input  [31:0] io_acc_rd_0_data_bits_0_18,
  input  [31:0] io_acc_rd_0_data_bits_0_19,
  input  [31:0] io_acc_rd_0_data_bits_0_20,
  input  [31:0] io_acc_rd_0_data_bits_0_21,
  input  [31:0] io_acc_rd_0_data_bits_0_22,
  input  [31:0] io_acc_rd_0_data_bits_0_23,
  input  [31:0] io_acc_rd_0_data_bits_0_24,
  input  [31:0] io_acc_rd_0_data_bits_0_25,
  input  [31:0] io_acc_rd_0_data_bits_0_26,
  input  [31:0] io_acc_rd_0_data_bits_0_27,
  input  [31:0] io_acc_rd_0_data_bits_0_28,
  input  [31:0] io_acc_rd_0_data_bits_0_29,
  input  [31:0] io_acc_rd_0_data_bits_0_30,
  input  [31:0] io_acc_rd_0_data_bits_0_31,
  output        io_acc_wr_0_valid,
  output [6:0]  io_acc_wr_0_bits_idx,
  output [31:0] io_acc_wr_0_bits_data_0_0,
  output [31:0] io_acc_wr_0_bits_data_0_1,
  output [31:0] io_acc_wr_0_bits_data_0_2,
  output [31:0] io_acc_wr_0_bits_data_0_3,
  output [31:0] io_acc_wr_0_bits_data_0_4,
  output [31:0] io_acc_wr_0_bits_data_0_5,
  output [31:0] io_acc_wr_0_bits_data_0_6,
  output [31:0] io_acc_wr_0_bits_data_0_7,
  output [31:0] io_acc_wr_0_bits_data_0_8,
  output [31:0] io_acc_wr_0_bits_data_0_9,
  output [31:0] io_acc_wr_0_bits_data_0_10,
  output [31:0] io_acc_wr_0_bits_data_0_11,
  output [31:0] io_acc_wr_0_bits_data_0_12,
  output [31:0] io_acc_wr_0_bits_data_0_13,
  output [31:0] io_acc_wr_0_bits_data_0_14,
  output [31:0] io_acc_wr_0_bits_data_0_15,
  output [31:0] io_acc_wr_0_bits_data_0_16,
  output [31:0] io_acc_wr_0_bits_data_0_17,
  output [31:0] io_acc_wr_0_bits_data_0_18,
  output [31:0] io_acc_wr_0_bits_data_0_19,
  output [31:0] io_acc_wr_0_bits_data_0_20,
  output [31:0] io_acc_wr_0_bits_data_0_21,
  output [31:0] io_acc_wr_0_bits_data_0_22,
  output [31:0] io_acc_wr_0_bits_data_0_23,
  output [31:0] io_acc_wr_0_bits_data_0_24,
  output [31:0] io_acc_wr_0_bits_data_0_25,
  output [31:0] io_acc_wr_0_bits_data_0_26,
  output [31:0] io_acc_wr_0_bits_data_0_27,
  output [31:0] io_acc_wr_0_bits_data_0_28,
  output [31:0] io_acc_wr_0_bits_data_0_29,
  output [31:0] io_acc_wr_0_bits_data_0_30,
  output [31:0] io_acc_wr_0_bits_data_0_31,
  input         io_out_rd_0_data_valid,
  output        io_out_wr_0_valid,
  output [6:0]  io_out_wr_0_bits_idx,
  output [7:0]  io_out_wr_0_bits_data_0_0,
  output [7:0]  io_out_wr_0_bits_data_0_1,
  output [7:0]  io_out_wr_0_bits_data_0_2,
  output [7:0]  io_out_wr_0_bits_data_0_3,
  output [7:0]  io_out_wr_0_bits_data_0_4,
  output [7:0]  io_out_wr_0_bits_data_0_5,
  output [7:0]  io_out_wr_0_bits_data_0_6,
  output [7:0]  io_out_wr_0_bits_data_0_7,
  output [7:0]  io_out_wr_0_bits_data_0_8,
  output [7:0]  io_out_wr_0_bits_data_0_9,
  output [7:0]  io_out_wr_0_bits_data_0_10,
  output [7:0]  io_out_wr_0_bits_data_0_11,
  output [7:0]  io_out_wr_0_bits_data_0_12,
  output [7:0]  io_out_wr_0_bits_data_0_13,
  output [7:0]  io_out_wr_0_bits_data_0_14,
  output [7:0]  io_out_wr_0_bits_data_0_15,
  output [7:0]  io_out_wr_0_bits_data_0_16,
  output [7:0]  io_out_wr_0_bits_data_0_17,
  output [7:0]  io_out_wr_0_bits_data_0_18,
  output [7:0]  io_out_wr_0_bits_data_0_19,
  output [7:0]  io_out_wr_0_bits_data_0_20,
  output [7:0]  io_out_wr_0_bits_data_0_21,
  output [7:0]  io_out_wr_0_bits_data_0_22,
  output [7:0]  io_out_wr_0_bits_data_0_23,
  output [7:0]  io_out_wr_0_bits_data_0_24,
  output [7:0]  io_out_wr_0_bits_data_0_25,
  output [7:0]  io_out_wr_0_bits_data_0_26,
  output [7:0]  io_out_wr_0_bits_data_0_27,
  output [7:0]  io_out_wr_0_bits_data_0_28,
  output [7:0]  io_out_wr_0_bits_data_0_29,
  output [7:0]  io_out_wr_0_bits_data_0_30,
  output [7:0]  io_out_wr_0_bits_data_0_31
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
`endif // RANDOMIZE_REG_INIT
  wire  index_generator_clock; // @[TensorAlu.scala 205:31]
  wire  index_generator_reset; // @[TensorAlu.scala 205:31]
  wire  index_generator_io_start; // @[TensorAlu.scala 205:31]
  wire  index_generator_io_last; // @[TensorAlu.scala 205:31]
  wire  index_generator_io_dec_alu_use_imm; // @[TensorAlu.scala 205:31]
  wire [10:0] index_generator_io_dec_src_1; // @[TensorAlu.scala 205:31]
  wire [10:0] index_generator_io_dec_src_0; // @[TensorAlu.scala 205:31]
  wire [10:0] index_generator_io_dec_dst_1; // @[TensorAlu.scala 205:31]
  wire [10:0] index_generator_io_dec_dst_0; // @[TensorAlu.scala 205:31]
  wire [13:0] index_generator_io_dec_lp_1; // @[TensorAlu.scala 205:31]
  wire [13:0] index_generator_io_dec_lp_0; // @[TensorAlu.scala 205:31]
  wire [13:0] index_generator_io_dec_uop_end; // @[TensorAlu.scala 205:31]
  wire [12:0] index_generator_io_dec_uop_begin; // @[TensorAlu.scala 205:31]
  wire  index_generator_io_valid; // @[TensorAlu.scala 205:31]
  wire  index_generator_io_src_valid; // @[TensorAlu.scala 205:31]
  wire [6:0] index_generator_io_dst_idx; // @[TensorAlu.scala 205:31]
  wire [6:0] index_generator_io_src_idx; // @[TensorAlu.scala 205:31]
  wire [6:0] index_generator_io_uop_idx; // @[TensorAlu.scala 205:31]
  wire  alu_clock; // @[TensorAlu.scala 301:21]
  wire [2:0] alu_io_opcode; // @[TensorAlu.scala 301:21]
  wire  alu_io_acc_a_data_valid; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_0; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_1; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_2; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_3; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_4; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_5; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_6; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_7; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_8; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_9; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_10; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_11; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_12; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_13; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_14; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_15; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_16; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_17; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_18; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_19; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_20; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_21; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_22; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_23; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_24; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_25; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_26; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_27; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_28; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_29; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_30; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_a_data_bits_0_31; // @[TensorAlu.scala 301:21]
  wire  alu_io_acc_b_data_valid; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_0; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_1; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_2; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_3; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_4; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_5; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_6; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_7; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_8; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_9; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_10; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_11; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_12; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_13; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_14; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_15; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_16; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_17; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_18; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_19; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_20; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_21; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_22; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_23; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_24; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_25; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_26; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_27; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_28; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_29; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_30; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_b_data_bits_0_31; // @[TensorAlu.scala 301:21]
  wire  alu_io_acc_y_data_valid; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_0; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_1; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_2; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_3; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_4; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_5; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_6; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_7; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_8; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_9; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_10; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_11; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_12; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_13; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_14; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_15; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_16; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_17; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_18; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_19; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_20; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_21; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_22; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_23; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_24; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_25; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_26; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_27; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_28; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_29; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_30; // @[TensorAlu.scala 301:21]
  wire [31:0] alu_io_acc_y_data_bits_0_31; // @[TensorAlu.scala 301:21]
  wire  alu_io_out_data_valid; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_0; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_1; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_2; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_3; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_4; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_5; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_6; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_7; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_8; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_9; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_10; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_11; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_12; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_13; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_14; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_15; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_16; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_17; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_18; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_19; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_20; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_21; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_22; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_23; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_24; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_25; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_26; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_27; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_28; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_29; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_30; // @[TensorAlu.scala 301:21]
  wire [7:0] alu_io_out_data_bits_0_31; // @[TensorAlu.scala 301:21]
  reg [1:0] state; // @[TensorAlu.scala 202:22]
  reg [3:0] inflight; // @[TensorAlu.scala 203:25]
  wire  _T = state == 2'h0; // @[TensorAlu.scala 210:14]
  wire  _T_5 = inflight == 4'h0; // @[TensorAlu.scala 214:42]
  wire  _T_6 = state == 2'h2 & inflight == 4'h0; // @[TensorAlu.scala 214:30]
  wire  _GEN_3 = state == 2'h1 & index_generator_io_last ? 1'h0 : _T_6; // @[TensorAlu.scala 209:11 212:57]
  reg  valid_r1; // @[Reg.scala 28:20]
  wire  _GEN_6 = index_generator_io_valid; // @[Reg.scala 29:18 28:20 29:22]
  reg  valid_r2; // @[TensorAlu.scala 227:25]
  reg  valid_r3; // @[TensorAlu.scala 228:25]
  reg  valid_r4; // @[TensorAlu.scala 229:25]
  wire  _T_7 = index_generator_io_valid & valid_r4; // @[TensorAlu.scala 231:33]
  wire  _T_10 = ~reset; // @[TensorAlu.scala 233:11]
  wire [3:0] _inflight_T_1 = inflight + 4'h1; // @[TensorAlu.scala 234:26]
  wire [3:0] _inflight_T_3 = inflight - 4'h1; // @[TensorAlu.scala 237:26]
  wire [3:0] _GEN_7 = valid_r4 ? _inflight_T_3 : inflight; // @[TensorAlu.scala 235:24 237:14 203:25]
  reg  src_valid_r1; // @[Reg.scala 28:20]
  wire  _GEN_11 = index_generator_io_src_valid; // @[Reg.scala 29:18 28:20 29:22]
  reg  src_valid_r2; // @[TensorAlu.scala 248:29]
  reg  src_valid_r3; // @[TensorAlu.scala 249:29]
  reg [6:0] dst_idx_r1; // @[Reg.scala 16:16]
  reg [6:0] src_idx_r1; // @[Reg.scala 16:16]
  wire [10:0] u2 = {{1'd0}, io_uop_data_bits_u2}; // @[TensorAlu.scala 260:{40,40}]
  wire [17:0] _src_offset_T = {u2, 7'h0}; // @[TensorAlu.scala 263:24]
  wire [17:0] _GEN_14 = {{7'd0}, io_uop_data_bits_u1}; // @[TensorAlu.scala 263:30]
  wire [17:0] src_offset = _src_offset_T | _GEN_14; // @[TensorAlu.scala 263:30]
  reg  io_acc_rd_0_idx_valid_REG; // @[TensorAlu.scala 268:40]
  wire [17:0] _GEN_15 = {{11'd0}, src_idx_r1}; // @[TensorAlu.scala 271:35]
  wire [17:0] new_src_idx_r1 = _GEN_15 + src_offset; // @[TensorAlu.scala 271:35]
  reg [17:0] src_idx_r2; // @[TensorAlu.scala 272:27]
  reg [17:0] src_idx_r3; // @[TensorAlu.scala 273:27]
  wire [10:0] _GEN_16 = {{4'd0}, dst_idx_r1}; // @[TensorAlu.scala 275:35]
  wire [10:0] new_dst_idx_r1 = _GEN_16 + io_uop_data_bits_u0; // @[TensorAlu.scala 275:35]
  reg [10:0] dst_idx_r2; // @[TensorAlu.scala 276:27]
  reg [10:0] dst_idx_r3; // @[TensorAlu.scala 277:27]
  reg [10:0] dst_idx_r4; // @[TensorAlu.scala 278:27]
  reg [17:0] io_acc_rd_0_idx_bits_REG; // @[TensorAlu.scala 283:39]
  reg [31:0] save_src_0_0; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_1; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_2; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_3; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_4; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_5; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_6; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_7; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_8; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_9; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_10; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_11; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_12; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_13; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_14; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_15; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_16; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_17; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_18; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_19; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_20; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_21; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_22; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_23; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_24; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_25; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_26; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_27; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_28; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_29; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_30; // @[TensorAlu.scala 311:27]
  reg [31:0] save_src_0_31; // @[TensorAlu.scala 311:27]
  wire [31:0] _tensorImm_data_bits_0_0_T_1 = {16'hffff,io_dec_alu_imm}; // @[Cat.scala 31:58]
  wire [31:0] tensorImm_data_bits_0_0 = io_dec_alu_imm[15] ? _tensorImm_data_bits_0_0_T_1 : {{16'd0}, io_dec_alu_imm}; // @[TensorAlu.scala 319:17]
  wire  isSHR = io_dec_alu_op == 3'h3; // @[TensorAlu.scala 328:37]
  wire  neg_shift = isSHR & io_dec_alu_imm[15]; // @[TensorAlu.scala 329:27]
  reg  alu_io_acc_a_data_valid_REG; // @[TensorAlu.scala 338:39]
  wire  bypass_dst = valid_r3 & valid_r4 & dst_idx_r4 == dst_idx_r3; // @[TensorAlu.scala 386:41]
  wire [17:0] _GEN_17 = {{7'd0}, dst_idx_r4}; // @[TensorAlu.scala 387:60]
  wire  bypass_src = src_valid_r3 & valid_r4 & _GEN_17 == src_idx_r3; // @[TensorAlu.scala 387:45]
  wire  _GEN_18 = ~_T_7; // @[TensorAlu.scala 233:11]
  TensorAluIndexGenerator index_generator ( // @[TensorAlu.scala 205:31]
    .clock(index_generator_clock),
    .reset(index_generator_reset),
    .io_start(index_generator_io_start),
    .io_last(index_generator_io_last),
    .io_dec_alu_use_imm(index_generator_io_dec_alu_use_imm),
    .io_dec_src_1(index_generator_io_dec_src_1),
    .io_dec_src_0(index_generator_io_dec_src_0),
    .io_dec_dst_1(index_generator_io_dec_dst_1),
    .io_dec_dst_0(index_generator_io_dec_dst_0),
    .io_dec_lp_1(index_generator_io_dec_lp_1),
    .io_dec_lp_0(index_generator_io_dec_lp_0),
    .io_dec_uop_end(index_generator_io_dec_uop_end),
    .io_dec_uop_begin(index_generator_io_dec_uop_begin),
    .io_valid(index_generator_io_valid),
    .io_src_valid(index_generator_io_src_valid),
    .io_dst_idx(index_generator_io_dst_idx),
    .io_src_idx(index_generator_io_src_idx),
    .io_uop_idx(index_generator_io_uop_idx)
  );
  AluVector alu ( // @[TensorAlu.scala 301:21]
    .clock(alu_clock),
    .io_opcode(alu_io_opcode),
    .io_acc_a_data_valid(alu_io_acc_a_data_valid),
    .io_acc_a_data_bits_0_0(alu_io_acc_a_data_bits_0_0),
    .io_acc_a_data_bits_0_1(alu_io_acc_a_data_bits_0_1),
    .io_acc_a_data_bits_0_2(alu_io_acc_a_data_bits_0_2),
    .io_acc_a_data_bits_0_3(alu_io_acc_a_data_bits_0_3),
    .io_acc_a_data_bits_0_4(alu_io_acc_a_data_bits_0_4),
    .io_acc_a_data_bits_0_5(alu_io_acc_a_data_bits_0_5),
    .io_acc_a_data_bits_0_6(alu_io_acc_a_data_bits_0_6),
    .io_acc_a_data_bits_0_7(alu_io_acc_a_data_bits_0_7),
    .io_acc_a_data_bits_0_8(alu_io_acc_a_data_bits_0_8),
    .io_acc_a_data_bits_0_9(alu_io_acc_a_data_bits_0_9),
    .io_acc_a_data_bits_0_10(alu_io_acc_a_data_bits_0_10),
    .io_acc_a_data_bits_0_11(alu_io_acc_a_data_bits_0_11),
    .io_acc_a_data_bits_0_12(alu_io_acc_a_data_bits_0_12),
    .io_acc_a_data_bits_0_13(alu_io_acc_a_data_bits_0_13),
    .io_acc_a_data_bits_0_14(alu_io_acc_a_data_bits_0_14),
    .io_acc_a_data_bits_0_15(alu_io_acc_a_data_bits_0_15),
    .io_acc_a_data_bits_0_16(alu_io_acc_a_data_bits_0_16),
    .io_acc_a_data_bits_0_17(alu_io_acc_a_data_bits_0_17),
    .io_acc_a_data_bits_0_18(alu_io_acc_a_data_bits_0_18),
    .io_acc_a_data_bits_0_19(alu_io_acc_a_data_bits_0_19),
    .io_acc_a_data_bits_0_20(alu_io_acc_a_data_bits_0_20),
    .io_acc_a_data_bits_0_21(alu_io_acc_a_data_bits_0_21),
    .io_acc_a_data_bits_0_22(alu_io_acc_a_data_bits_0_22),
    .io_acc_a_data_bits_0_23(alu_io_acc_a_data_bits_0_23),
    .io_acc_a_data_bits_0_24(alu_io_acc_a_data_bits_0_24),
    .io_acc_a_data_bits_0_25(alu_io_acc_a_data_bits_0_25),
    .io_acc_a_data_bits_0_26(alu_io_acc_a_data_bits_0_26),
    .io_acc_a_data_bits_0_27(alu_io_acc_a_data_bits_0_27),
    .io_acc_a_data_bits_0_28(alu_io_acc_a_data_bits_0_28),
    .io_acc_a_data_bits_0_29(alu_io_acc_a_data_bits_0_29),
    .io_acc_a_data_bits_0_30(alu_io_acc_a_data_bits_0_30),
    .io_acc_a_data_bits_0_31(alu_io_acc_a_data_bits_0_31),
    .io_acc_b_data_valid(alu_io_acc_b_data_valid),
    .io_acc_b_data_bits_0_0(alu_io_acc_b_data_bits_0_0),
    .io_acc_b_data_bits_0_1(alu_io_acc_b_data_bits_0_1),
    .io_acc_b_data_bits_0_2(alu_io_acc_b_data_bits_0_2),
    .io_acc_b_data_bits_0_3(alu_io_acc_b_data_bits_0_3),
    .io_acc_b_data_bits_0_4(alu_io_acc_b_data_bits_0_4),
    .io_acc_b_data_bits_0_5(alu_io_acc_b_data_bits_0_5),
    .io_acc_b_data_bits_0_6(alu_io_acc_b_data_bits_0_6),
    .io_acc_b_data_bits_0_7(alu_io_acc_b_data_bits_0_7),
    .io_acc_b_data_bits_0_8(alu_io_acc_b_data_bits_0_8),
    .io_acc_b_data_bits_0_9(alu_io_acc_b_data_bits_0_9),
    .io_acc_b_data_bits_0_10(alu_io_acc_b_data_bits_0_10),
    .io_acc_b_data_bits_0_11(alu_io_acc_b_data_bits_0_11),
    .io_acc_b_data_bits_0_12(alu_io_acc_b_data_bits_0_12),
    .io_acc_b_data_bits_0_13(alu_io_acc_b_data_bits_0_13),
    .io_acc_b_data_bits_0_14(alu_io_acc_b_data_bits_0_14),
    .io_acc_b_data_bits_0_15(alu_io_acc_b_data_bits_0_15),
    .io_acc_b_data_bits_0_16(alu_io_acc_b_data_bits_0_16),
    .io_acc_b_data_bits_0_17(alu_io_acc_b_data_bits_0_17),
    .io_acc_b_data_bits_0_18(alu_io_acc_b_data_bits_0_18),
    .io_acc_b_data_bits_0_19(alu_io_acc_b_data_bits_0_19),
    .io_acc_b_data_bits_0_20(alu_io_acc_b_data_bits_0_20),
    .io_acc_b_data_bits_0_21(alu_io_acc_b_data_bits_0_21),
    .io_acc_b_data_bits_0_22(alu_io_acc_b_data_bits_0_22),
    .io_acc_b_data_bits_0_23(alu_io_acc_b_data_bits_0_23),
    .io_acc_b_data_bits_0_24(alu_io_acc_b_data_bits_0_24),
    .io_acc_b_data_bits_0_25(alu_io_acc_b_data_bits_0_25),
    .io_acc_b_data_bits_0_26(alu_io_acc_b_data_bits_0_26),
    .io_acc_b_data_bits_0_27(alu_io_acc_b_data_bits_0_27),
    .io_acc_b_data_bits_0_28(alu_io_acc_b_data_bits_0_28),
    .io_acc_b_data_bits_0_29(alu_io_acc_b_data_bits_0_29),
    .io_acc_b_data_bits_0_30(alu_io_acc_b_data_bits_0_30),
    .io_acc_b_data_bits_0_31(alu_io_acc_b_data_bits_0_31),
    .io_acc_y_data_valid(alu_io_acc_y_data_valid),
    .io_acc_y_data_bits_0_0(alu_io_acc_y_data_bits_0_0),
    .io_acc_y_data_bits_0_1(alu_io_acc_y_data_bits_0_1),
    .io_acc_y_data_bits_0_2(alu_io_acc_y_data_bits_0_2),
    .io_acc_y_data_bits_0_3(alu_io_acc_y_data_bits_0_3),
    .io_acc_y_data_bits_0_4(alu_io_acc_y_data_bits_0_4),
    .io_acc_y_data_bits_0_5(alu_io_acc_y_data_bits_0_5),
    .io_acc_y_data_bits_0_6(alu_io_acc_y_data_bits_0_6),
    .io_acc_y_data_bits_0_7(alu_io_acc_y_data_bits_0_7),
    .io_acc_y_data_bits_0_8(alu_io_acc_y_data_bits_0_8),
    .io_acc_y_data_bits_0_9(alu_io_acc_y_data_bits_0_9),
    .io_acc_y_data_bits_0_10(alu_io_acc_y_data_bits_0_10),
    .io_acc_y_data_bits_0_11(alu_io_acc_y_data_bits_0_11),
    .io_acc_y_data_bits_0_12(alu_io_acc_y_data_bits_0_12),
    .io_acc_y_data_bits_0_13(alu_io_acc_y_data_bits_0_13),
    .io_acc_y_data_bits_0_14(alu_io_acc_y_data_bits_0_14),
    .io_acc_y_data_bits_0_15(alu_io_acc_y_data_bits_0_15),
    .io_acc_y_data_bits_0_16(alu_io_acc_y_data_bits_0_16),
    .io_acc_y_data_bits_0_17(alu_io_acc_y_data_bits_0_17),
    .io_acc_y_data_bits_0_18(alu_io_acc_y_data_bits_0_18),
    .io_acc_y_data_bits_0_19(alu_io_acc_y_data_bits_0_19),
    .io_acc_y_data_bits_0_20(alu_io_acc_y_data_bits_0_20),
    .io_acc_y_data_bits_0_21(alu_io_acc_y_data_bits_0_21),
    .io_acc_y_data_bits_0_22(alu_io_acc_y_data_bits_0_22),
    .io_acc_y_data_bits_0_23(alu_io_acc_y_data_bits_0_23),
    .io_acc_y_data_bits_0_24(alu_io_acc_y_data_bits_0_24),
    .io_acc_y_data_bits_0_25(alu_io_acc_y_data_bits_0_25),
    .io_acc_y_data_bits_0_26(alu_io_acc_y_data_bits_0_26),
    .io_acc_y_data_bits_0_27(alu_io_acc_y_data_bits_0_27),
    .io_acc_y_data_bits_0_28(alu_io_acc_y_data_bits_0_28),
    .io_acc_y_data_bits_0_29(alu_io_acc_y_data_bits_0_29),
    .io_acc_y_data_bits_0_30(alu_io_acc_y_data_bits_0_30),
    .io_acc_y_data_bits_0_31(alu_io_acc_y_data_bits_0_31),
    .io_out_data_valid(alu_io_out_data_valid),
    .io_out_data_bits_0_0(alu_io_out_data_bits_0_0),
    .io_out_data_bits_0_1(alu_io_out_data_bits_0_1),
    .io_out_data_bits_0_2(alu_io_out_data_bits_0_2),
    .io_out_data_bits_0_3(alu_io_out_data_bits_0_3),
    .io_out_data_bits_0_4(alu_io_out_data_bits_0_4),
    .io_out_data_bits_0_5(alu_io_out_data_bits_0_5),
    .io_out_data_bits_0_6(alu_io_out_data_bits_0_6),
    .io_out_data_bits_0_7(alu_io_out_data_bits_0_7),
    .io_out_data_bits_0_8(alu_io_out_data_bits_0_8),
    .io_out_data_bits_0_9(alu_io_out_data_bits_0_9),
    .io_out_data_bits_0_10(alu_io_out_data_bits_0_10),
    .io_out_data_bits_0_11(alu_io_out_data_bits_0_11),
    .io_out_data_bits_0_12(alu_io_out_data_bits_0_12),
    .io_out_data_bits_0_13(alu_io_out_data_bits_0_13),
    .io_out_data_bits_0_14(alu_io_out_data_bits_0_14),
    .io_out_data_bits_0_15(alu_io_out_data_bits_0_15),
    .io_out_data_bits_0_16(alu_io_out_data_bits_0_16),
    .io_out_data_bits_0_17(alu_io_out_data_bits_0_17),
    .io_out_data_bits_0_18(alu_io_out_data_bits_0_18),
    .io_out_data_bits_0_19(alu_io_out_data_bits_0_19),
    .io_out_data_bits_0_20(alu_io_out_data_bits_0_20),
    .io_out_data_bits_0_21(alu_io_out_data_bits_0_21),
    .io_out_data_bits_0_22(alu_io_out_data_bits_0_22),
    .io_out_data_bits_0_23(alu_io_out_data_bits_0_23),
    .io_out_data_bits_0_24(alu_io_out_data_bits_0_24),
    .io_out_data_bits_0_25(alu_io_out_data_bits_0_25),
    .io_out_data_bits_0_26(alu_io_out_data_bits_0_26),
    .io_out_data_bits_0_27(alu_io_out_data_bits_0_27),
    .io_out_data_bits_0_28(alu_io_out_data_bits_0_28),
    .io_out_data_bits_0_29(alu_io_out_data_bits_0_29),
    .io_out_data_bits_0_30(alu_io_out_data_bits_0_30),
    .io_out_data_bits_0_31(alu_io_out_data_bits_0_31)
  );
  assign io_done = state == 2'h0 & io_start ? 1'h0 : _GEN_3; // @[TensorAlu.scala 209:11 210:37]
  assign io_uop_idx_valid = index_generator_io_valid | index_generator_io_src_valid; // @[TensorAlu.scala 223:48]
  assign io_uop_idx_bits = index_generator_io_uop_idx; // @[TensorAlu.scala 224:19]
  assign io_acc_rd_0_idx_valid = io_acc_rd_0_idx_valid_REG; // @[TensorAlu.scala 268:30]
  assign io_acc_rd_0_idx_bits = io_acc_rd_0_idx_bits_REG[6:0]; // @[TensorAlu.scala 283:29]
  assign io_acc_wr_0_valid = valid_r4; // @[TensorAlu.scala 360:26]
  assign io_acc_wr_0_bits_idx = dst_idx_r4[6:0]; // @[TensorAlu.scala 361:29]
  assign io_acc_wr_0_bits_data_0_0 = alu_io_acc_y_data_bits_0_0; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_1 = alu_io_acc_y_data_bits_0_1; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_2 = alu_io_acc_y_data_bits_0_2; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_3 = alu_io_acc_y_data_bits_0_3; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_4 = alu_io_acc_y_data_bits_0_4; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_5 = alu_io_acc_y_data_bits_0_5; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_6 = alu_io_acc_y_data_bits_0_6; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_7 = alu_io_acc_y_data_bits_0_7; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_8 = alu_io_acc_y_data_bits_0_8; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_9 = alu_io_acc_y_data_bits_0_9; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_10 = alu_io_acc_y_data_bits_0_10; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_11 = alu_io_acc_y_data_bits_0_11; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_12 = alu_io_acc_y_data_bits_0_12; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_13 = alu_io_acc_y_data_bits_0_13; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_14 = alu_io_acc_y_data_bits_0_14; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_15 = alu_io_acc_y_data_bits_0_15; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_16 = alu_io_acc_y_data_bits_0_16; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_17 = alu_io_acc_y_data_bits_0_17; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_18 = alu_io_acc_y_data_bits_0_18; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_19 = alu_io_acc_y_data_bits_0_19; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_20 = alu_io_acc_y_data_bits_0_20; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_21 = alu_io_acc_y_data_bits_0_21; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_22 = alu_io_acc_y_data_bits_0_22; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_23 = alu_io_acc_y_data_bits_0_23; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_24 = alu_io_acc_y_data_bits_0_24; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_25 = alu_io_acc_y_data_bits_0_25; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_26 = alu_io_acc_y_data_bits_0_26; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_27 = alu_io_acc_y_data_bits_0_27; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_28 = alu_io_acc_y_data_bits_0_28; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_29 = alu_io_acc_y_data_bits_0_29; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_30 = alu_io_acc_y_data_bits_0_30; // @[TensorAlu.scala 367:62]
  assign io_acc_wr_0_bits_data_0_31 = alu_io_acc_y_data_bits_0_31; // @[TensorAlu.scala 367:62]
  assign io_out_wr_0_valid = valid_r4; // @[TensorAlu.scala 381:22]
  assign io_out_wr_0_bits_idx = dst_idx_r4[6:0]; // @[TensorAlu.scala 382:25]
  assign io_out_wr_0_bits_data_0_0 = alu_io_out_data_bits_0_0; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_1 = alu_io_out_data_bits_0_1; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_2 = alu_io_out_data_bits_0_2; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_3 = alu_io_out_data_bits_0_3; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_4 = alu_io_out_data_bits_0_4; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_5 = alu_io_out_data_bits_0_5; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_6 = alu_io_out_data_bits_0_6; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_7 = alu_io_out_data_bits_0_7; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_8 = alu_io_out_data_bits_0_8; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_9 = alu_io_out_data_bits_0_9; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_10 = alu_io_out_data_bits_0_10; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_11 = alu_io_out_data_bits_0_11; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_12 = alu_io_out_data_bits_0_12; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_13 = alu_io_out_data_bits_0_13; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_14 = alu_io_out_data_bits_0_14; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_15 = alu_io_out_data_bits_0_15; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_16 = alu_io_out_data_bits_0_16; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_17 = alu_io_out_data_bits_0_17; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_18 = alu_io_out_data_bits_0_18; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_19 = alu_io_out_data_bits_0_19; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_20 = alu_io_out_data_bits_0_20; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_21 = alu_io_out_data_bits_0_21; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_22 = alu_io_out_data_bits_0_22; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_23 = alu_io_out_data_bits_0_23; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_24 = alu_io_out_data_bits_0_24; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_25 = alu_io_out_data_bits_0_25; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_26 = alu_io_out_data_bits_0_26; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_27 = alu_io_out_data_bits_0_27; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_28 = alu_io_out_data_bits_0_28; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_29 = alu_io_out_data_bits_0_29; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_30 = alu_io_out_data_bits_0_30; // @[TensorAlu.scala 289:21 375:66]
  assign io_out_wr_0_bits_data_0_31 = alu_io_out_data_bits_0_31; // @[TensorAlu.scala 289:21 375:66]
  assign index_generator_clock = clock;
  assign index_generator_reset = reset;
  assign index_generator_io_start = io_start; // @[TensorAlu.scala 219:28]
  assign index_generator_io_dec_alu_use_imm = io_dec_alu_use_imm; // @[TensorAlu.scala 220:26]
  assign index_generator_io_dec_src_1 = io_dec_src_1; // @[TensorAlu.scala 220:26]
  assign index_generator_io_dec_src_0 = io_dec_src_0; // @[TensorAlu.scala 220:26]
  assign index_generator_io_dec_dst_1 = io_dec_dst_1; // @[TensorAlu.scala 220:26]
  assign index_generator_io_dec_dst_0 = io_dec_dst_0; // @[TensorAlu.scala 220:26]
  assign index_generator_io_dec_lp_1 = io_dec_lp_1; // @[TensorAlu.scala 220:26]
  assign index_generator_io_dec_lp_0 = io_dec_lp_0; // @[TensorAlu.scala 220:26]
  assign index_generator_io_dec_uop_end = io_dec_uop_end; // @[TensorAlu.scala 220:26]
  assign index_generator_io_dec_uop_begin = io_dec_uop_begin; // @[TensorAlu.scala 220:26]
  assign alu_clock = clock;
  assign alu_io_opcode = neg_shift ? 3'h4 : io_dec_alu_op; // @[TensorAlu.scala 330:27]
  assign alu_io_acc_a_data_valid = alu_io_acc_a_data_valid_REG; // @[TensorAlu.scala 338:29]
  assign alu_io_acc_a_data_bits_0_0 = io_acc_rd_0_data_bits_0_0; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_1 = io_acc_rd_0_data_bits_0_1; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_2 = io_acc_rd_0_data_bits_0_2; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_3 = io_acc_rd_0_data_bits_0_3; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_4 = io_acc_rd_0_data_bits_0_4; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_5 = io_acc_rd_0_data_bits_0_5; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_6 = io_acc_rd_0_data_bits_0_6; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_7 = io_acc_rd_0_data_bits_0_7; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_8 = io_acc_rd_0_data_bits_0_8; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_9 = io_acc_rd_0_data_bits_0_9; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_10 = io_acc_rd_0_data_bits_0_10; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_11 = io_acc_rd_0_data_bits_0_11; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_12 = io_acc_rd_0_data_bits_0_12; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_13 = io_acc_rd_0_data_bits_0_13; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_14 = io_acc_rd_0_data_bits_0_14; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_15 = io_acc_rd_0_data_bits_0_15; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_16 = io_acc_rd_0_data_bits_0_16; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_17 = io_acc_rd_0_data_bits_0_17; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_18 = io_acc_rd_0_data_bits_0_18; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_19 = io_acc_rd_0_data_bits_0_19; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_20 = io_acc_rd_0_data_bits_0_20; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_21 = io_acc_rd_0_data_bits_0_21; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_22 = io_acc_rd_0_data_bits_0_22; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_23 = io_acc_rd_0_data_bits_0_23; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_24 = io_acc_rd_0_data_bits_0_24; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_25 = io_acc_rd_0_data_bits_0_25; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_26 = io_acc_rd_0_data_bits_0_26; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_27 = io_acc_rd_0_data_bits_0_27; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_28 = io_acc_rd_0_data_bits_0_28; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_29 = io_acc_rd_0_data_bits_0_29; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_30 = io_acc_rd_0_data_bits_0_30; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_a_data_bits_0_31 = io_acc_rd_0_data_bits_0_31; // @[TensorAlu.scala 291:24 344:47]
  assign alu_io_acc_b_data_valid = valid_r3; // @[TensorAlu.scala 352:35]
  assign alu_io_acc_b_data_bits_0_0 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_0; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_1 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_1; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_2 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_2; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_3 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_3; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_4 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_4; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_5 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_5; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_6 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_6; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_7 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_7; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_8 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_8; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_9 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_9; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_10 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_10; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_11 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_11; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_12 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_12; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_13 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_13; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_14 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_14; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_15 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_15; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_16 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_16; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_17 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_17; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_18 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_18; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_19 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_19; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_20 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_20; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_21 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_21; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_22 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_22; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_23 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_23; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_24 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_24; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_25 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_25; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_26 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_26; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_27 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_27; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_28 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_28; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_29 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_29; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_30 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_30; // @[TensorAlu.scala 355:34]
  assign alu_io_acc_b_data_bits_0_31 = io_dec_alu_use_imm ? tensorImm_data_bits_0_0 : save_src_0_31; // @[TensorAlu.scala 355:34]
  always @(posedge clock) begin
    if (reset) begin // @[TensorAlu.scala 202:22]
      state <= 2'h0; // @[TensorAlu.scala 202:22]
    end else if (state == 2'h0 & io_start) begin // @[TensorAlu.scala 210:37]
      state <= 2'h1; // @[TensorAlu.scala 211:11]
    end else if (state == 2'h1 & index_generator_io_last) begin // @[TensorAlu.scala 212:57]
      state <= 2'h2; // @[TensorAlu.scala 213:11]
    end else if (state == 2'h2 & inflight == 4'h0) begin // @[TensorAlu.scala 214:51]
      state <= 2'h0; // @[TensorAlu.scala 215:11]
    end
    if (reset) begin // @[TensorAlu.scala 203:25]
      inflight <= 4'h0; // @[TensorAlu.scala 203:25]
    end else if (_T) begin // @[TensorAlu.scala 239:25]
      inflight <= 4'h0; // @[TensorAlu.scala 241:14]
    end else if (!(index_generator_io_valid & valid_r4)) begin // @[TensorAlu.scala 231:46]
      if (index_generator_io_valid) begin // @[TensorAlu.scala 232:40]
        inflight <= _inflight_T_1; // @[TensorAlu.scala 234:14]
      end else begin
        inflight <= _GEN_7;
      end
    end
    if (reset) begin // @[Reg.scala 28:20]
      valid_r1 <= 1'h0; // @[Reg.scala 28:20]
    end else begin
      valid_r1 <= _GEN_6;
    end
    if (reset) begin // @[TensorAlu.scala 227:25]
      valid_r2 <= 1'h0; // @[TensorAlu.scala 227:25]
    end else begin
      valid_r2 <= valid_r1; // @[TensorAlu.scala 227:25]
    end
    if (reset) begin // @[TensorAlu.scala 228:25]
      valid_r3 <= 1'h0; // @[TensorAlu.scala 228:25]
    end else begin
      valid_r3 <= valid_r2; // @[TensorAlu.scala 228:25]
    end
    if (reset) begin // @[TensorAlu.scala 229:25]
      valid_r4 <= 1'h0; // @[TensorAlu.scala 229:25]
    end else begin
      valid_r4 <= valid_r3; // @[TensorAlu.scala 229:25]
    end
    if (reset) begin // @[Reg.scala 28:20]
      src_valid_r1 <= 1'h0; // @[Reg.scala 28:20]
    end else begin
      src_valid_r1 <= _GEN_11;
    end
    if (reset) begin // @[TensorAlu.scala 248:29]
      src_valid_r2 <= 1'h0; // @[TensorAlu.scala 248:29]
    end else begin
      src_valid_r2 <= src_valid_r1; // @[TensorAlu.scala 248:29]
    end
    if (reset) begin // @[TensorAlu.scala 249:29]
      src_valid_r3 <= 1'h0; // @[TensorAlu.scala 249:29]
    end else begin
      src_valid_r3 <= src_valid_r2; // @[TensorAlu.scala 249:29]
    end
    dst_idx_r1 <= index_generator_io_dst_idx; // @[Reg.scala 16:16 17:{18,22}]
    src_idx_r1 <= index_generator_io_src_idx; // @[Reg.scala 16:16 17:{18,22}]
    io_acc_rd_0_idx_valid_REG <= valid_r1 | src_valid_r1; // @[TensorAlu.scala 266:32]
    src_idx_r2 <= _GEN_15 + src_offset; // @[TensorAlu.scala 271:35]
    src_idx_r3 <= src_idx_r2; // @[TensorAlu.scala 273:27]
    dst_idx_r2 <= _GEN_16 + io_uop_data_bits_u0; // @[TensorAlu.scala 275:35]
    dst_idx_r3 <= dst_idx_r2; // @[TensorAlu.scala 277:27]
    dst_idx_r4 <= dst_idx_r3; // @[TensorAlu.scala 278:27]
    if (src_valid_r1 | io_dec_alu_use_imm) begin // @[TensorAlu.scala 281:25]
      io_acc_rd_0_idx_bits_REG <= new_src_idx_r1;
    end else begin
      io_acc_rd_0_idx_bits_REG <= {{7'd0}, new_dst_idx_r1};
    end
    save_src_0_0 <= io_acc_rd_0_data_bits_0_0; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_1 <= io_acc_rd_0_data_bits_0_1; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_2 <= io_acc_rd_0_data_bits_0_2; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_3 <= io_acc_rd_0_data_bits_0_3; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_4 <= io_acc_rd_0_data_bits_0_4; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_5 <= io_acc_rd_0_data_bits_0_5; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_6 <= io_acc_rd_0_data_bits_0_6; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_7 <= io_acc_rd_0_data_bits_0_7; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_8 <= io_acc_rd_0_data_bits_0_8; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_9 <= io_acc_rd_0_data_bits_0_9; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_10 <= io_acc_rd_0_data_bits_0_10; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_11 <= io_acc_rd_0_data_bits_0_11; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_12 <= io_acc_rd_0_data_bits_0_12; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_13 <= io_acc_rd_0_data_bits_0_13; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_14 <= io_acc_rd_0_data_bits_0_14; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_15 <= io_acc_rd_0_data_bits_0_15; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_16 <= io_acc_rd_0_data_bits_0_16; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_17 <= io_acc_rd_0_data_bits_0_17; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_18 <= io_acc_rd_0_data_bits_0_18; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_19 <= io_acc_rd_0_data_bits_0_19; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_20 <= io_acc_rd_0_data_bits_0_20; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_21 <= io_acc_rd_0_data_bits_0_21; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_22 <= io_acc_rd_0_data_bits_0_22; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_23 <= io_acc_rd_0_data_bits_0_23; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_24 <= io_acc_rd_0_data_bits_0_24; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_25 <= io_acc_rd_0_data_bits_0_25; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_26 <= io_acc_rd_0_data_bits_0_26; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_27 <= io_acc_rd_0_data_bits_0_27; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_28 <= io_acc_rd_0_data_bits_0_28; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_29 <= io_acc_rd_0_data_bits_0_29; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_30 <= io_acc_rd_0_data_bits_0_30; // @[TensorAlu.scala 290:24 307:47]
    save_src_0_31 <= io_acc_rd_0_data_bits_0_31; // @[TensorAlu.scala 290:24 307:47]
    alu_io_acc_a_data_valid_REG <= valid_r2; // @[TensorAlu.scala 338:39]
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_7 & index_generator_io_valid & ~reset & ~(inflight != 4'hf)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorAlu.scala:233 assert(inflight =/= ((1<<inflightBits)-1).U)\n"); // @[TensorAlu.scala 233:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_18 & ~index_generator_io_valid & valid_r4 & _T_10 & ~(inflight != 4'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TensorAlu.scala:236 assert(inflight =/= 0.U)\n"); // @[TensorAlu.scala 236:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & _T_10 & ~_T_5) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TensorAlu.scala:240 assert(inflight === 0.U)\n"); // @[TensorAlu.scala 240:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(io_acc_rd_0_data_valid == (valid_r3 | src_valid_r3))) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorAlu.scala:284 assert(io.acc.rd(idx).data.valid === (valid_r3 || src_valid_r3))\n"
            ); // @[TensorAlu.scala 284:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~valid_r3 | io_acc_rd_0_data_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorAlu.scala:336 assert(!valid_r3 || io.acc.rd(idx).data.valid)\n"); // @[TensorAlu.scala 336:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(alu_io_acc_y_data_valid == valid_r4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorAlu.scala:359 assert(alu.io.acc_y.data.valid === valid_r4)\n"); // @[TensorAlu.scala 359:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(alu_io_out_data_valid == valid_r4)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorAlu.scala:372 assert(alu.io.out.data.valid === valid_r4)\n"); // @[TensorAlu.scala 372:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~bypass_dst)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Bypass required on dst_idx read TensorAlu.dst_idx_r3: Reg[UInt] RAW with write TensorAlu.dst_idx_r4: Reg[UInt]\n\n    at TensorAlu.scala:390 assert(!bypass_dst, s\"Bypass required on dst_idx read $dst_idx_r3 RAW with write $dst_idx_r4\\n\")\n"
            ); // @[TensorAlu.scala 390:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & ~(~bypass_src)) begin
          $fwrite(32'h80000002,
            "Assertion failed: Bypass required on src_idx read TensorAlu.src_idx_r3: Reg[UInt] RAW with write TensorAlu.dst_idx_r4: Reg[UInt]\n\n    at TensorAlu.scala:391 assert(!bypass_src, s\"Bypass required on src_idx read $src_idx_r3 RAW with write $dst_idx_r4\\n\")\n"
            ); // @[TensorAlu.scala 391:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflight = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  valid_r1 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  valid_r2 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  valid_r3 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  valid_r4 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  src_valid_r1 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  src_valid_r2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  src_valid_r3 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  dst_idx_r1 = _RAND_9[6:0];
  _RAND_10 = {1{`RANDOM}};
  src_idx_r1 = _RAND_10[6:0];
  _RAND_11 = {1{`RANDOM}};
  io_acc_rd_0_idx_valid_REG = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  src_idx_r2 = _RAND_12[17:0];
  _RAND_13 = {1{`RANDOM}};
  src_idx_r3 = _RAND_13[17:0];
  _RAND_14 = {1{`RANDOM}};
  dst_idx_r2 = _RAND_14[10:0];
  _RAND_15 = {1{`RANDOM}};
  dst_idx_r3 = _RAND_15[10:0];
  _RAND_16 = {1{`RANDOM}};
  dst_idx_r4 = _RAND_16[10:0];
  _RAND_17 = {1{`RANDOM}};
  io_acc_rd_0_idx_bits_REG = _RAND_17[17:0];
  _RAND_18 = {1{`RANDOM}};
  save_src_0_0 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  save_src_0_1 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  save_src_0_2 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  save_src_0_3 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  save_src_0_4 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  save_src_0_5 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  save_src_0_6 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  save_src_0_7 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  save_src_0_8 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  save_src_0_9 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  save_src_0_10 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  save_src_0_11 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  save_src_0_12 = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  save_src_0_13 = _RAND_31[31:0];
  _RAND_32 = {1{`RANDOM}};
  save_src_0_14 = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  save_src_0_15 = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  save_src_0_16 = _RAND_34[31:0];
  _RAND_35 = {1{`RANDOM}};
  save_src_0_17 = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  save_src_0_18 = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  save_src_0_19 = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  save_src_0_20 = _RAND_38[31:0];
  _RAND_39 = {1{`RANDOM}};
  save_src_0_21 = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  save_src_0_22 = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  save_src_0_23 = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  save_src_0_24 = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  save_src_0_25 = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  save_src_0_26 = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  save_src_0_27 = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  save_src_0_28 = _RAND_46[31:0];
  _RAND_47 = {1{`RANDOM}};
  save_src_0_29 = _RAND_47[31:0];
  _RAND_48 = {1{`RANDOM}};
  save_src_0_30 = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  save_src_0_31 = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  alu_io_acc_a_data_valid_REG = _RAND_50[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~_T_7 & index_generator_io_valid & ~reset) begin
      assert(inflight != 4'hf); // @[TensorAlu.scala 233:11]
    end
    //
    if (_GEN_18 & ~index_generator_io_valid & valid_r4 & _T_10) begin
      assert(inflight != 4'h0); // @[TensorAlu.scala 236:11]
    end
    //
    if (_T & _T_10) begin
      assert(_T_5); // @[TensorAlu.scala 240:11]
    end
    //
    if (_T_10) begin
      assert(io_acc_rd_0_data_valid == (valid_r3 | src_valid_r3)); // @[TensorAlu.scala 284:11]
    end
    //
    if (_T_10) begin
      assert(~valid_r3 | io_acc_rd_0_data_valid); // @[TensorAlu.scala 336:11]
    end
    //
    if (_T_10) begin
      assert(alu_io_acc_y_data_valid == valid_r4); // @[TensorAlu.scala 359:11]
    end
    //
    if (_T_10) begin
      assert(alu_io_out_data_valid == valid_r4); // @[TensorAlu.scala 372:11]
    end
    //
    if (_T_10) begin
      assert(~bypass_dst); // @[TensorAlu.scala 390:9]
    end
    //
    if (_T_10) begin
      assert(~bypass_src); // @[TensorAlu.scala 391:9]
    end
  end
endmodule
module TwoPortMem_1(
  input          clock,
  input          io_wr_en,
  input  [15:0]  io_wr_addr,
  input  [127:0] io_wr_data,
  input          io_rd_en,
  input  [15:0]  io_rd_addr,
  output [127:0] io_rd_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [127:0] mem [0:31]; // @[SyncQueue.scala 496:24]
  wire  mem_io_rd_data_MPORT_en; // @[SyncQueue.scala 496:24]
  wire [4:0] mem_io_rd_data_MPORT_addr; // @[SyncQueue.scala 496:24]
  wire [127:0] mem_io_rd_data_MPORT_data; // @[SyncQueue.scala 496:24]
  wire [127:0] mem_MPORT_data; // @[SyncQueue.scala 496:24]
  wire [4:0] mem_MPORT_addr; // @[SyncQueue.scala 496:24]
  wire  mem_MPORT_mask; // @[SyncQueue.scala 496:24]
  wire  mem_MPORT_en; // @[SyncQueue.scala 496:24]
  reg  mem_io_rd_data_MPORT_en_pipe_0;
  reg [4:0] mem_io_rd_data_MPORT_addr_pipe_0;
  assign mem_io_rd_data_MPORT_en = mem_io_rd_data_MPORT_en_pipe_0;
  assign mem_io_rd_data_MPORT_addr = mem_io_rd_data_MPORT_addr_pipe_0;
  assign mem_io_rd_data_MPORT_data = mem[mem_io_rd_data_MPORT_addr]; // @[SyncQueue.scala 496:24]
  assign mem_MPORT_data = io_wr_data;
  assign mem_MPORT_addr = io_wr_addr[4:0];
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_wr_en;
  assign io_rd_data = mem_io_rd_data_MPORT_data; // @[SyncQueue.scala 502:20 503:16]
  always @(posedge clock) begin
    if (mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[SyncQueue.scala 496:24]
    end
    mem_io_rd_data_MPORT_en_pipe_0 <= io_rd_en;
    if (io_rd_en) begin
      mem_io_rd_data_MPORT_addr_pipe_0 <= io_rd_addr[4:0];
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    mem[initvar] = _RAND_0[127:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_io_rd_data_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  mem_io_rd_data_MPORT_addr_pipe_0 = _RAND_2[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module OneCycleQueue_1(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [127:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [127:0] io_deq_bits,
  output [5:0]   io_count
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  ram0_clock; // @[SyncQueue.scala 377:20]
  wire  ram0_io_wr_en; // @[SyncQueue.scala 377:20]
  wire [15:0] ram0_io_wr_addr; // @[SyncQueue.scala 377:20]
  wire [127:0] ram0_io_wr_data; // @[SyncQueue.scala 377:20]
  wire  ram0_io_rd_en; // @[SyncQueue.scala 377:20]
  wire [15:0] ram0_io_rd_addr; // @[SyncQueue.scala 377:20]
  wire [127:0] ram0_io_rd_data; // @[SyncQueue.scala 377:20]
  reg [4:0] value; // @[Counter.scala 62:40]
  reg [4:0] value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[SyncQueue.scala 380:27]
  wire  ptr_match = value == value_1; // @[SyncQueue.scala 383:33]
  wire  empty = ptr_match & ~maybe_full; // @[SyncQueue.scala 384:25]
  wire  full = ptr_match & maybe_full; // @[SyncQueue.scala 385:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  wrap = value_1 == 5'h1f; // @[Counter.scala 74:24]
  wire [4:0] _value_T_1 = value_1 + 5'h1; // @[Counter.scala 78:24]
  wire [4:0] _value_T_3 = value + 5'h1; // @[Counter.scala 78:24]
  wire  _firstRead_T_1 = do_enq & io_count == 6'h0; // @[SyncQueue.scala 403:43]
  reg  firstRead; // @[Reg.scala 28:20]
  wire  _io_deq_valid_T_1 = ~firstRead; // @[SyncQueue.scala 404:29]
  wire [4:0] _GEN_4 = wrap ? 5'h0 : _value_T_1; // @[SyncQueue.scala 413:17 414:14 416:14]
  wire [4:0] _GEN_5 = do_deq ? _GEN_4 : value_1; // @[SyncQueue.scala 411:23 419:12]
  wire [4:0] rdAddr = firstRead ? value_1 : _GEN_5; // @[SyncQueue.scala 409:19 410:12]
  wire [4:0] ptr_diff = value - value_1; // @[SyncQueue.scala 430:32]
  wire [5:0] _io_count_T_1 = maybe_full & ptr_match ? 6'h20 : 6'h0; // @[SyncQueue.scala 432:20]
  wire [5:0] _GEN_7 = {{1'd0}, ptr_diff}; // @[SyncQueue.scala 432:62]
  TwoPortMem_1 ram0 ( // @[SyncQueue.scala 377:20]
    .clock(ram0_clock),
    .io_wr_en(ram0_io_wr_en),
    .io_wr_addr(ram0_io_wr_addr),
    .io_wr_data(ram0_io_wr_data),
    .io_rd_en(ram0_io_rd_en),
    .io_rd_addr(ram0_io_rd_addr),
    .io_rd_data(ram0_io_rd_data)
  );
  assign io_enq_ready = ~full; // @[SyncQueue.scala 405:19]
  assign io_deq_valid = ~empty & ~firstRead; // @[SyncQueue.scala 404:26]
  assign io_deq_bits = ram0_io_rd_data; // @[SyncQueue.scala 426:15]
  assign io_count = _io_count_T_1 | _GEN_7; // @[SyncQueue.scala 432:62]
  assign ram0_clock = clock;
  assign ram0_io_wr_en = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  assign ram0_io_wr_addr = {{11'd0}, value}; // @[SyncQueue.scala 423:19]
  assign ram0_io_wr_data = io_enq_bits; // @[SyncQueue.scala 422:19]
  assign ram0_io_rd_en = do_deq | firstRead; // @[SyncQueue.scala 424:27]
  assign ram0_io_rd_addr = {{11'd0}, rdAddr}; // @[SyncQueue.scala 425:19]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 62:40]
      value <= 5'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[SyncQueue.scala 399:17]
      value <= _value_T_3; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[SyncQueue.scala 391:16]
      value_1 <= _value_T_1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[SyncQueue.scala 380:27]
      maybe_full <= 1'h0; // @[SyncQueue.scala 380:27]
    end else if (do_enq != do_deq) begin // @[SyncQueue.scala 395:27]
      maybe_full <= do_enq; // @[SyncQueue.scala 396:16]
    end
    if (reset) begin // @[Reg.scala 28:20]
      firstRead <= 1'h0; // @[Reg.scala 28:20]
    end else begin
      firstRead <= _firstRead_T_1;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(_io_deq_valid_T_1 | ~do_deq)) begin
          $fwrite(32'h80000002,
            "Assertion failed: -F- Cannot have deq with first read as queue output is not valid yet\n    at SyncQueue.scala:406 assert(!firstRead || !do_deq, \"-F- Cannot have deq with first read as queue output is not valid yet\")\n"
            ); // @[SyncQueue.scala 406:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  value_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  maybe_full = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  firstRead = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(_io_deq_valid_T_1 | ~do_deq); // @[SyncQueue.scala 406:9]
    end
  end
endmodule
module SyncQueue2PortMemImpl_1(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [127:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [127:0] io_deq_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  memoryQueue_clock; // @[SyncQueue.scala 172:27]
  wire  memoryQueue_reset; // @[SyncQueue.scala 172:27]
  wire  memoryQueue_io_enq_ready; // @[SyncQueue.scala 172:27]
  wire  memoryQueue_io_enq_valid; // @[SyncQueue.scala 172:27]
  wire [127:0] memoryQueue_io_enq_bits; // @[SyncQueue.scala 172:27]
  wire  memoryQueue_io_deq_ready; // @[SyncQueue.scala 172:27]
  wire  memoryQueue_io_deq_valid; // @[SyncQueue.scala 172:27]
  wire [127:0] memoryQueue_io_deq_bits; // @[SyncQueue.scala 172:27]
  wire [5:0] memoryQueue_io_count; // @[SyncQueue.scala 172:27]
  wire  buffer_clock; // @[SyncQueue.scala 173:22]
  wire  buffer_reset; // @[SyncQueue.scala 173:22]
  wire  buffer_io_enq_ready; // @[SyncQueue.scala 173:22]
  wire  buffer_io_enq_valid; // @[SyncQueue.scala 173:22]
  wire [127:0] buffer_io_enq_bits; // @[SyncQueue.scala 173:22]
  wire  buffer_io_deq_ready; // @[SyncQueue.scala 173:22]
  wire  buffer_io_deq_valid; // @[SyncQueue.scala 173:22]
  wire [127:0] buffer_io_deq_bits; // @[SyncQueue.scala 173:22]
  wire  memoryQueueHasValues = memoryQueue_io_count != 6'h0; // @[SyncQueue.scala 175:51]
  wire  _memoryQueue_io_enq_valid_T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _countNext_T_1 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire  _countNext_T_2 = _memoryQueue_io_enq_valid_T | _countNext_T_1; // @[SyncQueue.scala 190:26]
  reg [5:0] countNext; // @[Reg.scala 28:20]
  wire  _T_3 = _memoryQueue_io_enq_valid_T & ~_countNext_T_1; // @[SyncQueue.scala 191:21]
  wire [5:0] _count_T_1 = countNext + 6'h1; // @[SyncQueue.scala 193:24]
  wire  _T_11 = ~_memoryQueue_io_enq_valid_T & _countNext_T_1; // @[SyncQueue.scala 194:28]
  wire [5:0] _count_T_3 = countNext - 6'h1; // @[SyncQueue.scala 196:24]
  wire  _T_6 = ~reset; // @[SyncQueue.scala 192:11]
  OneCycleQueue_1 memoryQueue ( // @[SyncQueue.scala 172:27]
    .clock(memoryQueue_clock),
    .reset(memoryQueue_reset),
    .io_enq_ready(memoryQueue_io_enq_ready),
    .io_enq_valid(memoryQueue_io_enq_valid),
    .io_enq_bits(memoryQueue_io_enq_bits),
    .io_deq_ready(memoryQueue_io_deq_ready),
    .io_deq_valid(memoryQueue_io_deq_valid),
    .io_deq_bits(memoryQueue_io_deq_bits),
    .io_count(memoryQueue_io_count)
  );
  Queue_5 buffer ( // @[SyncQueue.scala 173:22]
    .clock(buffer_clock),
    .reset(buffer_reset),
    .io_enq_ready(buffer_io_enq_ready),
    .io_enq_valid(buffer_io_enq_valid),
    .io_enq_bits(buffer_io_enq_bits),
    .io_deq_ready(buffer_io_deq_ready),
    .io_deq_valid(buffer_io_deq_valid),
    .io_deq_bits(buffer_io_deq_bits)
  );
  assign io_enq_ready = countNext != 6'h20; // @[SyncQueue.scala 202:30]
  assign io_deq_valid = countNext != 6'h0; // @[SyncQueue.scala 203:30]
  assign io_deq_bits = buffer_io_deq_bits; // @[SyncQueue.scala 181:10]
  assign memoryQueue_clock = clock;
  assign memoryQueue_reset = reset;
  assign memoryQueue_io_enq_valid = _memoryQueue_io_enq_valid_T & (~buffer_io_enq_ready | memoryQueueHasValues); // @[SyncQueue.scala 183:43]
  assign memoryQueue_io_enq_bits = io_enq_bits; // @[SyncQueue.scala 182:27]
  assign memoryQueue_io_deq_ready = buffer_io_enq_ready; // @[SyncQueue.scala 184:28]
  assign buffer_clock = clock;
  assign buffer_reset = reset;
  assign buffer_io_enq_valid = memoryQueueHasValues ? memoryQueue_io_deq_valid : io_enq_valid; // @[SyncQueue.scala 176:26]
  assign buffer_io_enq_bits = memoryQueueHasValues ? memoryQueue_io_deq_bits : io_enq_bits; // @[SyncQueue.scala 177:25]
  assign buffer_io_deq_ready = io_deq_ready; // @[SyncQueue.scala 181:10]
  always @(posedge clock) begin
    if (reset) begin // @[Reg.scala 28:20]
      countNext <= 6'h0; // @[Reg.scala 28:20]
    end else if (_countNext_T_2) begin // @[Reg.scala 29:18]
      if (_memoryQueue_io_enq_valid_T & ~_countNext_T_1) begin // @[SyncQueue.scala 191:38]
        countNext <= _count_T_1; // @[SyncQueue.scala 193:11]
      end else if (~_memoryQueue_io_enq_valid_T & _countNext_T_1) begin // @[SyncQueue.scala 194:44]
        countNext <= _count_T_3; // @[SyncQueue.scala 196:11]
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_3 & ~reset & ~(countNext < 6'h20)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at SyncQueue.scala:192 assert(countNext < entries.U)\n"); // @[SyncQueue.scala 192:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T_3 & _T_11 & _T_6 & ~(countNext > 6'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at SyncQueue.scala:195 assert(countNext > 0.U)\n"); // @[SyncQueue.scala 195:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6 & ~(io_deq_valid == buffer_io_deq_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at SyncQueue.scala:204 assert(io.deq.valid === buffer.io.deq.valid)\n"); // @[SyncQueue.scala 204:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6 & ~(io_enq_ready == buffer_io_enq_ready | memoryQueue_io_enq_ready)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at SyncQueue.scala:205 assert(io.enq.ready === buffer.io.enq.ready || memoryQueue.io.enq.ready)\n"
            ); // @[SyncQueue.scala 205:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  countNext = _RAND_0[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T_3 & ~reset) begin
      assert(countNext < 6'h20); // @[SyncQueue.scala 192:11]
    end
    //
    if (~_T_3 & _T_11 & _T_6) begin
      assert(countNext > 6'h0); // @[SyncQueue.scala 195:11]
    end
    //
    if (_T_6) begin
      assert(io_deq_valid == buffer_io_deq_valid); // @[SyncQueue.scala 204:9]
    end
    //
    if (_T_6) begin
      assert(io_enq_ready == buffer_io_enq_ready | memoryQueue_io_enq_ready); // @[SyncQueue.scala 205:9]
    end
  end
endmodule
module SyncQueue2PortMem_1(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [127:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [127:0] io_deq_bits
);
  wire  queue_clock; // @[SyncQueue.scala 151:23]
  wire  queue_reset; // @[SyncQueue.scala 151:23]
  wire  queue_io_enq_ready; // @[SyncQueue.scala 151:23]
  wire  queue_io_enq_valid; // @[SyncQueue.scala 151:23]
  wire [127:0] queue_io_enq_bits; // @[SyncQueue.scala 151:23]
  wire  queue_io_deq_ready; // @[SyncQueue.scala 151:23]
  wire  queue_io_deq_valid; // @[SyncQueue.scala 151:23]
  wire [127:0] queue_io_deq_bits; // @[SyncQueue.scala 151:23]
  SyncQueue2PortMemImpl_1 queue ( // @[SyncQueue.scala 151:23]
    .clock(queue_clock),
    .reset(queue_reset),
    .io_enq_ready(queue_io_enq_ready),
    .io_enq_valid(queue_io_enq_valid),
    .io_enq_bits(queue_io_enq_bits),
    .io_deq_ready(queue_io_deq_ready),
    .io_deq_valid(queue_io_deq_valid),
    .io_deq_bits(queue_io_deq_bits)
  );
  assign io_enq_ready = queue_io_enq_ready; // @[SyncQueue.scala 152:8]
  assign io_deq_valid = queue_io_deq_valid; // @[SyncQueue.scala 152:8]
  assign io_deq_bits = queue_io_deq_bits; // @[SyncQueue.scala 152:8]
  assign queue_clock = clock;
  assign queue_reset = reset;
  assign queue_io_enq_valid = io_enq_valid; // @[SyncQueue.scala 152:8]
  assign queue_io_enq_bits = io_enq_bits; // @[SyncQueue.scala 152:8]
  assign queue_io_deq_ready = io_deq_ready; // @[SyncQueue.scala 152:8]
endmodule
module SyncQueue_1(
  input          clock,
  input          reset,
  output         io_enq_ready,
  input          io_enq_valid,
  input  [127:0] io_enq_bits,
  input          io_deq_ready,
  output         io_deq_valid,
  output [127:0] io_deq_bits
);
  wire  queue_clock; // @[SyncQueue.scala 47:23]
  wire  queue_reset; // @[SyncQueue.scala 47:23]
  wire  queue_io_enq_ready; // @[SyncQueue.scala 47:23]
  wire  queue_io_enq_valid; // @[SyncQueue.scala 47:23]
  wire [127:0] queue_io_enq_bits; // @[SyncQueue.scala 47:23]
  wire  queue_io_deq_ready; // @[SyncQueue.scala 47:23]
  wire  queue_io_deq_valid; // @[SyncQueue.scala 47:23]
  wire [127:0] queue_io_deq_bits; // @[SyncQueue.scala 47:23]
  SyncQueue2PortMem_1 queue ( // @[SyncQueue.scala 47:23]
    .clock(queue_clock),
    .reset(queue_reset),
    .io_enq_ready(queue_io_enq_ready),
    .io_enq_valid(queue_io_enq_valid),
    .io_enq_bits(queue_io_enq_bits),
    .io_deq_ready(queue_io_deq_ready),
    .io_deq_valid(queue_io_deq_valid),
    .io_deq_bits(queue_io_deq_bits)
  );
  assign io_enq_ready = queue_io_enq_ready; // @[SyncQueue.scala 48:8]
  assign io_deq_valid = queue_io_deq_valid; // @[SyncQueue.scala 48:8]
  assign io_deq_bits = queue_io_deq_bits; // @[SyncQueue.scala 48:8]
  assign queue_clock = clock;
  assign queue_reset = reset;
  assign queue_io_enq_valid = io_enq_valid; // @[SyncQueue.scala 48:8]
  assign queue_io_enq_bits = io_enq_bits; // @[SyncQueue.scala 48:8]
  assign queue_io_deq_ready = io_deq_ready; // @[SyncQueue.scala 48:8]
endmodule
module ComputeDecode(
  input  [127:0] io_inst,
  output         io_push_next,
  output         io_push_prev,
  output         io_pop_next,
  output         io_pop_prev,
  output         io_isLoadAcc,
  output         io_isLoadUop,
  output         io_isSync,
  output         io_isAlu,
  output         io_isGemm,
  output         io_isFinish
);
  wire [15:0] dec_xsize = io_inst[95:80]; // @[Decode.scala 199:29]
  wire [127:0] _io_isLoadAcc_T = io_inst & 128'h387; // @[Decode.scala 204:27]
  wire  _io_isLoadAcc_T_1 = 128'h180 == _io_isLoadAcc_T; // @[Decode.scala 204:27]
  wire  _io_isLoadAcc_T_2 = dec_xsize != 16'h0; // @[Decode.scala 204:48]
  wire  _io_isLoadUop_T_1 = 128'h0 == _io_isLoadAcc_T; // @[Decode.scala 205:27]
  wire [127:0] _io_isAlu_T = io_inst & 128'h7000000000000000000000000007; // @[Decode.scala 207:23]
  wire [127:0] _io_isGemm_T = io_inst & 128'h7; // @[Decode.scala 208:24]
  assign io_push_next = io_inst[6]; // @[Decode.scala 199:29]
  assign io_push_prev = io_inst[5]; // @[Decode.scala 199:29]
  assign io_pop_next = io_inst[4]; // @[Decode.scala 199:29]
  assign io_pop_prev = io_inst[3]; // @[Decode.scala 199:29]
  assign io_isLoadAcc = 128'h180 == _io_isLoadAcc_T & dec_xsize != 16'h0; // @[Decode.scala 204:36]
  assign io_isLoadUop = 128'h0 == _io_isLoadAcc_T & _io_isLoadAcc_T_2; // @[Decode.scala 205:36]
  assign io_isSync = (_io_isLoadAcc_T_1 | _io_isLoadUop_T_1) & dec_xsize == 16'h0; // @[Decode.scala 206:54]
  assign io_isAlu = 128'h4 == _io_isAlu_T | 128'h1000000000000000000000000004 == _io_isAlu_T | 128'h2000000000000000000000000004
     == _io_isAlu_T | 128'h3000000000000000000000000004 == _io_isAlu_T; // @[Decode.scala 207:70]
  assign io_isGemm = 128'h2 == _io_isGemm_T; // @[Decode.scala 208:24]
  assign io_isFinish = 128'h3 == _io_isGemm_T; // @[Decode.scala 209:26]
endmodule
module Compute(
  input          clock,
  input          reset,
  input          io_i_post_0,
  input          io_i_post_1,
  output         io_o_post_0,
  output         io_o_post_1,
  output         io_inst_ready,
  input          io_inst_valid,
  input  [127:0] io_inst_bits,
  input  [31:0]  io_uop_baddr,
  input  [31:0]  io_acc_baddr,
  input          io_vme_rd_0_cmd_ready,
  output         io_vme_rd_0_cmd_valid,
  output [31:0]  io_vme_rd_0_cmd_bits_addr,
  output [3:0]   io_vme_rd_0_cmd_bits_len,
  output [20:0]  io_vme_rd_0_cmd_bits_tag,
  input          io_vme_rd_0_data_valid,
  input  [63:0]  io_vme_rd_0_data_bits_data,
  input  [20:0]  io_vme_rd_0_data_bits_tag,
  input          io_vme_rd_0_data_bits_last,
  input          io_vme_rd_1_cmd_ready,
  output         io_vme_rd_1_cmd_valid,
  output [31:0]  io_vme_rd_1_cmd_bits_addr,
  output [3:0]   io_vme_rd_1_cmd_bits_len,
  output [20:0]  io_vme_rd_1_cmd_bits_tag,
  input          io_vme_rd_1_data_valid,
  input  [63:0]  io_vme_rd_1_data_bits_data,
  input  [20:0]  io_vme_rd_1_data_bits_tag,
  output         io_inp_rd_0_idx_valid,
  output [6:0]   io_inp_rd_0_idx_bits,
  input          io_inp_rd_0_data_valid,
  input  [7:0]   io_inp_rd_0_data_bits_0_0,
  input  [7:0]   io_inp_rd_0_data_bits_0_1,
  input  [7:0]   io_inp_rd_0_data_bits_0_2,
  input  [7:0]   io_inp_rd_0_data_bits_0_3,
  input  [7:0]   io_inp_rd_0_data_bits_0_4,
  input  [7:0]   io_inp_rd_0_data_bits_0_5,
  input  [7:0]   io_inp_rd_0_data_bits_0_6,
  input  [7:0]   io_inp_rd_0_data_bits_0_7,
  input  [7:0]   io_inp_rd_0_data_bits_0_8,
  input  [7:0]   io_inp_rd_0_data_bits_0_9,
  input  [7:0]   io_inp_rd_0_data_bits_0_10,
  input  [7:0]   io_inp_rd_0_data_bits_0_11,
  input  [7:0]   io_inp_rd_0_data_bits_0_12,
  input  [7:0]   io_inp_rd_0_data_bits_0_13,
  input  [7:0]   io_inp_rd_0_data_bits_0_14,
  input  [7:0]   io_inp_rd_0_data_bits_0_15,
  output         io_wgt_rd_0_idx_valid,
  output [5:0]   io_wgt_rd_0_idx_bits,
  input          io_wgt_rd_0_data_valid,
  input  [7:0]   io_wgt_rd_0_data_bits_0_0,
  input  [7:0]   io_wgt_rd_0_data_bits_0_1,
  input  [7:0]   io_wgt_rd_0_data_bits_0_2,
  input  [7:0]   io_wgt_rd_0_data_bits_0_3,
  input  [7:0]   io_wgt_rd_0_data_bits_0_4,
  input  [7:0]   io_wgt_rd_0_data_bits_0_5,
  input  [7:0]   io_wgt_rd_0_data_bits_0_6,
  input  [7:0]   io_wgt_rd_0_data_bits_0_7,
  input  [7:0]   io_wgt_rd_0_data_bits_0_8,
  input  [7:0]   io_wgt_rd_0_data_bits_0_9,
  input  [7:0]   io_wgt_rd_0_data_bits_0_10,
  input  [7:0]   io_wgt_rd_0_data_bits_0_11,
  input  [7:0]   io_wgt_rd_0_data_bits_0_12,
  input  [7:0]   io_wgt_rd_0_data_bits_0_13,
  input  [7:0]   io_wgt_rd_0_data_bits_0_14,
  input  [7:0]   io_wgt_rd_0_data_bits_0_15,
  input  [7:0]   io_wgt_rd_0_data_bits_1_0,
  input  [7:0]   io_wgt_rd_0_data_bits_1_1,
  input  [7:0]   io_wgt_rd_0_data_bits_1_2,
  input  [7:0]   io_wgt_rd_0_data_bits_1_3,
  input  [7:0]   io_wgt_rd_0_data_bits_1_4,
  input  [7:0]   io_wgt_rd_0_data_bits_1_5,
  input  [7:0]   io_wgt_rd_0_data_bits_1_6,
  input  [7:0]   io_wgt_rd_0_data_bits_1_7,
  input  [7:0]   io_wgt_rd_0_data_bits_1_8,
  input  [7:0]   io_wgt_rd_0_data_bits_1_9,
  input  [7:0]   io_wgt_rd_0_data_bits_1_10,
  input  [7:0]   io_wgt_rd_0_data_bits_1_11,
  input  [7:0]   io_wgt_rd_0_data_bits_1_12,
  input  [7:0]   io_wgt_rd_0_data_bits_1_13,
  input  [7:0]   io_wgt_rd_0_data_bits_1_14,
  input  [7:0]   io_wgt_rd_0_data_bits_1_15,
  input  [7:0]   io_wgt_rd_0_data_bits_2_0,
  input  [7:0]   io_wgt_rd_0_data_bits_2_1,
  input  [7:0]   io_wgt_rd_0_data_bits_2_2,
  input  [7:0]   io_wgt_rd_0_data_bits_2_3,
  input  [7:0]   io_wgt_rd_0_data_bits_2_4,
  input  [7:0]   io_wgt_rd_0_data_bits_2_5,
  input  [7:0]   io_wgt_rd_0_data_bits_2_6,
  input  [7:0]   io_wgt_rd_0_data_bits_2_7,
  input  [7:0]   io_wgt_rd_0_data_bits_2_8,
  input  [7:0]   io_wgt_rd_0_data_bits_2_9,
  input  [7:0]   io_wgt_rd_0_data_bits_2_10,
  input  [7:0]   io_wgt_rd_0_data_bits_2_11,
  input  [7:0]   io_wgt_rd_0_data_bits_2_12,
  input  [7:0]   io_wgt_rd_0_data_bits_2_13,
  input  [7:0]   io_wgt_rd_0_data_bits_2_14,
  input  [7:0]   io_wgt_rd_0_data_bits_2_15,
  input  [7:0]   io_wgt_rd_0_data_bits_3_0,
  input  [7:0]   io_wgt_rd_0_data_bits_3_1,
  input  [7:0]   io_wgt_rd_0_data_bits_3_2,
  input  [7:0]   io_wgt_rd_0_data_bits_3_3,
  input  [7:0]   io_wgt_rd_0_data_bits_3_4,
  input  [7:0]   io_wgt_rd_0_data_bits_3_5,
  input  [7:0]   io_wgt_rd_0_data_bits_3_6,
  input  [7:0]   io_wgt_rd_0_data_bits_3_7,
  input  [7:0]   io_wgt_rd_0_data_bits_3_8,
  input  [7:0]   io_wgt_rd_0_data_bits_3_9,
  input  [7:0]   io_wgt_rd_0_data_bits_3_10,
  input  [7:0]   io_wgt_rd_0_data_bits_3_11,
  input  [7:0]   io_wgt_rd_0_data_bits_3_12,
  input  [7:0]   io_wgt_rd_0_data_bits_3_13,
  input  [7:0]   io_wgt_rd_0_data_bits_3_14,
  input  [7:0]   io_wgt_rd_0_data_bits_3_15,
  input  [7:0]   io_wgt_rd_0_data_bits_4_0,
  input  [7:0]   io_wgt_rd_0_data_bits_4_1,
  input  [7:0]   io_wgt_rd_0_data_bits_4_2,
  input  [7:0]   io_wgt_rd_0_data_bits_4_3,
  input  [7:0]   io_wgt_rd_0_data_bits_4_4,
  input  [7:0]   io_wgt_rd_0_data_bits_4_5,
  input  [7:0]   io_wgt_rd_0_data_bits_4_6,
  input  [7:0]   io_wgt_rd_0_data_bits_4_7,
  input  [7:0]   io_wgt_rd_0_data_bits_4_8,
  input  [7:0]   io_wgt_rd_0_data_bits_4_9,
  input  [7:0]   io_wgt_rd_0_data_bits_4_10,
  input  [7:0]   io_wgt_rd_0_data_bits_4_11,
  input  [7:0]   io_wgt_rd_0_data_bits_4_12,
  input  [7:0]   io_wgt_rd_0_data_bits_4_13,
  input  [7:0]   io_wgt_rd_0_data_bits_4_14,
  input  [7:0]   io_wgt_rd_0_data_bits_4_15,
  input  [7:0]   io_wgt_rd_0_data_bits_5_0,
  input  [7:0]   io_wgt_rd_0_data_bits_5_1,
  input  [7:0]   io_wgt_rd_0_data_bits_5_2,
  input  [7:0]   io_wgt_rd_0_data_bits_5_3,
  input  [7:0]   io_wgt_rd_0_data_bits_5_4,
  input  [7:0]   io_wgt_rd_0_data_bits_5_5,
  input  [7:0]   io_wgt_rd_0_data_bits_5_6,
  input  [7:0]   io_wgt_rd_0_data_bits_5_7,
  input  [7:0]   io_wgt_rd_0_data_bits_5_8,
  input  [7:0]   io_wgt_rd_0_data_bits_5_9,
  input  [7:0]   io_wgt_rd_0_data_bits_5_10,
  input  [7:0]   io_wgt_rd_0_data_bits_5_11,
  input  [7:0]   io_wgt_rd_0_data_bits_5_12,
  input  [7:0]   io_wgt_rd_0_data_bits_5_13,
  input  [7:0]   io_wgt_rd_0_data_bits_5_14,
  input  [7:0]   io_wgt_rd_0_data_bits_5_15,
  input  [7:0]   io_wgt_rd_0_data_bits_6_0,
  input  [7:0]   io_wgt_rd_0_data_bits_6_1,
  input  [7:0]   io_wgt_rd_0_data_bits_6_2,
  input  [7:0]   io_wgt_rd_0_data_bits_6_3,
  input  [7:0]   io_wgt_rd_0_data_bits_6_4,
  input  [7:0]   io_wgt_rd_0_data_bits_6_5,
  input  [7:0]   io_wgt_rd_0_data_bits_6_6,
  input  [7:0]   io_wgt_rd_0_data_bits_6_7,
  input  [7:0]   io_wgt_rd_0_data_bits_6_8,
  input  [7:0]   io_wgt_rd_0_data_bits_6_9,
  input  [7:0]   io_wgt_rd_0_data_bits_6_10,
  input  [7:0]   io_wgt_rd_0_data_bits_6_11,
  input  [7:0]   io_wgt_rd_0_data_bits_6_12,
  input  [7:0]   io_wgt_rd_0_data_bits_6_13,
  input  [7:0]   io_wgt_rd_0_data_bits_6_14,
  input  [7:0]   io_wgt_rd_0_data_bits_6_15,
  input  [7:0]   io_wgt_rd_0_data_bits_7_0,
  input  [7:0]   io_wgt_rd_0_data_bits_7_1,
  input  [7:0]   io_wgt_rd_0_data_bits_7_2,
  input  [7:0]   io_wgt_rd_0_data_bits_7_3,
  input  [7:0]   io_wgt_rd_0_data_bits_7_4,
  input  [7:0]   io_wgt_rd_0_data_bits_7_5,
  input  [7:0]   io_wgt_rd_0_data_bits_7_6,
  input  [7:0]   io_wgt_rd_0_data_bits_7_7,
  input  [7:0]   io_wgt_rd_0_data_bits_7_8,
  input  [7:0]   io_wgt_rd_0_data_bits_7_9,
  input  [7:0]   io_wgt_rd_0_data_bits_7_10,
  input  [7:0]   io_wgt_rd_0_data_bits_7_11,
  input  [7:0]   io_wgt_rd_0_data_bits_7_12,
  input  [7:0]   io_wgt_rd_0_data_bits_7_13,
  input  [7:0]   io_wgt_rd_0_data_bits_7_14,
  input  [7:0]   io_wgt_rd_0_data_bits_7_15,
  input  [7:0]   io_wgt_rd_0_data_bits_8_0,
  input  [7:0]   io_wgt_rd_0_data_bits_8_1,
  input  [7:0]   io_wgt_rd_0_data_bits_8_2,
  input  [7:0]   io_wgt_rd_0_data_bits_8_3,
  input  [7:0]   io_wgt_rd_0_data_bits_8_4,
  input  [7:0]   io_wgt_rd_0_data_bits_8_5,
  input  [7:0]   io_wgt_rd_0_data_bits_8_6,
  input  [7:0]   io_wgt_rd_0_data_bits_8_7,
  input  [7:0]   io_wgt_rd_0_data_bits_8_8,
  input  [7:0]   io_wgt_rd_0_data_bits_8_9,
  input  [7:0]   io_wgt_rd_0_data_bits_8_10,
  input  [7:0]   io_wgt_rd_0_data_bits_8_11,
  input  [7:0]   io_wgt_rd_0_data_bits_8_12,
  input  [7:0]   io_wgt_rd_0_data_bits_8_13,
  input  [7:0]   io_wgt_rd_0_data_bits_8_14,
  input  [7:0]   io_wgt_rd_0_data_bits_8_15,
  input  [7:0]   io_wgt_rd_0_data_bits_9_0,
  input  [7:0]   io_wgt_rd_0_data_bits_9_1,
  input  [7:0]   io_wgt_rd_0_data_bits_9_2,
  input  [7:0]   io_wgt_rd_0_data_bits_9_3,
  input  [7:0]   io_wgt_rd_0_data_bits_9_4,
  input  [7:0]   io_wgt_rd_0_data_bits_9_5,
  input  [7:0]   io_wgt_rd_0_data_bits_9_6,
  input  [7:0]   io_wgt_rd_0_data_bits_9_7,
  input  [7:0]   io_wgt_rd_0_data_bits_9_8,
  input  [7:0]   io_wgt_rd_0_data_bits_9_9,
  input  [7:0]   io_wgt_rd_0_data_bits_9_10,
  input  [7:0]   io_wgt_rd_0_data_bits_9_11,
  input  [7:0]   io_wgt_rd_0_data_bits_9_12,
  input  [7:0]   io_wgt_rd_0_data_bits_9_13,
  input  [7:0]   io_wgt_rd_0_data_bits_9_14,
  input  [7:0]   io_wgt_rd_0_data_bits_9_15,
  input  [7:0]   io_wgt_rd_0_data_bits_10_0,
  input  [7:0]   io_wgt_rd_0_data_bits_10_1,
  input  [7:0]   io_wgt_rd_0_data_bits_10_2,
  input  [7:0]   io_wgt_rd_0_data_bits_10_3,
  input  [7:0]   io_wgt_rd_0_data_bits_10_4,
  input  [7:0]   io_wgt_rd_0_data_bits_10_5,
  input  [7:0]   io_wgt_rd_0_data_bits_10_6,
  input  [7:0]   io_wgt_rd_0_data_bits_10_7,
  input  [7:0]   io_wgt_rd_0_data_bits_10_8,
  input  [7:0]   io_wgt_rd_0_data_bits_10_9,
  input  [7:0]   io_wgt_rd_0_data_bits_10_10,
  input  [7:0]   io_wgt_rd_0_data_bits_10_11,
  input  [7:0]   io_wgt_rd_0_data_bits_10_12,
  input  [7:0]   io_wgt_rd_0_data_bits_10_13,
  input  [7:0]   io_wgt_rd_0_data_bits_10_14,
  input  [7:0]   io_wgt_rd_0_data_bits_10_15,
  input  [7:0]   io_wgt_rd_0_data_bits_11_0,
  input  [7:0]   io_wgt_rd_0_data_bits_11_1,
  input  [7:0]   io_wgt_rd_0_data_bits_11_2,
  input  [7:0]   io_wgt_rd_0_data_bits_11_3,
  input  [7:0]   io_wgt_rd_0_data_bits_11_4,
  input  [7:0]   io_wgt_rd_0_data_bits_11_5,
  input  [7:0]   io_wgt_rd_0_data_bits_11_6,
  input  [7:0]   io_wgt_rd_0_data_bits_11_7,
  input  [7:0]   io_wgt_rd_0_data_bits_11_8,
  input  [7:0]   io_wgt_rd_0_data_bits_11_9,
  input  [7:0]   io_wgt_rd_0_data_bits_11_10,
  input  [7:0]   io_wgt_rd_0_data_bits_11_11,
  input  [7:0]   io_wgt_rd_0_data_bits_11_12,
  input  [7:0]   io_wgt_rd_0_data_bits_11_13,
  input  [7:0]   io_wgt_rd_0_data_bits_11_14,
  input  [7:0]   io_wgt_rd_0_data_bits_11_15,
  input  [7:0]   io_wgt_rd_0_data_bits_12_0,
  input  [7:0]   io_wgt_rd_0_data_bits_12_1,
  input  [7:0]   io_wgt_rd_0_data_bits_12_2,
  input  [7:0]   io_wgt_rd_0_data_bits_12_3,
  input  [7:0]   io_wgt_rd_0_data_bits_12_4,
  input  [7:0]   io_wgt_rd_0_data_bits_12_5,
  input  [7:0]   io_wgt_rd_0_data_bits_12_6,
  input  [7:0]   io_wgt_rd_0_data_bits_12_7,
  input  [7:0]   io_wgt_rd_0_data_bits_12_8,
  input  [7:0]   io_wgt_rd_0_data_bits_12_9,
  input  [7:0]   io_wgt_rd_0_data_bits_12_10,
  input  [7:0]   io_wgt_rd_0_data_bits_12_11,
  input  [7:0]   io_wgt_rd_0_data_bits_12_12,
  input  [7:0]   io_wgt_rd_0_data_bits_12_13,
  input  [7:0]   io_wgt_rd_0_data_bits_12_14,
  input  [7:0]   io_wgt_rd_0_data_bits_12_15,
  input  [7:0]   io_wgt_rd_0_data_bits_13_0,
  input  [7:0]   io_wgt_rd_0_data_bits_13_1,
  input  [7:0]   io_wgt_rd_0_data_bits_13_2,
  input  [7:0]   io_wgt_rd_0_data_bits_13_3,
  input  [7:0]   io_wgt_rd_0_data_bits_13_4,
  input  [7:0]   io_wgt_rd_0_data_bits_13_5,
  input  [7:0]   io_wgt_rd_0_data_bits_13_6,
  input  [7:0]   io_wgt_rd_0_data_bits_13_7,
  input  [7:0]   io_wgt_rd_0_data_bits_13_8,
  input  [7:0]   io_wgt_rd_0_data_bits_13_9,
  input  [7:0]   io_wgt_rd_0_data_bits_13_10,
  input  [7:0]   io_wgt_rd_0_data_bits_13_11,
  input  [7:0]   io_wgt_rd_0_data_bits_13_12,
  input  [7:0]   io_wgt_rd_0_data_bits_13_13,
  input  [7:0]   io_wgt_rd_0_data_bits_13_14,
  input  [7:0]   io_wgt_rd_0_data_bits_13_15,
  input  [7:0]   io_wgt_rd_0_data_bits_14_0,
  input  [7:0]   io_wgt_rd_0_data_bits_14_1,
  input  [7:0]   io_wgt_rd_0_data_bits_14_2,
  input  [7:0]   io_wgt_rd_0_data_bits_14_3,
  input  [7:0]   io_wgt_rd_0_data_bits_14_4,
  input  [7:0]   io_wgt_rd_0_data_bits_14_5,
  input  [7:0]   io_wgt_rd_0_data_bits_14_6,
  input  [7:0]   io_wgt_rd_0_data_bits_14_7,
  input  [7:0]   io_wgt_rd_0_data_bits_14_8,
  input  [7:0]   io_wgt_rd_0_data_bits_14_9,
  input  [7:0]   io_wgt_rd_0_data_bits_14_10,
  input  [7:0]   io_wgt_rd_0_data_bits_14_11,
  input  [7:0]   io_wgt_rd_0_data_bits_14_12,
  input  [7:0]   io_wgt_rd_0_data_bits_14_13,
  input  [7:0]   io_wgt_rd_0_data_bits_14_14,
  input  [7:0]   io_wgt_rd_0_data_bits_14_15,
  input  [7:0]   io_wgt_rd_0_data_bits_15_0,
  input  [7:0]   io_wgt_rd_0_data_bits_15_1,
  input  [7:0]   io_wgt_rd_0_data_bits_15_2,
  input  [7:0]   io_wgt_rd_0_data_bits_15_3,
  input  [7:0]   io_wgt_rd_0_data_bits_15_4,
  input  [7:0]   io_wgt_rd_0_data_bits_15_5,
  input  [7:0]   io_wgt_rd_0_data_bits_15_6,
  input  [7:0]   io_wgt_rd_0_data_bits_15_7,
  input  [7:0]   io_wgt_rd_0_data_bits_15_8,
  input  [7:0]   io_wgt_rd_0_data_bits_15_9,
  input  [7:0]   io_wgt_rd_0_data_bits_15_10,
  input  [7:0]   io_wgt_rd_0_data_bits_15_11,
  input  [7:0]   io_wgt_rd_0_data_bits_15_12,
  input  [7:0]   io_wgt_rd_0_data_bits_15_13,
  input  [7:0]   io_wgt_rd_0_data_bits_15_14,
  input  [7:0]   io_wgt_rd_0_data_bits_15_15,
  input  [7:0]   io_wgt_rd_0_data_bits_16_0,
  input  [7:0]   io_wgt_rd_0_data_bits_16_1,
  input  [7:0]   io_wgt_rd_0_data_bits_16_2,
  input  [7:0]   io_wgt_rd_0_data_bits_16_3,
  input  [7:0]   io_wgt_rd_0_data_bits_16_4,
  input  [7:0]   io_wgt_rd_0_data_bits_16_5,
  input  [7:0]   io_wgt_rd_0_data_bits_16_6,
  input  [7:0]   io_wgt_rd_0_data_bits_16_7,
  input  [7:0]   io_wgt_rd_0_data_bits_16_8,
  input  [7:0]   io_wgt_rd_0_data_bits_16_9,
  input  [7:0]   io_wgt_rd_0_data_bits_16_10,
  input  [7:0]   io_wgt_rd_0_data_bits_16_11,
  input  [7:0]   io_wgt_rd_0_data_bits_16_12,
  input  [7:0]   io_wgt_rd_0_data_bits_16_13,
  input  [7:0]   io_wgt_rd_0_data_bits_16_14,
  input  [7:0]   io_wgt_rd_0_data_bits_16_15,
  input  [7:0]   io_wgt_rd_0_data_bits_17_0,
  input  [7:0]   io_wgt_rd_0_data_bits_17_1,
  input  [7:0]   io_wgt_rd_0_data_bits_17_2,
  input  [7:0]   io_wgt_rd_0_data_bits_17_3,
  input  [7:0]   io_wgt_rd_0_data_bits_17_4,
  input  [7:0]   io_wgt_rd_0_data_bits_17_5,
  input  [7:0]   io_wgt_rd_0_data_bits_17_6,
  input  [7:0]   io_wgt_rd_0_data_bits_17_7,
  input  [7:0]   io_wgt_rd_0_data_bits_17_8,
  input  [7:0]   io_wgt_rd_0_data_bits_17_9,
  input  [7:0]   io_wgt_rd_0_data_bits_17_10,
  input  [7:0]   io_wgt_rd_0_data_bits_17_11,
  input  [7:0]   io_wgt_rd_0_data_bits_17_12,
  input  [7:0]   io_wgt_rd_0_data_bits_17_13,
  input  [7:0]   io_wgt_rd_0_data_bits_17_14,
  input  [7:0]   io_wgt_rd_0_data_bits_17_15,
  input  [7:0]   io_wgt_rd_0_data_bits_18_0,
  input  [7:0]   io_wgt_rd_0_data_bits_18_1,
  input  [7:0]   io_wgt_rd_0_data_bits_18_2,
  input  [7:0]   io_wgt_rd_0_data_bits_18_3,
  input  [7:0]   io_wgt_rd_0_data_bits_18_4,
  input  [7:0]   io_wgt_rd_0_data_bits_18_5,
  input  [7:0]   io_wgt_rd_0_data_bits_18_6,
  input  [7:0]   io_wgt_rd_0_data_bits_18_7,
  input  [7:0]   io_wgt_rd_0_data_bits_18_8,
  input  [7:0]   io_wgt_rd_0_data_bits_18_9,
  input  [7:0]   io_wgt_rd_0_data_bits_18_10,
  input  [7:0]   io_wgt_rd_0_data_bits_18_11,
  input  [7:0]   io_wgt_rd_0_data_bits_18_12,
  input  [7:0]   io_wgt_rd_0_data_bits_18_13,
  input  [7:0]   io_wgt_rd_0_data_bits_18_14,
  input  [7:0]   io_wgt_rd_0_data_bits_18_15,
  input  [7:0]   io_wgt_rd_0_data_bits_19_0,
  input  [7:0]   io_wgt_rd_0_data_bits_19_1,
  input  [7:0]   io_wgt_rd_0_data_bits_19_2,
  input  [7:0]   io_wgt_rd_0_data_bits_19_3,
  input  [7:0]   io_wgt_rd_0_data_bits_19_4,
  input  [7:0]   io_wgt_rd_0_data_bits_19_5,
  input  [7:0]   io_wgt_rd_0_data_bits_19_6,
  input  [7:0]   io_wgt_rd_0_data_bits_19_7,
  input  [7:0]   io_wgt_rd_0_data_bits_19_8,
  input  [7:0]   io_wgt_rd_0_data_bits_19_9,
  input  [7:0]   io_wgt_rd_0_data_bits_19_10,
  input  [7:0]   io_wgt_rd_0_data_bits_19_11,
  input  [7:0]   io_wgt_rd_0_data_bits_19_12,
  input  [7:0]   io_wgt_rd_0_data_bits_19_13,
  input  [7:0]   io_wgt_rd_0_data_bits_19_14,
  input  [7:0]   io_wgt_rd_0_data_bits_19_15,
  input  [7:0]   io_wgt_rd_0_data_bits_20_0,
  input  [7:0]   io_wgt_rd_0_data_bits_20_1,
  input  [7:0]   io_wgt_rd_0_data_bits_20_2,
  input  [7:0]   io_wgt_rd_0_data_bits_20_3,
  input  [7:0]   io_wgt_rd_0_data_bits_20_4,
  input  [7:0]   io_wgt_rd_0_data_bits_20_5,
  input  [7:0]   io_wgt_rd_0_data_bits_20_6,
  input  [7:0]   io_wgt_rd_0_data_bits_20_7,
  input  [7:0]   io_wgt_rd_0_data_bits_20_8,
  input  [7:0]   io_wgt_rd_0_data_bits_20_9,
  input  [7:0]   io_wgt_rd_0_data_bits_20_10,
  input  [7:0]   io_wgt_rd_0_data_bits_20_11,
  input  [7:0]   io_wgt_rd_0_data_bits_20_12,
  input  [7:0]   io_wgt_rd_0_data_bits_20_13,
  input  [7:0]   io_wgt_rd_0_data_bits_20_14,
  input  [7:0]   io_wgt_rd_0_data_bits_20_15,
  input  [7:0]   io_wgt_rd_0_data_bits_21_0,
  input  [7:0]   io_wgt_rd_0_data_bits_21_1,
  input  [7:0]   io_wgt_rd_0_data_bits_21_2,
  input  [7:0]   io_wgt_rd_0_data_bits_21_3,
  input  [7:0]   io_wgt_rd_0_data_bits_21_4,
  input  [7:0]   io_wgt_rd_0_data_bits_21_5,
  input  [7:0]   io_wgt_rd_0_data_bits_21_6,
  input  [7:0]   io_wgt_rd_0_data_bits_21_7,
  input  [7:0]   io_wgt_rd_0_data_bits_21_8,
  input  [7:0]   io_wgt_rd_0_data_bits_21_9,
  input  [7:0]   io_wgt_rd_0_data_bits_21_10,
  input  [7:0]   io_wgt_rd_0_data_bits_21_11,
  input  [7:0]   io_wgt_rd_0_data_bits_21_12,
  input  [7:0]   io_wgt_rd_0_data_bits_21_13,
  input  [7:0]   io_wgt_rd_0_data_bits_21_14,
  input  [7:0]   io_wgt_rd_0_data_bits_21_15,
  input  [7:0]   io_wgt_rd_0_data_bits_22_0,
  input  [7:0]   io_wgt_rd_0_data_bits_22_1,
  input  [7:0]   io_wgt_rd_0_data_bits_22_2,
  input  [7:0]   io_wgt_rd_0_data_bits_22_3,
  input  [7:0]   io_wgt_rd_0_data_bits_22_4,
  input  [7:0]   io_wgt_rd_0_data_bits_22_5,
  input  [7:0]   io_wgt_rd_0_data_bits_22_6,
  input  [7:0]   io_wgt_rd_0_data_bits_22_7,
  input  [7:0]   io_wgt_rd_0_data_bits_22_8,
  input  [7:0]   io_wgt_rd_0_data_bits_22_9,
  input  [7:0]   io_wgt_rd_0_data_bits_22_10,
  input  [7:0]   io_wgt_rd_0_data_bits_22_11,
  input  [7:0]   io_wgt_rd_0_data_bits_22_12,
  input  [7:0]   io_wgt_rd_0_data_bits_22_13,
  input  [7:0]   io_wgt_rd_0_data_bits_22_14,
  input  [7:0]   io_wgt_rd_0_data_bits_22_15,
  input  [7:0]   io_wgt_rd_0_data_bits_23_0,
  input  [7:0]   io_wgt_rd_0_data_bits_23_1,
  input  [7:0]   io_wgt_rd_0_data_bits_23_2,
  input  [7:0]   io_wgt_rd_0_data_bits_23_3,
  input  [7:0]   io_wgt_rd_0_data_bits_23_4,
  input  [7:0]   io_wgt_rd_0_data_bits_23_5,
  input  [7:0]   io_wgt_rd_0_data_bits_23_6,
  input  [7:0]   io_wgt_rd_0_data_bits_23_7,
  input  [7:0]   io_wgt_rd_0_data_bits_23_8,
  input  [7:0]   io_wgt_rd_0_data_bits_23_9,
  input  [7:0]   io_wgt_rd_0_data_bits_23_10,
  input  [7:0]   io_wgt_rd_0_data_bits_23_11,
  input  [7:0]   io_wgt_rd_0_data_bits_23_12,
  input  [7:0]   io_wgt_rd_0_data_bits_23_13,
  input  [7:0]   io_wgt_rd_0_data_bits_23_14,
  input  [7:0]   io_wgt_rd_0_data_bits_23_15,
  input  [7:0]   io_wgt_rd_0_data_bits_24_0,
  input  [7:0]   io_wgt_rd_0_data_bits_24_1,
  input  [7:0]   io_wgt_rd_0_data_bits_24_2,
  input  [7:0]   io_wgt_rd_0_data_bits_24_3,
  input  [7:0]   io_wgt_rd_0_data_bits_24_4,
  input  [7:0]   io_wgt_rd_0_data_bits_24_5,
  input  [7:0]   io_wgt_rd_0_data_bits_24_6,
  input  [7:0]   io_wgt_rd_0_data_bits_24_7,
  input  [7:0]   io_wgt_rd_0_data_bits_24_8,
  input  [7:0]   io_wgt_rd_0_data_bits_24_9,
  input  [7:0]   io_wgt_rd_0_data_bits_24_10,
  input  [7:0]   io_wgt_rd_0_data_bits_24_11,
  input  [7:0]   io_wgt_rd_0_data_bits_24_12,
  input  [7:0]   io_wgt_rd_0_data_bits_24_13,
  input  [7:0]   io_wgt_rd_0_data_bits_24_14,
  input  [7:0]   io_wgt_rd_0_data_bits_24_15,
  input  [7:0]   io_wgt_rd_0_data_bits_25_0,
  input  [7:0]   io_wgt_rd_0_data_bits_25_1,
  input  [7:0]   io_wgt_rd_0_data_bits_25_2,
  input  [7:0]   io_wgt_rd_0_data_bits_25_3,
  input  [7:0]   io_wgt_rd_0_data_bits_25_4,
  input  [7:0]   io_wgt_rd_0_data_bits_25_5,
  input  [7:0]   io_wgt_rd_0_data_bits_25_6,
  input  [7:0]   io_wgt_rd_0_data_bits_25_7,
  input  [7:0]   io_wgt_rd_0_data_bits_25_8,
  input  [7:0]   io_wgt_rd_0_data_bits_25_9,
  input  [7:0]   io_wgt_rd_0_data_bits_25_10,
  input  [7:0]   io_wgt_rd_0_data_bits_25_11,
  input  [7:0]   io_wgt_rd_0_data_bits_25_12,
  input  [7:0]   io_wgt_rd_0_data_bits_25_13,
  input  [7:0]   io_wgt_rd_0_data_bits_25_14,
  input  [7:0]   io_wgt_rd_0_data_bits_25_15,
  input  [7:0]   io_wgt_rd_0_data_bits_26_0,
  input  [7:0]   io_wgt_rd_0_data_bits_26_1,
  input  [7:0]   io_wgt_rd_0_data_bits_26_2,
  input  [7:0]   io_wgt_rd_0_data_bits_26_3,
  input  [7:0]   io_wgt_rd_0_data_bits_26_4,
  input  [7:0]   io_wgt_rd_0_data_bits_26_5,
  input  [7:0]   io_wgt_rd_0_data_bits_26_6,
  input  [7:0]   io_wgt_rd_0_data_bits_26_7,
  input  [7:0]   io_wgt_rd_0_data_bits_26_8,
  input  [7:0]   io_wgt_rd_0_data_bits_26_9,
  input  [7:0]   io_wgt_rd_0_data_bits_26_10,
  input  [7:0]   io_wgt_rd_0_data_bits_26_11,
  input  [7:0]   io_wgt_rd_0_data_bits_26_12,
  input  [7:0]   io_wgt_rd_0_data_bits_26_13,
  input  [7:0]   io_wgt_rd_0_data_bits_26_14,
  input  [7:0]   io_wgt_rd_0_data_bits_26_15,
  input  [7:0]   io_wgt_rd_0_data_bits_27_0,
  input  [7:0]   io_wgt_rd_0_data_bits_27_1,
  input  [7:0]   io_wgt_rd_0_data_bits_27_2,
  input  [7:0]   io_wgt_rd_0_data_bits_27_3,
  input  [7:0]   io_wgt_rd_0_data_bits_27_4,
  input  [7:0]   io_wgt_rd_0_data_bits_27_5,
  input  [7:0]   io_wgt_rd_0_data_bits_27_6,
  input  [7:0]   io_wgt_rd_0_data_bits_27_7,
  input  [7:0]   io_wgt_rd_0_data_bits_27_8,
  input  [7:0]   io_wgt_rd_0_data_bits_27_9,
  input  [7:0]   io_wgt_rd_0_data_bits_27_10,
  input  [7:0]   io_wgt_rd_0_data_bits_27_11,
  input  [7:0]   io_wgt_rd_0_data_bits_27_12,
  input  [7:0]   io_wgt_rd_0_data_bits_27_13,
  input  [7:0]   io_wgt_rd_0_data_bits_27_14,
  input  [7:0]   io_wgt_rd_0_data_bits_27_15,
  input  [7:0]   io_wgt_rd_0_data_bits_28_0,
  input  [7:0]   io_wgt_rd_0_data_bits_28_1,
  input  [7:0]   io_wgt_rd_0_data_bits_28_2,
  input  [7:0]   io_wgt_rd_0_data_bits_28_3,
  input  [7:0]   io_wgt_rd_0_data_bits_28_4,
  input  [7:0]   io_wgt_rd_0_data_bits_28_5,
  input  [7:0]   io_wgt_rd_0_data_bits_28_6,
  input  [7:0]   io_wgt_rd_0_data_bits_28_7,
  input  [7:0]   io_wgt_rd_0_data_bits_28_8,
  input  [7:0]   io_wgt_rd_0_data_bits_28_9,
  input  [7:0]   io_wgt_rd_0_data_bits_28_10,
  input  [7:0]   io_wgt_rd_0_data_bits_28_11,
  input  [7:0]   io_wgt_rd_0_data_bits_28_12,
  input  [7:0]   io_wgt_rd_0_data_bits_28_13,
  input  [7:0]   io_wgt_rd_0_data_bits_28_14,
  input  [7:0]   io_wgt_rd_0_data_bits_28_15,
  input  [7:0]   io_wgt_rd_0_data_bits_29_0,
  input  [7:0]   io_wgt_rd_0_data_bits_29_1,
  input  [7:0]   io_wgt_rd_0_data_bits_29_2,
  input  [7:0]   io_wgt_rd_0_data_bits_29_3,
  input  [7:0]   io_wgt_rd_0_data_bits_29_4,
  input  [7:0]   io_wgt_rd_0_data_bits_29_5,
  input  [7:0]   io_wgt_rd_0_data_bits_29_6,
  input  [7:0]   io_wgt_rd_0_data_bits_29_7,
  input  [7:0]   io_wgt_rd_0_data_bits_29_8,
  input  [7:0]   io_wgt_rd_0_data_bits_29_9,
  input  [7:0]   io_wgt_rd_0_data_bits_29_10,
  input  [7:0]   io_wgt_rd_0_data_bits_29_11,
  input  [7:0]   io_wgt_rd_0_data_bits_29_12,
  input  [7:0]   io_wgt_rd_0_data_bits_29_13,
  input  [7:0]   io_wgt_rd_0_data_bits_29_14,
  input  [7:0]   io_wgt_rd_0_data_bits_29_15,
  input  [7:0]   io_wgt_rd_0_data_bits_30_0,
  input  [7:0]   io_wgt_rd_0_data_bits_30_1,
  input  [7:0]   io_wgt_rd_0_data_bits_30_2,
  input  [7:0]   io_wgt_rd_0_data_bits_30_3,
  input  [7:0]   io_wgt_rd_0_data_bits_30_4,
  input  [7:0]   io_wgt_rd_0_data_bits_30_5,
  input  [7:0]   io_wgt_rd_0_data_bits_30_6,
  input  [7:0]   io_wgt_rd_0_data_bits_30_7,
  input  [7:0]   io_wgt_rd_0_data_bits_30_8,
  input  [7:0]   io_wgt_rd_0_data_bits_30_9,
  input  [7:0]   io_wgt_rd_0_data_bits_30_10,
  input  [7:0]   io_wgt_rd_0_data_bits_30_11,
  input  [7:0]   io_wgt_rd_0_data_bits_30_12,
  input  [7:0]   io_wgt_rd_0_data_bits_30_13,
  input  [7:0]   io_wgt_rd_0_data_bits_30_14,
  input  [7:0]   io_wgt_rd_0_data_bits_30_15,
  input  [7:0]   io_wgt_rd_0_data_bits_31_0,
  input  [7:0]   io_wgt_rd_0_data_bits_31_1,
  input  [7:0]   io_wgt_rd_0_data_bits_31_2,
  input  [7:0]   io_wgt_rd_0_data_bits_31_3,
  input  [7:0]   io_wgt_rd_0_data_bits_31_4,
  input  [7:0]   io_wgt_rd_0_data_bits_31_5,
  input  [7:0]   io_wgt_rd_0_data_bits_31_6,
  input  [7:0]   io_wgt_rd_0_data_bits_31_7,
  input  [7:0]   io_wgt_rd_0_data_bits_31_8,
  input  [7:0]   io_wgt_rd_0_data_bits_31_9,
  input  [7:0]   io_wgt_rd_0_data_bits_31_10,
  input  [7:0]   io_wgt_rd_0_data_bits_31_11,
  input  [7:0]   io_wgt_rd_0_data_bits_31_12,
  input  [7:0]   io_wgt_rd_0_data_bits_31_13,
  input  [7:0]   io_wgt_rd_0_data_bits_31_14,
  input  [7:0]   io_wgt_rd_0_data_bits_31_15,
  output         io_out_wr_0_valid,
  output [6:0]   io_out_wr_0_bits_idx,
  output [7:0]   io_out_wr_0_bits_data_0_0,
  output [7:0]   io_out_wr_0_bits_data_0_1,
  output [7:0]   io_out_wr_0_bits_data_0_2,
  output [7:0]   io_out_wr_0_bits_data_0_3,
  output [7:0]   io_out_wr_0_bits_data_0_4,
  output [7:0]   io_out_wr_0_bits_data_0_5,
  output [7:0]   io_out_wr_0_bits_data_0_6,
  output [7:0]   io_out_wr_0_bits_data_0_7,
  output [7:0]   io_out_wr_0_bits_data_0_8,
  output [7:0]   io_out_wr_0_bits_data_0_9,
  output [7:0]   io_out_wr_0_bits_data_0_10,
  output [7:0]   io_out_wr_0_bits_data_0_11,
  output [7:0]   io_out_wr_0_bits_data_0_12,
  output [7:0]   io_out_wr_0_bits_data_0_13,
  output [7:0]   io_out_wr_0_bits_data_0_14,
  output [7:0]   io_out_wr_0_bits_data_0_15,
  output [7:0]   io_out_wr_0_bits_data_0_16,
  output [7:0]   io_out_wr_0_bits_data_0_17,
  output [7:0]   io_out_wr_0_bits_data_0_18,
  output [7:0]   io_out_wr_0_bits_data_0_19,
  output [7:0]   io_out_wr_0_bits_data_0_20,
  output [7:0]   io_out_wr_0_bits_data_0_21,
  output [7:0]   io_out_wr_0_bits_data_0_22,
  output [7:0]   io_out_wr_0_bits_data_0_23,
  output [7:0]   io_out_wr_0_bits_data_0_24,
  output [7:0]   io_out_wr_0_bits_data_0_25,
  output [7:0]   io_out_wr_0_bits_data_0_26,
  output [7:0]   io_out_wr_0_bits_data_0_27,
  output [7:0]   io_out_wr_0_bits_data_0_28,
  output [7:0]   io_out_wr_0_bits_data_0_29,
  output [7:0]   io_out_wr_0_bits_data_0_30,
  output [7:0]   io_out_wr_0_bits_data_0_31,
  output         io_finish,
  output         io_acc_wr_event
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  s_0_clock; // @[Compute.scala 58:11]
  wire  s_0_reset; // @[Compute.scala 58:11]
  wire  s_0_io_spost; // @[Compute.scala 58:11]
  wire  s_0_io_swait; // @[Compute.scala 58:11]
  wire  s_0_io_sready; // @[Compute.scala 58:11]
  wire  s_1_clock; // @[Compute.scala 58:11]
  wire  s_1_reset; // @[Compute.scala 58:11]
  wire  s_1_io_spost; // @[Compute.scala 58:11]
  wire  s_1_io_swait; // @[Compute.scala 58:11]
  wire  s_1_io_sready; // @[Compute.scala 58:11]
  wire  loadUop_clock; // @[Compute.scala 61:23]
  wire  loadUop_reset; // @[Compute.scala 61:23]
  wire  loadUop_io_start; // @[Compute.scala 61:23]
  wire  loadUop_io_done; // @[Compute.scala 61:23]
  wire [127:0] loadUop_io_inst; // @[Compute.scala 61:23]
  wire [31:0] loadUop_io_baddr; // @[Compute.scala 61:23]
  wire  loadUop_io_vme_rd_cmd_ready; // @[Compute.scala 61:23]
  wire  loadUop_io_vme_rd_cmd_valid; // @[Compute.scala 61:23]
  wire [31:0] loadUop_io_vme_rd_cmd_bits_addr; // @[Compute.scala 61:23]
  wire [3:0] loadUop_io_vme_rd_cmd_bits_len; // @[Compute.scala 61:23]
  wire [20:0] loadUop_io_vme_rd_cmd_bits_tag; // @[Compute.scala 61:23]
  wire  loadUop_io_vme_rd_data_valid; // @[Compute.scala 61:23]
  wire [63:0] loadUop_io_vme_rd_data_bits_data; // @[Compute.scala 61:23]
  wire [20:0] loadUop_io_vme_rd_data_bits_tag; // @[Compute.scala 61:23]
  wire  loadUop_io_vme_rd_data_bits_last; // @[Compute.scala 61:23]
  wire  loadUop_io_uop_idx_valid; // @[Compute.scala 61:23]
  wire [6:0] loadUop_io_uop_idx_bits; // @[Compute.scala 61:23]
  wire  loadUop_io_uop_data_valid; // @[Compute.scala 61:23]
  wire [9:0] loadUop_io_uop_data_bits_u2; // @[Compute.scala 61:23]
  wire [10:0] loadUop_io_uop_data_bits_u1; // @[Compute.scala 61:23]
  wire [10:0] loadUop_io_uop_data_bits_u0; // @[Compute.scala 61:23]
  wire  tensorAcc_clock; // @[Compute.scala 62:25]
  wire  tensorAcc_reset; // @[Compute.scala 62:25]
  wire  tensorAcc_io_start; // @[Compute.scala 62:25]
  wire  tensorAcc_io_done; // @[Compute.scala 62:25]
  wire [127:0] tensorAcc_io_inst; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_baddr; // @[Compute.scala 62:25]
  wire  tensorAcc_io_vme_rd_cmd_ready; // @[Compute.scala 62:25]
  wire  tensorAcc_io_vme_rd_cmd_valid; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_vme_rd_cmd_bits_addr; // @[Compute.scala 62:25]
  wire [3:0] tensorAcc_io_vme_rd_cmd_bits_len; // @[Compute.scala 62:25]
  wire [20:0] tensorAcc_io_vme_rd_cmd_bits_tag; // @[Compute.scala 62:25]
  wire  tensorAcc_io_vme_rd_data_valid; // @[Compute.scala 62:25]
  wire [63:0] tensorAcc_io_vme_rd_data_bits_data; // @[Compute.scala 62:25]
  wire [20:0] tensorAcc_io_vme_rd_data_bits_tag; // @[Compute.scala 62:25]
  wire  tensorAcc_io_tensor_rd_0_idx_valid; // @[Compute.scala 62:25]
  wire [6:0] tensorAcc_io_tensor_rd_0_idx_bits; // @[Compute.scala 62:25]
  wire  tensorAcc_io_tensor_rd_0_data_valid; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_0; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_1; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_2; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_3; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_4; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_5; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_6; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_7; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_8; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_9; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_10; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_11; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_12; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_13; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_14; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_15; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_16; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_17; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_18; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_19; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_20; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_21; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_22; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_23; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_24; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_25; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_26; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_27; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_28; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_29; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_30; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_rd_0_data_bits_0_31; // @[Compute.scala 62:25]
  wire  tensorAcc_io_tensor_wr_0_valid; // @[Compute.scala 62:25]
  wire [6:0] tensorAcc_io_tensor_wr_0_bits_idx; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_0; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_1; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_2; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_3; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_4; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_5; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_6; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_7; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_8; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_9; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_10; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_11; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_12; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_13; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_14; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_15; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_16; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_17; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_18; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_19; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_20; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_21; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_22; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_23; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_24; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_25; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_26; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_27; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_28; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_29; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_30; // @[Compute.scala 62:25]
  wire [31:0] tensorAcc_io_tensor_wr_0_bits_data_0_31; // @[Compute.scala 62:25]
  wire  tensorGemm_clock; // @[Compute.scala 63:26]
  wire  tensorGemm_reset; // @[Compute.scala 63:26]
  wire  tensorGemm_io_start; // @[Compute.scala 63:26]
  wire  tensorGemm_io_done; // @[Compute.scala 63:26]
  wire [9:0] tensorGemm_io_dec_wgt_1; // @[Compute.scala 63:26]
  wire [9:0] tensorGemm_io_dec_wgt_0; // @[Compute.scala 63:26]
  wire [10:0] tensorGemm_io_dec_inp_1; // @[Compute.scala 63:26]
  wire [10:0] tensorGemm_io_dec_inp_0; // @[Compute.scala 63:26]
  wire [10:0] tensorGemm_io_dec_acc_1; // @[Compute.scala 63:26]
  wire [10:0] tensorGemm_io_dec_acc_0; // @[Compute.scala 63:26]
  wire  tensorGemm_io_dec_empty_0; // @[Compute.scala 63:26]
  wire [13:0] tensorGemm_io_dec_lp_1; // @[Compute.scala 63:26]
  wire [13:0] tensorGemm_io_dec_lp_0; // @[Compute.scala 63:26]
  wire [13:0] tensorGemm_io_dec_uop_end; // @[Compute.scala 63:26]
  wire [12:0] tensorGemm_io_dec_uop_begin; // @[Compute.scala 63:26]
  wire  tensorGemm_io_dec_reset; // @[Compute.scala 63:26]
  wire  tensorGemm_io_dec_push_next; // @[Compute.scala 63:26]
  wire  tensorGemm_io_dec_push_prev; // @[Compute.scala 63:26]
  wire  tensorGemm_io_dec_pop_next; // @[Compute.scala 63:26]
  wire  tensorGemm_io_dec_pop_prev; // @[Compute.scala 63:26]
  wire [2:0] tensorGemm_io_dec_op; // @[Compute.scala 63:26]
  wire  tensorGemm_io_uop_idx_valid; // @[Compute.scala 63:26]
  wire [6:0] tensorGemm_io_uop_idx_bits; // @[Compute.scala 63:26]
  wire  tensorGemm_io_uop_data_valid; // @[Compute.scala 63:26]
  wire [9:0] tensorGemm_io_uop_data_bits_u2; // @[Compute.scala 63:26]
  wire [10:0] tensorGemm_io_uop_data_bits_u1; // @[Compute.scala 63:26]
  wire [10:0] tensorGemm_io_uop_data_bits_u0; // @[Compute.scala 63:26]
  wire  tensorGemm_io_inp_rd_0_idx_valid; // @[Compute.scala 63:26]
  wire [6:0] tensorGemm_io_inp_rd_0_idx_bits; // @[Compute.scala 63:26]
  wire  tensorGemm_io_inp_rd_0_data_valid; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_inp_rd_0_data_bits_0_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_inp_rd_0_data_bits_0_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_inp_rd_0_data_bits_0_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_inp_rd_0_data_bits_0_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_inp_rd_0_data_bits_0_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_inp_rd_0_data_bits_0_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_inp_rd_0_data_bits_0_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_inp_rd_0_data_bits_0_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_inp_rd_0_data_bits_0_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_inp_rd_0_data_bits_0_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_inp_rd_0_data_bits_0_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_inp_rd_0_data_bits_0_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_inp_rd_0_data_bits_0_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_inp_rd_0_data_bits_0_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_inp_rd_0_data_bits_0_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_inp_rd_0_data_bits_0_15; // @[Compute.scala 63:26]
  wire  tensorGemm_io_wgt_rd_0_idx_valid; // @[Compute.scala 63:26]
  wire [5:0] tensorGemm_io_wgt_rd_0_idx_bits; // @[Compute.scala 63:26]
  wire  tensorGemm_io_wgt_rd_0_data_valid; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_0_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_0_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_0_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_0_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_0_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_0_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_0_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_0_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_0_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_0_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_0_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_0_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_0_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_0_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_0_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_0_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_1_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_1_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_1_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_1_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_1_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_1_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_1_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_1_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_1_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_1_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_1_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_1_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_1_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_1_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_1_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_1_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_2_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_2_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_2_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_2_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_2_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_2_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_2_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_2_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_2_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_2_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_2_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_2_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_2_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_2_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_2_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_2_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_3_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_3_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_3_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_3_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_3_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_3_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_3_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_3_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_3_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_3_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_3_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_3_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_3_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_3_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_3_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_3_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_4_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_4_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_4_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_4_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_4_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_4_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_4_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_4_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_4_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_4_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_4_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_4_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_4_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_4_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_4_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_4_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_5_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_5_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_5_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_5_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_5_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_5_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_5_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_5_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_5_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_5_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_5_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_5_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_5_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_5_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_5_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_5_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_6_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_6_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_6_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_6_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_6_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_6_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_6_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_6_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_6_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_6_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_6_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_6_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_6_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_6_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_6_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_6_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_7_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_7_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_7_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_7_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_7_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_7_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_7_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_7_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_7_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_7_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_7_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_7_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_7_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_7_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_7_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_7_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_8_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_8_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_8_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_8_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_8_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_8_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_8_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_8_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_8_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_8_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_8_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_8_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_8_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_8_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_8_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_8_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_9_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_9_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_9_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_9_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_9_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_9_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_9_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_9_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_9_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_9_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_9_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_9_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_9_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_9_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_9_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_9_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_10_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_10_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_10_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_10_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_10_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_10_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_10_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_10_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_10_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_10_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_10_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_10_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_10_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_10_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_10_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_10_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_11_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_11_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_11_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_11_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_11_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_11_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_11_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_11_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_11_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_11_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_11_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_11_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_11_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_11_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_11_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_11_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_12_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_12_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_12_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_12_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_12_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_12_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_12_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_12_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_12_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_12_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_12_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_12_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_12_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_12_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_12_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_12_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_13_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_13_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_13_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_13_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_13_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_13_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_13_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_13_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_13_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_13_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_13_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_13_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_13_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_13_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_13_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_13_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_14_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_14_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_14_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_14_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_14_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_14_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_14_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_14_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_14_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_14_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_14_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_14_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_14_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_14_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_14_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_14_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_15_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_15_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_15_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_15_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_15_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_15_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_15_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_15_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_15_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_15_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_15_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_15_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_15_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_15_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_15_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_15_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_16_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_16_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_16_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_16_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_16_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_16_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_16_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_16_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_16_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_16_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_16_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_16_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_16_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_16_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_16_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_16_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_17_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_17_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_17_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_17_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_17_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_17_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_17_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_17_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_17_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_17_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_17_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_17_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_17_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_17_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_17_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_17_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_18_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_18_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_18_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_18_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_18_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_18_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_18_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_18_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_18_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_18_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_18_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_18_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_18_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_18_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_18_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_18_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_19_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_19_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_19_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_19_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_19_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_19_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_19_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_19_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_19_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_19_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_19_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_19_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_19_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_19_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_19_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_19_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_20_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_20_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_20_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_20_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_20_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_20_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_20_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_20_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_20_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_20_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_20_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_20_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_20_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_20_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_20_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_20_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_21_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_21_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_21_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_21_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_21_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_21_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_21_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_21_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_21_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_21_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_21_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_21_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_21_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_21_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_21_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_21_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_22_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_22_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_22_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_22_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_22_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_22_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_22_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_22_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_22_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_22_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_22_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_22_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_22_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_22_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_22_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_22_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_23_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_23_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_23_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_23_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_23_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_23_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_23_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_23_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_23_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_23_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_23_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_23_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_23_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_23_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_23_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_23_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_24_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_24_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_24_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_24_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_24_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_24_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_24_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_24_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_24_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_24_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_24_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_24_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_24_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_24_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_24_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_24_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_25_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_25_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_25_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_25_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_25_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_25_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_25_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_25_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_25_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_25_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_25_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_25_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_25_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_25_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_25_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_25_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_26_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_26_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_26_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_26_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_26_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_26_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_26_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_26_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_26_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_26_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_26_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_26_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_26_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_26_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_26_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_26_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_27_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_27_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_27_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_27_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_27_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_27_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_27_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_27_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_27_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_27_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_27_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_27_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_27_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_27_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_27_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_27_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_28_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_28_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_28_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_28_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_28_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_28_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_28_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_28_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_28_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_28_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_28_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_28_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_28_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_28_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_28_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_28_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_29_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_29_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_29_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_29_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_29_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_29_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_29_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_29_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_29_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_29_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_29_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_29_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_29_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_29_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_29_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_29_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_30_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_30_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_30_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_30_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_30_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_30_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_30_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_30_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_30_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_30_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_30_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_30_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_30_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_30_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_30_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_30_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_31_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_31_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_31_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_31_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_31_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_31_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_31_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_31_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_31_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_31_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_31_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_31_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_31_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_31_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_31_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_wgt_rd_0_data_bits_31_15; // @[Compute.scala 63:26]
  wire  tensorGemm_io_acc_rd_0_idx_valid; // @[Compute.scala 63:26]
  wire [6:0] tensorGemm_io_acc_rd_0_idx_bits; // @[Compute.scala 63:26]
  wire  tensorGemm_io_acc_rd_0_data_valid; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_0; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_1; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_2; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_3; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_4; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_5; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_6; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_7; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_8; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_9; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_10; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_11; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_12; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_13; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_14; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_15; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_16; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_17; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_18; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_19; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_20; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_21; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_22; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_23; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_24; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_25; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_26; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_27; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_28; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_29; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_30; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_rd_0_data_bits_0_31; // @[Compute.scala 63:26]
  wire  tensorGemm_io_acc_wr_0_valid; // @[Compute.scala 63:26]
  wire [6:0] tensorGemm_io_acc_wr_0_bits_idx; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_0; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_1; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_2; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_3; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_4; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_5; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_6; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_7; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_8; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_9; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_10; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_11; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_12; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_13; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_14; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_15; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_16; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_17; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_18; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_19; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_20; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_21; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_22; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_23; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_24; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_25; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_26; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_27; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_28; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_29; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_30; // @[Compute.scala 63:26]
  wire [31:0] tensorGemm_io_acc_wr_0_bits_data_0_31; // @[Compute.scala 63:26]
  wire  tensorGemm_io_out_rd_0_data_valid; // @[Compute.scala 63:26]
  wire  tensorGemm_io_out_wr_0_valid; // @[Compute.scala 63:26]
  wire [6:0] tensorGemm_io_out_wr_0_bits_idx; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_0; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_1; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_2; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_3; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_4; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_5; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_6; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_7; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_8; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_9; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_10; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_11; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_12; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_13; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_14; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_15; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_16; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_17; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_18; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_19; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_20; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_21; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_22; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_23; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_24; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_25; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_26; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_27; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_28; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_29; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_30; // @[Compute.scala 63:26]
  wire [7:0] tensorGemm_io_out_wr_0_bits_data_0_31; // @[Compute.scala 63:26]
  wire  tensorAlu_clock; // @[Compute.scala 64:25]
  wire  tensorAlu_reset; // @[Compute.scala 64:25]
  wire  tensorAlu_io_start; // @[Compute.scala 64:25]
  wire  tensorAlu_io_done; // @[Compute.scala 64:25]
  wire [15:0] tensorAlu_io_dec_alu_imm; // @[Compute.scala 64:25]
  wire  tensorAlu_io_dec_alu_use_imm; // @[Compute.scala 64:25]
  wire [2:0] tensorAlu_io_dec_alu_op; // @[Compute.scala 64:25]
  wire [10:0] tensorAlu_io_dec_src_1; // @[Compute.scala 64:25]
  wire [10:0] tensorAlu_io_dec_src_0; // @[Compute.scala 64:25]
  wire [10:0] tensorAlu_io_dec_dst_1; // @[Compute.scala 64:25]
  wire [10:0] tensorAlu_io_dec_dst_0; // @[Compute.scala 64:25]
  wire [13:0] tensorAlu_io_dec_lp_1; // @[Compute.scala 64:25]
  wire [13:0] tensorAlu_io_dec_lp_0; // @[Compute.scala 64:25]
  wire [13:0] tensorAlu_io_dec_uop_end; // @[Compute.scala 64:25]
  wire [12:0] tensorAlu_io_dec_uop_begin; // @[Compute.scala 64:25]
  wire  tensorAlu_io_uop_idx_valid; // @[Compute.scala 64:25]
  wire [6:0] tensorAlu_io_uop_idx_bits; // @[Compute.scala 64:25]
  wire [9:0] tensorAlu_io_uop_data_bits_u2; // @[Compute.scala 64:25]
  wire [10:0] tensorAlu_io_uop_data_bits_u1; // @[Compute.scala 64:25]
  wire [10:0] tensorAlu_io_uop_data_bits_u0; // @[Compute.scala 64:25]
  wire  tensorAlu_io_acc_rd_0_idx_valid; // @[Compute.scala 64:25]
  wire [6:0] tensorAlu_io_acc_rd_0_idx_bits; // @[Compute.scala 64:25]
  wire  tensorAlu_io_acc_rd_0_data_valid; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_0; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_1; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_2; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_3; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_4; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_5; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_6; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_7; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_8; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_9; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_10; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_11; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_12; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_13; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_14; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_15; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_16; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_17; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_18; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_19; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_20; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_21; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_22; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_23; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_24; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_25; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_26; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_27; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_28; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_29; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_30; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_rd_0_data_bits_0_31; // @[Compute.scala 64:25]
  wire  tensorAlu_io_acc_wr_0_valid; // @[Compute.scala 64:25]
  wire [6:0] tensorAlu_io_acc_wr_0_bits_idx; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_0; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_1; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_2; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_3; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_4; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_5; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_6; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_7; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_8; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_9; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_10; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_11; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_12; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_13; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_14; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_15; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_16; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_17; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_18; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_19; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_20; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_21; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_22; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_23; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_24; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_25; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_26; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_27; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_28; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_29; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_30; // @[Compute.scala 64:25]
  wire [31:0] tensorAlu_io_acc_wr_0_bits_data_0_31; // @[Compute.scala 64:25]
  wire  tensorAlu_io_out_rd_0_data_valid; // @[Compute.scala 64:25]
  wire  tensorAlu_io_out_wr_0_valid; // @[Compute.scala 64:25]
  wire [6:0] tensorAlu_io_out_wr_0_bits_idx; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_0; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_1; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_2; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_3; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_4; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_5; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_6; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_7; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_8; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_9; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_10; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_11; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_12; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_13; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_14; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_15; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_16; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_17; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_18; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_19; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_20; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_21; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_22; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_23; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_24; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_25; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_26; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_27; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_28; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_29; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_30; // @[Compute.scala 64:25]
  wire [7:0] tensorAlu_io_out_wr_0_bits_data_0_31; // @[Compute.scala 64:25]
  wire  inst_q_clock; // @[Compute.scala 69:22]
  wire  inst_q_reset; // @[Compute.scala 69:22]
  wire  inst_q_io_enq_ready; // @[Compute.scala 69:22]
  wire  inst_q_io_enq_valid; // @[Compute.scala 69:22]
  wire [127:0] inst_q_io_enq_bits; // @[Compute.scala 69:22]
  wire  inst_q_io_deq_ready; // @[Compute.scala 69:22]
  wire  inst_q_io_deq_valid; // @[Compute.scala 69:22]
  wire [127:0] inst_q_io_deq_bits; // @[Compute.scala 69:22]
  wire [127:0] dec_io_inst; // @[Compute.scala 72:19]
  wire  dec_io_push_next; // @[Compute.scala 72:19]
  wire  dec_io_push_prev; // @[Compute.scala 72:19]
  wire  dec_io_pop_next; // @[Compute.scala 72:19]
  wire  dec_io_pop_prev; // @[Compute.scala 72:19]
  wire  dec_io_isLoadAcc; // @[Compute.scala 72:19]
  wire  dec_io_isLoadUop; // @[Compute.scala 72:19]
  wire  dec_io_isSync; // @[Compute.scala 72:19]
  wire  dec_io_isAlu; // @[Compute.scala 72:19]
  wire  dec_io_isGemm; // @[Compute.scala 72:19]
  wire  dec_io_isFinish; // @[Compute.scala 72:19]
  reg [1:0] state; // @[Compute.scala 55:22]
  wire [4:0] inst_type = {dec_io_isFinish,dec_io_isAlu,dec_io_isGemm,dec_io_isLoadAcc,dec_io_isLoadUop}; // @[Cat.scala 31:58]
  wire  _sprev_T = dec_io_pop_prev ? s_0_io_sready : 1'h1; // @[Compute.scala 82:40]
  wire  sprev = inst_q_io_deq_valid & _sprev_T; // @[Compute.scala 82:35]
  wire  _snext_T = dec_io_pop_next ? s_1_io_sready : 1'h1; // @[Compute.scala 83:40]
  wire  snext = inst_q_io_deq_valid & _snext_T; // @[Compute.scala 83:35]
  wire  start = snext & sprev; // @[Compute.scala 84:21]
  wire  _done_T_3 = 5'h2 == inst_type ? tensorAcc_io_done : 5'h1 == inst_type & loadUop_io_done; // @[Mux.scala 81:58]
  wire  _done_T_5 = 5'h4 == inst_type ? tensorGemm_io_done : _done_T_3; // @[Mux.scala 81:58]
  wire  _done_T_7 = 5'h8 == inst_type ? tensorAlu_io_done : _done_T_5; // @[Mux.scala 81:58]
  wire  done = 5'h10 == inst_type | _done_T_7; // @[Mux.scala 81:58]
  wire [1:0] _GEN_0 = |inst_type ? 2'h2 : state; // @[Compute.scala 104:35 105:17 55:22]
  wire [1:0] _GEN_3 = done ? 2'h0 : state; // @[Compute.scala 113:18 114:15 55:22]
  wire  _inst_q_io_deq_ready_T_1 = state == 2'h2 & done; // @[Compute.scala 121:42]
  wire  _inst_q_io_deq_ready_T_3 = state == 2'h2 & done | state == 2'h1; // @[Compute.scala 121:50]
  wire  _loadUop_io_start_T_1 = state == 2'h0 & start; // @[Compute.scala 124:39]
  wire  _T_8 = ~reset; // @[Compute.scala 129:9]
  reg  tensorAcc_io_tensor_rd_0_idx_REG; // @[Compute.scala 150:14]
  reg  tensorAcc_io_tensor_wr_0_REG; // @[Compute.scala 154:14]
  reg  tensorGemm_io_start_REG; // @[Compute.scala 162:33]
  wire [127:0] _tensorGemm_io_dec_WIRE_1 = inst_q_io_deq_bits;
  reg  tensorGemm_io_acc_rd_0_data_valid_REG; // @[Compute.scala 170:55]
  reg  tensorAlu_io_start_REG; // @[Compute.scala 180:32]
  reg  tensorAlu_io_acc_rd_0_data_valid_REG; // @[Compute.scala 186:55]
  reg  io_out_wr_0_valid_REG; // @[Compute.scala 208:12]
  reg  io_out_wr_0_bits_idx_REG; // @[Compute.scala 210:12]
  reg  outDataBits_0_REG; // @[Compute.scala 221:14]
  wire [63:0] srcGemFlat_hi_lo = {tensorGemm_io_out_wr_0_bits_data_0_23,tensorGemm_io_out_wr_0_bits_data_0_22,
    tensorGemm_io_out_wr_0_bits_data_0_21,tensorGemm_io_out_wr_0_bits_data_0_20,tensorGemm_io_out_wr_0_bits_data_0_19,
    tensorGemm_io_out_wr_0_bits_data_0_18,tensorGemm_io_out_wr_0_bits_data_0_17,tensorGemm_io_out_wr_0_bits_data_0_16}; // @[Compute.scala 219:56]
  wire [63:0] srcGemFlat_lo_lo = {tensorGemm_io_out_wr_0_bits_data_0_7,tensorGemm_io_out_wr_0_bits_data_0_6,
    tensorGemm_io_out_wr_0_bits_data_0_5,tensorGemm_io_out_wr_0_bits_data_0_4,tensorGemm_io_out_wr_0_bits_data_0_3,
    tensorGemm_io_out_wr_0_bits_data_0_2,tensorGemm_io_out_wr_0_bits_data_0_1,tensorGemm_io_out_wr_0_bits_data_0_0}; // @[Compute.scala 219:56]
  wire [127:0] srcGemFlat_lo = {tensorGemm_io_out_wr_0_bits_data_0_15,tensorGemm_io_out_wr_0_bits_data_0_14,
    tensorGemm_io_out_wr_0_bits_data_0_13,tensorGemm_io_out_wr_0_bits_data_0_12,tensorGemm_io_out_wr_0_bits_data_0_11,
    tensorGemm_io_out_wr_0_bits_data_0_10,tensorGemm_io_out_wr_0_bits_data_0_9,tensorGemm_io_out_wr_0_bits_data_0_8,
    srcGemFlat_lo_lo}; // @[Compute.scala 219:56]
  wire [255:0] srcGemFlat = {tensorGemm_io_out_wr_0_bits_data_0_31,tensorGemm_io_out_wr_0_bits_data_0_30,
    tensorGemm_io_out_wr_0_bits_data_0_29,tensorGemm_io_out_wr_0_bits_data_0_28,tensorGemm_io_out_wr_0_bits_data_0_27,
    tensorGemm_io_out_wr_0_bits_data_0_26,tensorGemm_io_out_wr_0_bits_data_0_25,tensorGemm_io_out_wr_0_bits_data_0_24,
    srcGemFlat_hi_lo,srcGemFlat_lo}; // @[Compute.scala 219:56]
  wire [63:0] srcAluFlat_hi_lo = {tensorAlu_io_out_wr_0_bits_data_0_23,tensorAlu_io_out_wr_0_bits_data_0_22,
    tensorAlu_io_out_wr_0_bits_data_0_21,tensorAlu_io_out_wr_0_bits_data_0_20,tensorAlu_io_out_wr_0_bits_data_0_19,
    tensorAlu_io_out_wr_0_bits_data_0_18,tensorAlu_io_out_wr_0_bits_data_0_17,tensorAlu_io_out_wr_0_bits_data_0_16}; // @[Compute.scala 218:55]
  wire [63:0] srcAluFlat_lo_lo = {tensorAlu_io_out_wr_0_bits_data_0_7,tensorAlu_io_out_wr_0_bits_data_0_6,
    tensorAlu_io_out_wr_0_bits_data_0_5,tensorAlu_io_out_wr_0_bits_data_0_4,tensorAlu_io_out_wr_0_bits_data_0_3,
    tensorAlu_io_out_wr_0_bits_data_0_2,tensorAlu_io_out_wr_0_bits_data_0_1,tensorAlu_io_out_wr_0_bits_data_0_0}; // @[Compute.scala 218:55]
  wire [127:0] srcAluFlat_lo = {tensorAlu_io_out_wr_0_bits_data_0_15,tensorAlu_io_out_wr_0_bits_data_0_14,
    tensorAlu_io_out_wr_0_bits_data_0_13,tensorAlu_io_out_wr_0_bits_data_0_12,tensorAlu_io_out_wr_0_bits_data_0_11,
    tensorAlu_io_out_wr_0_bits_data_0_10,tensorAlu_io_out_wr_0_bits_data_0_9,tensorAlu_io_out_wr_0_bits_data_0_8,
    srcAluFlat_lo_lo}; // @[Compute.scala 218:55]
  wire [255:0] srcAluFlat = {tensorAlu_io_out_wr_0_bits_data_0_31,tensorAlu_io_out_wr_0_bits_data_0_30,
    tensorAlu_io_out_wr_0_bits_data_0_29,tensorAlu_io_out_wr_0_bits_data_0_28,tensorAlu_io_out_wr_0_bits_data_0_27,
    tensorAlu_io_out_wr_0_bits_data_0_26,tensorAlu_io_out_wr_0_bits_data_0_25,tensorAlu_io_out_wr_0_bits_data_0_24,
    srcAluFlat_hi_lo,srcAluFlat_lo}; // @[Compute.scala 218:55]
  wire [255:0] outDataBits_0 = outDataBits_0_REG ? srcGemFlat : srcAluFlat; // @[Compute.scala 220:28]
  Semaphore s_0 ( // @[Compute.scala 58:11]
    .clock(s_0_clock),
    .reset(s_0_reset),
    .io_spost(s_0_io_spost),
    .io_swait(s_0_io_swait),
    .io_sready(s_0_io_sready)
  );
  Semaphore s_1 ( // @[Compute.scala 58:11]
    .clock(s_1_clock),
    .reset(s_1_reset),
    .io_spost(s_1_io_spost),
    .io_swait(s_1_io_swait),
    .io_sready(s_1_io_sready)
  );
  LoadUopTop loadUop ( // @[Compute.scala 61:23]
    .clock(loadUop_clock),
    .reset(loadUop_reset),
    .io_start(loadUop_io_start),
    .io_done(loadUop_io_done),
    .io_inst(loadUop_io_inst),
    .io_baddr(loadUop_io_baddr),
    .io_vme_rd_cmd_ready(loadUop_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(loadUop_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(loadUop_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(loadUop_io_vme_rd_cmd_bits_len),
    .io_vme_rd_cmd_bits_tag(loadUop_io_vme_rd_cmd_bits_tag),
    .io_vme_rd_data_valid(loadUop_io_vme_rd_data_valid),
    .io_vme_rd_data_bits_data(loadUop_io_vme_rd_data_bits_data),
    .io_vme_rd_data_bits_tag(loadUop_io_vme_rd_data_bits_tag),
    .io_vme_rd_data_bits_last(loadUop_io_vme_rd_data_bits_last),
    .io_uop_idx_valid(loadUop_io_uop_idx_valid),
    .io_uop_idx_bits(loadUop_io_uop_idx_bits),
    .io_uop_data_valid(loadUop_io_uop_data_valid),
    .io_uop_data_bits_u2(loadUop_io_uop_data_bits_u2),
    .io_uop_data_bits_u1(loadUop_io_uop_data_bits_u1),
    .io_uop_data_bits_u0(loadUop_io_uop_data_bits_u0)
  );
  TensorLoadAcc tensorAcc ( // @[Compute.scala 62:25]
    .clock(tensorAcc_clock),
    .reset(tensorAcc_reset),
    .io_start(tensorAcc_io_start),
    .io_done(tensorAcc_io_done),
    .io_inst(tensorAcc_io_inst),
    .io_baddr(tensorAcc_io_baddr),
    .io_vme_rd_cmd_ready(tensorAcc_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(tensorAcc_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(tensorAcc_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(tensorAcc_io_vme_rd_cmd_bits_len),
    .io_vme_rd_cmd_bits_tag(tensorAcc_io_vme_rd_cmd_bits_tag),
    .io_vme_rd_data_valid(tensorAcc_io_vme_rd_data_valid),
    .io_vme_rd_data_bits_data(tensorAcc_io_vme_rd_data_bits_data),
    .io_vme_rd_data_bits_tag(tensorAcc_io_vme_rd_data_bits_tag),
    .io_tensor_rd_0_idx_valid(tensorAcc_io_tensor_rd_0_idx_valid),
    .io_tensor_rd_0_idx_bits(tensorAcc_io_tensor_rd_0_idx_bits),
    .io_tensor_rd_0_data_valid(tensorAcc_io_tensor_rd_0_data_valid),
    .io_tensor_rd_0_data_bits_0_0(tensorAcc_io_tensor_rd_0_data_bits_0_0),
    .io_tensor_rd_0_data_bits_0_1(tensorAcc_io_tensor_rd_0_data_bits_0_1),
    .io_tensor_rd_0_data_bits_0_2(tensorAcc_io_tensor_rd_0_data_bits_0_2),
    .io_tensor_rd_0_data_bits_0_3(tensorAcc_io_tensor_rd_0_data_bits_0_3),
    .io_tensor_rd_0_data_bits_0_4(tensorAcc_io_tensor_rd_0_data_bits_0_4),
    .io_tensor_rd_0_data_bits_0_5(tensorAcc_io_tensor_rd_0_data_bits_0_5),
    .io_tensor_rd_0_data_bits_0_6(tensorAcc_io_tensor_rd_0_data_bits_0_6),
    .io_tensor_rd_0_data_bits_0_7(tensorAcc_io_tensor_rd_0_data_bits_0_7),
    .io_tensor_rd_0_data_bits_0_8(tensorAcc_io_tensor_rd_0_data_bits_0_8),
    .io_tensor_rd_0_data_bits_0_9(tensorAcc_io_tensor_rd_0_data_bits_0_9),
    .io_tensor_rd_0_data_bits_0_10(tensorAcc_io_tensor_rd_0_data_bits_0_10),
    .io_tensor_rd_0_data_bits_0_11(tensorAcc_io_tensor_rd_0_data_bits_0_11),
    .io_tensor_rd_0_data_bits_0_12(tensorAcc_io_tensor_rd_0_data_bits_0_12),
    .io_tensor_rd_0_data_bits_0_13(tensorAcc_io_tensor_rd_0_data_bits_0_13),
    .io_tensor_rd_0_data_bits_0_14(tensorAcc_io_tensor_rd_0_data_bits_0_14),
    .io_tensor_rd_0_data_bits_0_15(tensorAcc_io_tensor_rd_0_data_bits_0_15),
    .io_tensor_rd_0_data_bits_0_16(tensorAcc_io_tensor_rd_0_data_bits_0_16),
    .io_tensor_rd_0_data_bits_0_17(tensorAcc_io_tensor_rd_0_data_bits_0_17),
    .io_tensor_rd_0_data_bits_0_18(tensorAcc_io_tensor_rd_0_data_bits_0_18),
    .io_tensor_rd_0_data_bits_0_19(tensorAcc_io_tensor_rd_0_data_bits_0_19),
    .io_tensor_rd_0_data_bits_0_20(tensorAcc_io_tensor_rd_0_data_bits_0_20),
    .io_tensor_rd_0_data_bits_0_21(tensorAcc_io_tensor_rd_0_data_bits_0_21),
    .io_tensor_rd_0_data_bits_0_22(tensorAcc_io_tensor_rd_0_data_bits_0_22),
    .io_tensor_rd_0_data_bits_0_23(tensorAcc_io_tensor_rd_0_data_bits_0_23),
    .io_tensor_rd_0_data_bits_0_24(tensorAcc_io_tensor_rd_0_data_bits_0_24),
    .io_tensor_rd_0_data_bits_0_25(tensorAcc_io_tensor_rd_0_data_bits_0_25),
    .io_tensor_rd_0_data_bits_0_26(tensorAcc_io_tensor_rd_0_data_bits_0_26),
    .io_tensor_rd_0_data_bits_0_27(tensorAcc_io_tensor_rd_0_data_bits_0_27),
    .io_tensor_rd_0_data_bits_0_28(tensorAcc_io_tensor_rd_0_data_bits_0_28),
    .io_tensor_rd_0_data_bits_0_29(tensorAcc_io_tensor_rd_0_data_bits_0_29),
    .io_tensor_rd_0_data_bits_0_30(tensorAcc_io_tensor_rd_0_data_bits_0_30),
    .io_tensor_rd_0_data_bits_0_31(tensorAcc_io_tensor_rd_0_data_bits_0_31),
    .io_tensor_wr_0_valid(tensorAcc_io_tensor_wr_0_valid),
    .io_tensor_wr_0_bits_idx(tensorAcc_io_tensor_wr_0_bits_idx),
    .io_tensor_wr_0_bits_data_0_0(tensorAcc_io_tensor_wr_0_bits_data_0_0),
    .io_tensor_wr_0_bits_data_0_1(tensorAcc_io_tensor_wr_0_bits_data_0_1),
    .io_tensor_wr_0_bits_data_0_2(tensorAcc_io_tensor_wr_0_bits_data_0_2),
    .io_tensor_wr_0_bits_data_0_3(tensorAcc_io_tensor_wr_0_bits_data_0_3),
    .io_tensor_wr_0_bits_data_0_4(tensorAcc_io_tensor_wr_0_bits_data_0_4),
    .io_tensor_wr_0_bits_data_0_5(tensorAcc_io_tensor_wr_0_bits_data_0_5),
    .io_tensor_wr_0_bits_data_0_6(tensorAcc_io_tensor_wr_0_bits_data_0_6),
    .io_tensor_wr_0_bits_data_0_7(tensorAcc_io_tensor_wr_0_bits_data_0_7),
    .io_tensor_wr_0_bits_data_0_8(tensorAcc_io_tensor_wr_0_bits_data_0_8),
    .io_tensor_wr_0_bits_data_0_9(tensorAcc_io_tensor_wr_0_bits_data_0_9),
    .io_tensor_wr_0_bits_data_0_10(tensorAcc_io_tensor_wr_0_bits_data_0_10),
    .io_tensor_wr_0_bits_data_0_11(tensorAcc_io_tensor_wr_0_bits_data_0_11),
    .io_tensor_wr_0_bits_data_0_12(tensorAcc_io_tensor_wr_0_bits_data_0_12),
    .io_tensor_wr_0_bits_data_0_13(tensorAcc_io_tensor_wr_0_bits_data_0_13),
    .io_tensor_wr_0_bits_data_0_14(tensorAcc_io_tensor_wr_0_bits_data_0_14),
    .io_tensor_wr_0_bits_data_0_15(tensorAcc_io_tensor_wr_0_bits_data_0_15),
    .io_tensor_wr_0_bits_data_0_16(tensorAcc_io_tensor_wr_0_bits_data_0_16),
    .io_tensor_wr_0_bits_data_0_17(tensorAcc_io_tensor_wr_0_bits_data_0_17),
    .io_tensor_wr_0_bits_data_0_18(tensorAcc_io_tensor_wr_0_bits_data_0_18),
    .io_tensor_wr_0_bits_data_0_19(tensorAcc_io_tensor_wr_0_bits_data_0_19),
    .io_tensor_wr_0_bits_data_0_20(tensorAcc_io_tensor_wr_0_bits_data_0_20),
    .io_tensor_wr_0_bits_data_0_21(tensorAcc_io_tensor_wr_0_bits_data_0_21),
    .io_tensor_wr_0_bits_data_0_22(tensorAcc_io_tensor_wr_0_bits_data_0_22),
    .io_tensor_wr_0_bits_data_0_23(tensorAcc_io_tensor_wr_0_bits_data_0_23),
    .io_tensor_wr_0_bits_data_0_24(tensorAcc_io_tensor_wr_0_bits_data_0_24),
    .io_tensor_wr_0_bits_data_0_25(tensorAcc_io_tensor_wr_0_bits_data_0_25),
    .io_tensor_wr_0_bits_data_0_26(tensorAcc_io_tensor_wr_0_bits_data_0_26),
    .io_tensor_wr_0_bits_data_0_27(tensorAcc_io_tensor_wr_0_bits_data_0_27),
    .io_tensor_wr_0_bits_data_0_28(tensorAcc_io_tensor_wr_0_bits_data_0_28),
    .io_tensor_wr_0_bits_data_0_29(tensorAcc_io_tensor_wr_0_bits_data_0_29),
    .io_tensor_wr_0_bits_data_0_30(tensorAcc_io_tensor_wr_0_bits_data_0_30),
    .io_tensor_wr_0_bits_data_0_31(tensorAcc_io_tensor_wr_0_bits_data_0_31)
  );
  TensorGemm tensorGemm ( // @[Compute.scala 63:26]
    .clock(tensorGemm_clock),
    .reset(tensorGemm_reset),
    .io_start(tensorGemm_io_start),
    .io_done(tensorGemm_io_done),
    .io_dec_wgt_1(tensorGemm_io_dec_wgt_1),
    .io_dec_wgt_0(tensorGemm_io_dec_wgt_0),
    .io_dec_inp_1(tensorGemm_io_dec_inp_1),
    .io_dec_inp_0(tensorGemm_io_dec_inp_0),
    .io_dec_acc_1(tensorGemm_io_dec_acc_1),
    .io_dec_acc_0(tensorGemm_io_dec_acc_0),
    .io_dec_empty_0(tensorGemm_io_dec_empty_0),
    .io_dec_lp_1(tensorGemm_io_dec_lp_1),
    .io_dec_lp_0(tensorGemm_io_dec_lp_0),
    .io_dec_uop_end(tensorGemm_io_dec_uop_end),
    .io_dec_uop_begin(tensorGemm_io_dec_uop_begin),
    .io_dec_reset(tensorGemm_io_dec_reset),
    .io_dec_push_next(tensorGemm_io_dec_push_next),
    .io_dec_push_prev(tensorGemm_io_dec_push_prev),
    .io_dec_pop_next(tensorGemm_io_dec_pop_next),
    .io_dec_pop_prev(tensorGemm_io_dec_pop_prev),
    .io_dec_op(tensorGemm_io_dec_op),
    .io_uop_idx_valid(tensorGemm_io_uop_idx_valid),
    .io_uop_idx_bits(tensorGemm_io_uop_idx_bits),
    .io_uop_data_valid(tensorGemm_io_uop_data_valid),
    .io_uop_data_bits_u2(tensorGemm_io_uop_data_bits_u2),
    .io_uop_data_bits_u1(tensorGemm_io_uop_data_bits_u1),
    .io_uop_data_bits_u0(tensorGemm_io_uop_data_bits_u0),
    .io_inp_rd_0_idx_valid(tensorGemm_io_inp_rd_0_idx_valid),
    .io_inp_rd_0_idx_bits(tensorGemm_io_inp_rd_0_idx_bits),
    .io_inp_rd_0_data_valid(tensorGemm_io_inp_rd_0_data_valid),
    .io_inp_rd_0_data_bits_0_0(tensorGemm_io_inp_rd_0_data_bits_0_0),
    .io_inp_rd_0_data_bits_0_1(tensorGemm_io_inp_rd_0_data_bits_0_1),
    .io_inp_rd_0_data_bits_0_2(tensorGemm_io_inp_rd_0_data_bits_0_2),
    .io_inp_rd_0_data_bits_0_3(tensorGemm_io_inp_rd_0_data_bits_0_3),
    .io_inp_rd_0_data_bits_0_4(tensorGemm_io_inp_rd_0_data_bits_0_4),
    .io_inp_rd_0_data_bits_0_5(tensorGemm_io_inp_rd_0_data_bits_0_5),
    .io_inp_rd_0_data_bits_0_6(tensorGemm_io_inp_rd_0_data_bits_0_6),
    .io_inp_rd_0_data_bits_0_7(tensorGemm_io_inp_rd_0_data_bits_0_7),
    .io_inp_rd_0_data_bits_0_8(tensorGemm_io_inp_rd_0_data_bits_0_8),
    .io_inp_rd_0_data_bits_0_9(tensorGemm_io_inp_rd_0_data_bits_0_9),
    .io_inp_rd_0_data_bits_0_10(tensorGemm_io_inp_rd_0_data_bits_0_10),
    .io_inp_rd_0_data_bits_0_11(tensorGemm_io_inp_rd_0_data_bits_0_11),
    .io_inp_rd_0_data_bits_0_12(tensorGemm_io_inp_rd_0_data_bits_0_12),
    .io_inp_rd_0_data_bits_0_13(tensorGemm_io_inp_rd_0_data_bits_0_13),
    .io_inp_rd_0_data_bits_0_14(tensorGemm_io_inp_rd_0_data_bits_0_14),
    .io_inp_rd_0_data_bits_0_15(tensorGemm_io_inp_rd_0_data_bits_0_15),
    .io_wgt_rd_0_idx_valid(tensorGemm_io_wgt_rd_0_idx_valid),
    .io_wgt_rd_0_idx_bits(tensorGemm_io_wgt_rd_0_idx_bits),
    .io_wgt_rd_0_data_valid(tensorGemm_io_wgt_rd_0_data_valid),
    .io_wgt_rd_0_data_bits_0_0(tensorGemm_io_wgt_rd_0_data_bits_0_0),
    .io_wgt_rd_0_data_bits_0_1(tensorGemm_io_wgt_rd_0_data_bits_0_1),
    .io_wgt_rd_0_data_bits_0_2(tensorGemm_io_wgt_rd_0_data_bits_0_2),
    .io_wgt_rd_0_data_bits_0_3(tensorGemm_io_wgt_rd_0_data_bits_0_3),
    .io_wgt_rd_0_data_bits_0_4(tensorGemm_io_wgt_rd_0_data_bits_0_4),
    .io_wgt_rd_0_data_bits_0_5(tensorGemm_io_wgt_rd_0_data_bits_0_5),
    .io_wgt_rd_0_data_bits_0_6(tensorGemm_io_wgt_rd_0_data_bits_0_6),
    .io_wgt_rd_0_data_bits_0_7(tensorGemm_io_wgt_rd_0_data_bits_0_7),
    .io_wgt_rd_0_data_bits_0_8(tensorGemm_io_wgt_rd_0_data_bits_0_8),
    .io_wgt_rd_0_data_bits_0_9(tensorGemm_io_wgt_rd_0_data_bits_0_9),
    .io_wgt_rd_0_data_bits_0_10(tensorGemm_io_wgt_rd_0_data_bits_0_10),
    .io_wgt_rd_0_data_bits_0_11(tensorGemm_io_wgt_rd_0_data_bits_0_11),
    .io_wgt_rd_0_data_bits_0_12(tensorGemm_io_wgt_rd_0_data_bits_0_12),
    .io_wgt_rd_0_data_bits_0_13(tensorGemm_io_wgt_rd_0_data_bits_0_13),
    .io_wgt_rd_0_data_bits_0_14(tensorGemm_io_wgt_rd_0_data_bits_0_14),
    .io_wgt_rd_0_data_bits_0_15(tensorGemm_io_wgt_rd_0_data_bits_0_15),
    .io_wgt_rd_0_data_bits_1_0(tensorGemm_io_wgt_rd_0_data_bits_1_0),
    .io_wgt_rd_0_data_bits_1_1(tensorGemm_io_wgt_rd_0_data_bits_1_1),
    .io_wgt_rd_0_data_bits_1_2(tensorGemm_io_wgt_rd_0_data_bits_1_2),
    .io_wgt_rd_0_data_bits_1_3(tensorGemm_io_wgt_rd_0_data_bits_1_3),
    .io_wgt_rd_0_data_bits_1_4(tensorGemm_io_wgt_rd_0_data_bits_1_4),
    .io_wgt_rd_0_data_bits_1_5(tensorGemm_io_wgt_rd_0_data_bits_1_5),
    .io_wgt_rd_0_data_bits_1_6(tensorGemm_io_wgt_rd_0_data_bits_1_6),
    .io_wgt_rd_0_data_bits_1_7(tensorGemm_io_wgt_rd_0_data_bits_1_7),
    .io_wgt_rd_0_data_bits_1_8(tensorGemm_io_wgt_rd_0_data_bits_1_8),
    .io_wgt_rd_0_data_bits_1_9(tensorGemm_io_wgt_rd_0_data_bits_1_9),
    .io_wgt_rd_0_data_bits_1_10(tensorGemm_io_wgt_rd_0_data_bits_1_10),
    .io_wgt_rd_0_data_bits_1_11(tensorGemm_io_wgt_rd_0_data_bits_1_11),
    .io_wgt_rd_0_data_bits_1_12(tensorGemm_io_wgt_rd_0_data_bits_1_12),
    .io_wgt_rd_0_data_bits_1_13(tensorGemm_io_wgt_rd_0_data_bits_1_13),
    .io_wgt_rd_0_data_bits_1_14(tensorGemm_io_wgt_rd_0_data_bits_1_14),
    .io_wgt_rd_0_data_bits_1_15(tensorGemm_io_wgt_rd_0_data_bits_1_15),
    .io_wgt_rd_0_data_bits_2_0(tensorGemm_io_wgt_rd_0_data_bits_2_0),
    .io_wgt_rd_0_data_bits_2_1(tensorGemm_io_wgt_rd_0_data_bits_2_1),
    .io_wgt_rd_0_data_bits_2_2(tensorGemm_io_wgt_rd_0_data_bits_2_2),
    .io_wgt_rd_0_data_bits_2_3(tensorGemm_io_wgt_rd_0_data_bits_2_3),
    .io_wgt_rd_0_data_bits_2_4(tensorGemm_io_wgt_rd_0_data_bits_2_4),
    .io_wgt_rd_0_data_bits_2_5(tensorGemm_io_wgt_rd_0_data_bits_2_5),
    .io_wgt_rd_0_data_bits_2_6(tensorGemm_io_wgt_rd_0_data_bits_2_6),
    .io_wgt_rd_0_data_bits_2_7(tensorGemm_io_wgt_rd_0_data_bits_2_7),
    .io_wgt_rd_0_data_bits_2_8(tensorGemm_io_wgt_rd_0_data_bits_2_8),
    .io_wgt_rd_0_data_bits_2_9(tensorGemm_io_wgt_rd_0_data_bits_2_9),
    .io_wgt_rd_0_data_bits_2_10(tensorGemm_io_wgt_rd_0_data_bits_2_10),
    .io_wgt_rd_0_data_bits_2_11(tensorGemm_io_wgt_rd_0_data_bits_2_11),
    .io_wgt_rd_0_data_bits_2_12(tensorGemm_io_wgt_rd_0_data_bits_2_12),
    .io_wgt_rd_0_data_bits_2_13(tensorGemm_io_wgt_rd_0_data_bits_2_13),
    .io_wgt_rd_0_data_bits_2_14(tensorGemm_io_wgt_rd_0_data_bits_2_14),
    .io_wgt_rd_0_data_bits_2_15(tensorGemm_io_wgt_rd_0_data_bits_2_15),
    .io_wgt_rd_0_data_bits_3_0(tensorGemm_io_wgt_rd_0_data_bits_3_0),
    .io_wgt_rd_0_data_bits_3_1(tensorGemm_io_wgt_rd_0_data_bits_3_1),
    .io_wgt_rd_0_data_bits_3_2(tensorGemm_io_wgt_rd_0_data_bits_3_2),
    .io_wgt_rd_0_data_bits_3_3(tensorGemm_io_wgt_rd_0_data_bits_3_3),
    .io_wgt_rd_0_data_bits_3_4(tensorGemm_io_wgt_rd_0_data_bits_3_4),
    .io_wgt_rd_0_data_bits_3_5(tensorGemm_io_wgt_rd_0_data_bits_3_5),
    .io_wgt_rd_0_data_bits_3_6(tensorGemm_io_wgt_rd_0_data_bits_3_6),
    .io_wgt_rd_0_data_bits_3_7(tensorGemm_io_wgt_rd_0_data_bits_3_7),
    .io_wgt_rd_0_data_bits_3_8(tensorGemm_io_wgt_rd_0_data_bits_3_8),
    .io_wgt_rd_0_data_bits_3_9(tensorGemm_io_wgt_rd_0_data_bits_3_9),
    .io_wgt_rd_0_data_bits_3_10(tensorGemm_io_wgt_rd_0_data_bits_3_10),
    .io_wgt_rd_0_data_bits_3_11(tensorGemm_io_wgt_rd_0_data_bits_3_11),
    .io_wgt_rd_0_data_bits_3_12(tensorGemm_io_wgt_rd_0_data_bits_3_12),
    .io_wgt_rd_0_data_bits_3_13(tensorGemm_io_wgt_rd_0_data_bits_3_13),
    .io_wgt_rd_0_data_bits_3_14(tensorGemm_io_wgt_rd_0_data_bits_3_14),
    .io_wgt_rd_0_data_bits_3_15(tensorGemm_io_wgt_rd_0_data_bits_3_15),
    .io_wgt_rd_0_data_bits_4_0(tensorGemm_io_wgt_rd_0_data_bits_4_0),
    .io_wgt_rd_0_data_bits_4_1(tensorGemm_io_wgt_rd_0_data_bits_4_1),
    .io_wgt_rd_0_data_bits_4_2(tensorGemm_io_wgt_rd_0_data_bits_4_2),
    .io_wgt_rd_0_data_bits_4_3(tensorGemm_io_wgt_rd_0_data_bits_4_3),
    .io_wgt_rd_0_data_bits_4_4(tensorGemm_io_wgt_rd_0_data_bits_4_4),
    .io_wgt_rd_0_data_bits_4_5(tensorGemm_io_wgt_rd_0_data_bits_4_5),
    .io_wgt_rd_0_data_bits_4_6(tensorGemm_io_wgt_rd_0_data_bits_4_6),
    .io_wgt_rd_0_data_bits_4_7(tensorGemm_io_wgt_rd_0_data_bits_4_7),
    .io_wgt_rd_0_data_bits_4_8(tensorGemm_io_wgt_rd_0_data_bits_4_8),
    .io_wgt_rd_0_data_bits_4_9(tensorGemm_io_wgt_rd_0_data_bits_4_9),
    .io_wgt_rd_0_data_bits_4_10(tensorGemm_io_wgt_rd_0_data_bits_4_10),
    .io_wgt_rd_0_data_bits_4_11(tensorGemm_io_wgt_rd_0_data_bits_4_11),
    .io_wgt_rd_0_data_bits_4_12(tensorGemm_io_wgt_rd_0_data_bits_4_12),
    .io_wgt_rd_0_data_bits_4_13(tensorGemm_io_wgt_rd_0_data_bits_4_13),
    .io_wgt_rd_0_data_bits_4_14(tensorGemm_io_wgt_rd_0_data_bits_4_14),
    .io_wgt_rd_0_data_bits_4_15(tensorGemm_io_wgt_rd_0_data_bits_4_15),
    .io_wgt_rd_0_data_bits_5_0(tensorGemm_io_wgt_rd_0_data_bits_5_0),
    .io_wgt_rd_0_data_bits_5_1(tensorGemm_io_wgt_rd_0_data_bits_5_1),
    .io_wgt_rd_0_data_bits_5_2(tensorGemm_io_wgt_rd_0_data_bits_5_2),
    .io_wgt_rd_0_data_bits_5_3(tensorGemm_io_wgt_rd_0_data_bits_5_3),
    .io_wgt_rd_0_data_bits_5_4(tensorGemm_io_wgt_rd_0_data_bits_5_4),
    .io_wgt_rd_0_data_bits_5_5(tensorGemm_io_wgt_rd_0_data_bits_5_5),
    .io_wgt_rd_0_data_bits_5_6(tensorGemm_io_wgt_rd_0_data_bits_5_6),
    .io_wgt_rd_0_data_bits_5_7(tensorGemm_io_wgt_rd_0_data_bits_5_7),
    .io_wgt_rd_0_data_bits_5_8(tensorGemm_io_wgt_rd_0_data_bits_5_8),
    .io_wgt_rd_0_data_bits_5_9(tensorGemm_io_wgt_rd_0_data_bits_5_9),
    .io_wgt_rd_0_data_bits_5_10(tensorGemm_io_wgt_rd_0_data_bits_5_10),
    .io_wgt_rd_0_data_bits_5_11(tensorGemm_io_wgt_rd_0_data_bits_5_11),
    .io_wgt_rd_0_data_bits_5_12(tensorGemm_io_wgt_rd_0_data_bits_5_12),
    .io_wgt_rd_0_data_bits_5_13(tensorGemm_io_wgt_rd_0_data_bits_5_13),
    .io_wgt_rd_0_data_bits_5_14(tensorGemm_io_wgt_rd_0_data_bits_5_14),
    .io_wgt_rd_0_data_bits_5_15(tensorGemm_io_wgt_rd_0_data_bits_5_15),
    .io_wgt_rd_0_data_bits_6_0(tensorGemm_io_wgt_rd_0_data_bits_6_0),
    .io_wgt_rd_0_data_bits_6_1(tensorGemm_io_wgt_rd_0_data_bits_6_1),
    .io_wgt_rd_0_data_bits_6_2(tensorGemm_io_wgt_rd_0_data_bits_6_2),
    .io_wgt_rd_0_data_bits_6_3(tensorGemm_io_wgt_rd_0_data_bits_6_3),
    .io_wgt_rd_0_data_bits_6_4(tensorGemm_io_wgt_rd_0_data_bits_6_4),
    .io_wgt_rd_0_data_bits_6_5(tensorGemm_io_wgt_rd_0_data_bits_6_5),
    .io_wgt_rd_0_data_bits_6_6(tensorGemm_io_wgt_rd_0_data_bits_6_6),
    .io_wgt_rd_0_data_bits_6_7(tensorGemm_io_wgt_rd_0_data_bits_6_7),
    .io_wgt_rd_0_data_bits_6_8(tensorGemm_io_wgt_rd_0_data_bits_6_8),
    .io_wgt_rd_0_data_bits_6_9(tensorGemm_io_wgt_rd_0_data_bits_6_9),
    .io_wgt_rd_0_data_bits_6_10(tensorGemm_io_wgt_rd_0_data_bits_6_10),
    .io_wgt_rd_0_data_bits_6_11(tensorGemm_io_wgt_rd_0_data_bits_6_11),
    .io_wgt_rd_0_data_bits_6_12(tensorGemm_io_wgt_rd_0_data_bits_6_12),
    .io_wgt_rd_0_data_bits_6_13(tensorGemm_io_wgt_rd_0_data_bits_6_13),
    .io_wgt_rd_0_data_bits_6_14(tensorGemm_io_wgt_rd_0_data_bits_6_14),
    .io_wgt_rd_0_data_bits_6_15(tensorGemm_io_wgt_rd_0_data_bits_6_15),
    .io_wgt_rd_0_data_bits_7_0(tensorGemm_io_wgt_rd_0_data_bits_7_0),
    .io_wgt_rd_0_data_bits_7_1(tensorGemm_io_wgt_rd_0_data_bits_7_1),
    .io_wgt_rd_0_data_bits_7_2(tensorGemm_io_wgt_rd_0_data_bits_7_2),
    .io_wgt_rd_0_data_bits_7_3(tensorGemm_io_wgt_rd_0_data_bits_7_3),
    .io_wgt_rd_0_data_bits_7_4(tensorGemm_io_wgt_rd_0_data_bits_7_4),
    .io_wgt_rd_0_data_bits_7_5(tensorGemm_io_wgt_rd_0_data_bits_7_5),
    .io_wgt_rd_0_data_bits_7_6(tensorGemm_io_wgt_rd_0_data_bits_7_6),
    .io_wgt_rd_0_data_bits_7_7(tensorGemm_io_wgt_rd_0_data_bits_7_7),
    .io_wgt_rd_0_data_bits_7_8(tensorGemm_io_wgt_rd_0_data_bits_7_8),
    .io_wgt_rd_0_data_bits_7_9(tensorGemm_io_wgt_rd_0_data_bits_7_9),
    .io_wgt_rd_0_data_bits_7_10(tensorGemm_io_wgt_rd_0_data_bits_7_10),
    .io_wgt_rd_0_data_bits_7_11(tensorGemm_io_wgt_rd_0_data_bits_7_11),
    .io_wgt_rd_0_data_bits_7_12(tensorGemm_io_wgt_rd_0_data_bits_7_12),
    .io_wgt_rd_0_data_bits_7_13(tensorGemm_io_wgt_rd_0_data_bits_7_13),
    .io_wgt_rd_0_data_bits_7_14(tensorGemm_io_wgt_rd_0_data_bits_7_14),
    .io_wgt_rd_0_data_bits_7_15(tensorGemm_io_wgt_rd_0_data_bits_7_15),
    .io_wgt_rd_0_data_bits_8_0(tensorGemm_io_wgt_rd_0_data_bits_8_0),
    .io_wgt_rd_0_data_bits_8_1(tensorGemm_io_wgt_rd_0_data_bits_8_1),
    .io_wgt_rd_0_data_bits_8_2(tensorGemm_io_wgt_rd_0_data_bits_8_2),
    .io_wgt_rd_0_data_bits_8_3(tensorGemm_io_wgt_rd_0_data_bits_8_3),
    .io_wgt_rd_0_data_bits_8_4(tensorGemm_io_wgt_rd_0_data_bits_8_4),
    .io_wgt_rd_0_data_bits_8_5(tensorGemm_io_wgt_rd_0_data_bits_8_5),
    .io_wgt_rd_0_data_bits_8_6(tensorGemm_io_wgt_rd_0_data_bits_8_6),
    .io_wgt_rd_0_data_bits_8_7(tensorGemm_io_wgt_rd_0_data_bits_8_7),
    .io_wgt_rd_0_data_bits_8_8(tensorGemm_io_wgt_rd_0_data_bits_8_8),
    .io_wgt_rd_0_data_bits_8_9(tensorGemm_io_wgt_rd_0_data_bits_8_9),
    .io_wgt_rd_0_data_bits_8_10(tensorGemm_io_wgt_rd_0_data_bits_8_10),
    .io_wgt_rd_0_data_bits_8_11(tensorGemm_io_wgt_rd_0_data_bits_8_11),
    .io_wgt_rd_0_data_bits_8_12(tensorGemm_io_wgt_rd_0_data_bits_8_12),
    .io_wgt_rd_0_data_bits_8_13(tensorGemm_io_wgt_rd_0_data_bits_8_13),
    .io_wgt_rd_0_data_bits_8_14(tensorGemm_io_wgt_rd_0_data_bits_8_14),
    .io_wgt_rd_0_data_bits_8_15(tensorGemm_io_wgt_rd_0_data_bits_8_15),
    .io_wgt_rd_0_data_bits_9_0(tensorGemm_io_wgt_rd_0_data_bits_9_0),
    .io_wgt_rd_0_data_bits_9_1(tensorGemm_io_wgt_rd_0_data_bits_9_1),
    .io_wgt_rd_0_data_bits_9_2(tensorGemm_io_wgt_rd_0_data_bits_9_2),
    .io_wgt_rd_0_data_bits_9_3(tensorGemm_io_wgt_rd_0_data_bits_9_3),
    .io_wgt_rd_0_data_bits_9_4(tensorGemm_io_wgt_rd_0_data_bits_9_4),
    .io_wgt_rd_0_data_bits_9_5(tensorGemm_io_wgt_rd_0_data_bits_9_5),
    .io_wgt_rd_0_data_bits_9_6(tensorGemm_io_wgt_rd_0_data_bits_9_6),
    .io_wgt_rd_0_data_bits_9_7(tensorGemm_io_wgt_rd_0_data_bits_9_7),
    .io_wgt_rd_0_data_bits_9_8(tensorGemm_io_wgt_rd_0_data_bits_9_8),
    .io_wgt_rd_0_data_bits_9_9(tensorGemm_io_wgt_rd_0_data_bits_9_9),
    .io_wgt_rd_0_data_bits_9_10(tensorGemm_io_wgt_rd_0_data_bits_9_10),
    .io_wgt_rd_0_data_bits_9_11(tensorGemm_io_wgt_rd_0_data_bits_9_11),
    .io_wgt_rd_0_data_bits_9_12(tensorGemm_io_wgt_rd_0_data_bits_9_12),
    .io_wgt_rd_0_data_bits_9_13(tensorGemm_io_wgt_rd_0_data_bits_9_13),
    .io_wgt_rd_0_data_bits_9_14(tensorGemm_io_wgt_rd_0_data_bits_9_14),
    .io_wgt_rd_0_data_bits_9_15(tensorGemm_io_wgt_rd_0_data_bits_9_15),
    .io_wgt_rd_0_data_bits_10_0(tensorGemm_io_wgt_rd_0_data_bits_10_0),
    .io_wgt_rd_0_data_bits_10_1(tensorGemm_io_wgt_rd_0_data_bits_10_1),
    .io_wgt_rd_0_data_bits_10_2(tensorGemm_io_wgt_rd_0_data_bits_10_2),
    .io_wgt_rd_0_data_bits_10_3(tensorGemm_io_wgt_rd_0_data_bits_10_3),
    .io_wgt_rd_0_data_bits_10_4(tensorGemm_io_wgt_rd_0_data_bits_10_4),
    .io_wgt_rd_0_data_bits_10_5(tensorGemm_io_wgt_rd_0_data_bits_10_5),
    .io_wgt_rd_0_data_bits_10_6(tensorGemm_io_wgt_rd_0_data_bits_10_6),
    .io_wgt_rd_0_data_bits_10_7(tensorGemm_io_wgt_rd_0_data_bits_10_7),
    .io_wgt_rd_0_data_bits_10_8(tensorGemm_io_wgt_rd_0_data_bits_10_8),
    .io_wgt_rd_0_data_bits_10_9(tensorGemm_io_wgt_rd_0_data_bits_10_9),
    .io_wgt_rd_0_data_bits_10_10(tensorGemm_io_wgt_rd_0_data_bits_10_10),
    .io_wgt_rd_0_data_bits_10_11(tensorGemm_io_wgt_rd_0_data_bits_10_11),
    .io_wgt_rd_0_data_bits_10_12(tensorGemm_io_wgt_rd_0_data_bits_10_12),
    .io_wgt_rd_0_data_bits_10_13(tensorGemm_io_wgt_rd_0_data_bits_10_13),
    .io_wgt_rd_0_data_bits_10_14(tensorGemm_io_wgt_rd_0_data_bits_10_14),
    .io_wgt_rd_0_data_bits_10_15(tensorGemm_io_wgt_rd_0_data_bits_10_15),
    .io_wgt_rd_0_data_bits_11_0(tensorGemm_io_wgt_rd_0_data_bits_11_0),
    .io_wgt_rd_0_data_bits_11_1(tensorGemm_io_wgt_rd_0_data_bits_11_1),
    .io_wgt_rd_0_data_bits_11_2(tensorGemm_io_wgt_rd_0_data_bits_11_2),
    .io_wgt_rd_0_data_bits_11_3(tensorGemm_io_wgt_rd_0_data_bits_11_3),
    .io_wgt_rd_0_data_bits_11_4(tensorGemm_io_wgt_rd_0_data_bits_11_4),
    .io_wgt_rd_0_data_bits_11_5(tensorGemm_io_wgt_rd_0_data_bits_11_5),
    .io_wgt_rd_0_data_bits_11_6(tensorGemm_io_wgt_rd_0_data_bits_11_6),
    .io_wgt_rd_0_data_bits_11_7(tensorGemm_io_wgt_rd_0_data_bits_11_7),
    .io_wgt_rd_0_data_bits_11_8(tensorGemm_io_wgt_rd_0_data_bits_11_8),
    .io_wgt_rd_0_data_bits_11_9(tensorGemm_io_wgt_rd_0_data_bits_11_9),
    .io_wgt_rd_0_data_bits_11_10(tensorGemm_io_wgt_rd_0_data_bits_11_10),
    .io_wgt_rd_0_data_bits_11_11(tensorGemm_io_wgt_rd_0_data_bits_11_11),
    .io_wgt_rd_0_data_bits_11_12(tensorGemm_io_wgt_rd_0_data_bits_11_12),
    .io_wgt_rd_0_data_bits_11_13(tensorGemm_io_wgt_rd_0_data_bits_11_13),
    .io_wgt_rd_0_data_bits_11_14(tensorGemm_io_wgt_rd_0_data_bits_11_14),
    .io_wgt_rd_0_data_bits_11_15(tensorGemm_io_wgt_rd_0_data_bits_11_15),
    .io_wgt_rd_0_data_bits_12_0(tensorGemm_io_wgt_rd_0_data_bits_12_0),
    .io_wgt_rd_0_data_bits_12_1(tensorGemm_io_wgt_rd_0_data_bits_12_1),
    .io_wgt_rd_0_data_bits_12_2(tensorGemm_io_wgt_rd_0_data_bits_12_2),
    .io_wgt_rd_0_data_bits_12_3(tensorGemm_io_wgt_rd_0_data_bits_12_3),
    .io_wgt_rd_0_data_bits_12_4(tensorGemm_io_wgt_rd_0_data_bits_12_4),
    .io_wgt_rd_0_data_bits_12_5(tensorGemm_io_wgt_rd_0_data_bits_12_5),
    .io_wgt_rd_0_data_bits_12_6(tensorGemm_io_wgt_rd_0_data_bits_12_6),
    .io_wgt_rd_0_data_bits_12_7(tensorGemm_io_wgt_rd_0_data_bits_12_7),
    .io_wgt_rd_0_data_bits_12_8(tensorGemm_io_wgt_rd_0_data_bits_12_8),
    .io_wgt_rd_0_data_bits_12_9(tensorGemm_io_wgt_rd_0_data_bits_12_9),
    .io_wgt_rd_0_data_bits_12_10(tensorGemm_io_wgt_rd_0_data_bits_12_10),
    .io_wgt_rd_0_data_bits_12_11(tensorGemm_io_wgt_rd_0_data_bits_12_11),
    .io_wgt_rd_0_data_bits_12_12(tensorGemm_io_wgt_rd_0_data_bits_12_12),
    .io_wgt_rd_0_data_bits_12_13(tensorGemm_io_wgt_rd_0_data_bits_12_13),
    .io_wgt_rd_0_data_bits_12_14(tensorGemm_io_wgt_rd_0_data_bits_12_14),
    .io_wgt_rd_0_data_bits_12_15(tensorGemm_io_wgt_rd_0_data_bits_12_15),
    .io_wgt_rd_0_data_bits_13_0(tensorGemm_io_wgt_rd_0_data_bits_13_0),
    .io_wgt_rd_0_data_bits_13_1(tensorGemm_io_wgt_rd_0_data_bits_13_1),
    .io_wgt_rd_0_data_bits_13_2(tensorGemm_io_wgt_rd_0_data_bits_13_2),
    .io_wgt_rd_0_data_bits_13_3(tensorGemm_io_wgt_rd_0_data_bits_13_3),
    .io_wgt_rd_0_data_bits_13_4(tensorGemm_io_wgt_rd_0_data_bits_13_4),
    .io_wgt_rd_0_data_bits_13_5(tensorGemm_io_wgt_rd_0_data_bits_13_5),
    .io_wgt_rd_0_data_bits_13_6(tensorGemm_io_wgt_rd_0_data_bits_13_6),
    .io_wgt_rd_0_data_bits_13_7(tensorGemm_io_wgt_rd_0_data_bits_13_7),
    .io_wgt_rd_0_data_bits_13_8(tensorGemm_io_wgt_rd_0_data_bits_13_8),
    .io_wgt_rd_0_data_bits_13_9(tensorGemm_io_wgt_rd_0_data_bits_13_9),
    .io_wgt_rd_0_data_bits_13_10(tensorGemm_io_wgt_rd_0_data_bits_13_10),
    .io_wgt_rd_0_data_bits_13_11(tensorGemm_io_wgt_rd_0_data_bits_13_11),
    .io_wgt_rd_0_data_bits_13_12(tensorGemm_io_wgt_rd_0_data_bits_13_12),
    .io_wgt_rd_0_data_bits_13_13(tensorGemm_io_wgt_rd_0_data_bits_13_13),
    .io_wgt_rd_0_data_bits_13_14(tensorGemm_io_wgt_rd_0_data_bits_13_14),
    .io_wgt_rd_0_data_bits_13_15(tensorGemm_io_wgt_rd_0_data_bits_13_15),
    .io_wgt_rd_0_data_bits_14_0(tensorGemm_io_wgt_rd_0_data_bits_14_0),
    .io_wgt_rd_0_data_bits_14_1(tensorGemm_io_wgt_rd_0_data_bits_14_1),
    .io_wgt_rd_0_data_bits_14_2(tensorGemm_io_wgt_rd_0_data_bits_14_2),
    .io_wgt_rd_0_data_bits_14_3(tensorGemm_io_wgt_rd_0_data_bits_14_3),
    .io_wgt_rd_0_data_bits_14_4(tensorGemm_io_wgt_rd_0_data_bits_14_4),
    .io_wgt_rd_0_data_bits_14_5(tensorGemm_io_wgt_rd_0_data_bits_14_5),
    .io_wgt_rd_0_data_bits_14_6(tensorGemm_io_wgt_rd_0_data_bits_14_6),
    .io_wgt_rd_0_data_bits_14_7(tensorGemm_io_wgt_rd_0_data_bits_14_7),
    .io_wgt_rd_0_data_bits_14_8(tensorGemm_io_wgt_rd_0_data_bits_14_8),
    .io_wgt_rd_0_data_bits_14_9(tensorGemm_io_wgt_rd_0_data_bits_14_9),
    .io_wgt_rd_0_data_bits_14_10(tensorGemm_io_wgt_rd_0_data_bits_14_10),
    .io_wgt_rd_0_data_bits_14_11(tensorGemm_io_wgt_rd_0_data_bits_14_11),
    .io_wgt_rd_0_data_bits_14_12(tensorGemm_io_wgt_rd_0_data_bits_14_12),
    .io_wgt_rd_0_data_bits_14_13(tensorGemm_io_wgt_rd_0_data_bits_14_13),
    .io_wgt_rd_0_data_bits_14_14(tensorGemm_io_wgt_rd_0_data_bits_14_14),
    .io_wgt_rd_0_data_bits_14_15(tensorGemm_io_wgt_rd_0_data_bits_14_15),
    .io_wgt_rd_0_data_bits_15_0(tensorGemm_io_wgt_rd_0_data_bits_15_0),
    .io_wgt_rd_0_data_bits_15_1(tensorGemm_io_wgt_rd_0_data_bits_15_1),
    .io_wgt_rd_0_data_bits_15_2(tensorGemm_io_wgt_rd_0_data_bits_15_2),
    .io_wgt_rd_0_data_bits_15_3(tensorGemm_io_wgt_rd_0_data_bits_15_3),
    .io_wgt_rd_0_data_bits_15_4(tensorGemm_io_wgt_rd_0_data_bits_15_4),
    .io_wgt_rd_0_data_bits_15_5(tensorGemm_io_wgt_rd_0_data_bits_15_5),
    .io_wgt_rd_0_data_bits_15_6(tensorGemm_io_wgt_rd_0_data_bits_15_6),
    .io_wgt_rd_0_data_bits_15_7(tensorGemm_io_wgt_rd_0_data_bits_15_7),
    .io_wgt_rd_0_data_bits_15_8(tensorGemm_io_wgt_rd_0_data_bits_15_8),
    .io_wgt_rd_0_data_bits_15_9(tensorGemm_io_wgt_rd_0_data_bits_15_9),
    .io_wgt_rd_0_data_bits_15_10(tensorGemm_io_wgt_rd_0_data_bits_15_10),
    .io_wgt_rd_0_data_bits_15_11(tensorGemm_io_wgt_rd_0_data_bits_15_11),
    .io_wgt_rd_0_data_bits_15_12(tensorGemm_io_wgt_rd_0_data_bits_15_12),
    .io_wgt_rd_0_data_bits_15_13(tensorGemm_io_wgt_rd_0_data_bits_15_13),
    .io_wgt_rd_0_data_bits_15_14(tensorGemm_io_wgt_rd_0_data_bits_15_14),
    .io_wgt_rd_0_data_bits_15_15(tensorGemm_io_wgt_rd_0_data_bits_15_15),
    .io_wgt_rd_0_data_bits_16_0(tensorGemm_io_wgt_rd_0_data_bits_16_0),
    .io_wgt_rd_0_data_bits_16_1(tensorGemm_io_wgt_rd_0_data_bits_16_1),
    .io_wgt_rd_0_data_bits_16_2(tensorGemm_io_wgt_rd_0_data_bits_16_2),
    .io_wgt_rd_0_data_bits_16_3(tensorGemm_io_wgt_rd_0_data_bits_16_3),
    .io_wgt_rd_0_data_bits_16_4(tensorGemm_io_wgt_rd_0_data_bits_16_4),
    .io_wgt_rd_0_data_bits_16_5(tensorGemm_io_wgt_rd_0_data_bits_16_5),
    .io_wgt_rd_0_data_bits_16_6(tensorGemm_io_wgt_rd_0_data_bits_16_6),
    .io_wgt_rd_0_data_bits_16_7(tensorGemm_io_wgt_rd_0_data_bits_16_7),
    .io_wgt_rd_0_data_bits_16_8(tensorGemm_io_wgt_rd_0_data_bits_16_8),
    .io_wgt_rd_0_data_bits_16_9(tensorGemm_io_wgt_rd_0_data_bits_16_9),
    .io_wgt_rd_0_data_bits_16_10(tensorGemm_io_wgt_rd_0_data_bits_16_10),
    .io_wgt_rd_0_data_bits_16_11(tensorGemm_io_wgt_rd_0_data_bits_16_11),
    .io_wgt_rd_0_data_bits_16_12(tensorGemm_io_wgt_rd_0_data_bits_16_12),
    .io_wgt_rd_0_data_bits_16_13(tensorGemm_io_wgt_rd_0_data_bits_16_13),
    .io_wgt_rd_0_data_bits_16_14(tensorGemm_io_wgt_rd_0_data_bits_16_14),
    .io_wgt_rd_0_data_bits_16_15(tensorGemm_io_wgt_rd_0_data_bits_16_15),
    .io_wgt_rd_0_data_bits_17_0(tensorGemm_io_wgt_rd_0_data_bits_17_0),
    .io_wgt_rd_0_data_bits_17_1(tensorGemm_io_wgt_rd_0_data_bits_17_1),
    .io_wgt_rd_0_data_bits_17_2(tensorGemm_io_wgt_rd_0_data_bits_17_2),
    .io_wgt_rd_0_data_bits_17_3(tensorGemm_io_wgt_rd_0_data_bits_17_3),
    .io_wgt_rd_0_data_bits_17_4(tensorGemm_io_wgt_rd_0_data_bits_17_4),
    .io_wgt_rd_0_data_bits_17_5(tensorGemm_io_wgt_rd_0_data_bits_17_5),
    .io_wgt_rd_0_data_bits_17_6(tensorGemm_io_wgt_rd_0_data_bits_17_6),
    .io_wgt_rd_0_data_bits_17_7(tensorGemm_io_wgt_rd_0_data_bits_17_7),
    .io_wgt_rd_0_data_bits_17_8(tensorGemm_io_wgt_rd_0_data_bits_17_8),
    .io_wgt_rd_0_data_bits_17_9(tensorGemm_io_wgt_rd_0_data_bits_17_9),
    .io_wgt_rd_0_data_bits_17_10(tensorGemm_io_wgt_rd_0_data_bits_17_10),
    .io_wgt_rd_0_data_bits_17_11(tensorGemm_io_wgt_rd_0_data_bits_17_11),
    .io_wgt_rd_0_data_bits_17_12(tensorGemm_io_wgt_rd_0_data_bits_17_12),
    .io_wgt_rd_0_data_bits_17_13(tensorGemm_io_wgt_rd_0_data_bits_17_13),
    .io_wgt_rd_0_data_bits_17_14(tensorGemm_io_wgt_rd_0_data_bits_17_14),
    .io_wgt_rd_0_data_bits_17_15(tensorGemm_io_wgt_rd_0_data_bits_17_15),
    .io_wgt_rd_0_data_bits_18_0(tensorGemm_io_wgt_rd_0_data_bits_18_0),
    .io_wgt_rd_0_data_bits_18_1(tensorGemm_io_wgt_rd_0_data_bits_18_1),
    .io_wgt_rd_0_data_bits_18_2(tensorGemm_io_wgt_rd_0_data_bits_18_2),
    .io_wgt_rd_0_data_bits_18_3(tensorGemm_io_wgt_rd_0_data_bits_18_3),
    .io_wgt_rd_0_data_bits_18_4(tensorGemm_io_wgt_rd_0_data_bits_18_4),
    .io_wgt_rd_0_data_bits_18_5(tensorGemm_io_wgt_rd_0_data_bits_18_5),
    .io_wgt_rd_0_data_bits_18_6(tensorGemm_io_wgt_rd_0_data_bits_18_6),
    .io_wgt_rd_0_data_bits_18_7(tensorGemm_io_wgt_rd_0_data_bits_18_7),
    .io_wgt_rd_0_data_bits_18_8(tensorGemm_io_wgt_rd_0_data_bits_18_8),
    .io_wgt_rd_0_data_bits_18_9(tensorGemm_io_wgt_rd_0_data_bits_18_9),
    .io_wgt_rd_0_data_bits_18_10(tensorGemm_io_wgt_rd_0_data_bits_18_10),
    .io_wgt_rd_0_data_bits_18_11(tensorGemm_io_wgt_rd_0_data_bits_18_11),
    .io_wgt_rd_0_data_bits_18_12(tensorGemm_io_wgt_rd_0_data_bits_18_12),
    .io_wgt_rd_0_data_bits_18_13(tensorGemm_io_wgt_rd_0_data_bits_18_13),
    .io_wgt_rd_0_data_bits_18_14(tensorGemm_io_wgt_rd_0_data_bits_18_14),
    .io_wgt_rd_0_data_bits_18_15(tensorGemm_io_wgt_rd_0_data_bits_18_15),
    .io_wgt_rd_0_data_bits_19_0(tensorGemm_io_wgt_rd_0_data_bits_19_0),
    .io_wgt_rd_0_data_bits_19_1(tensorGemm_io_wgt_rd_0_data_bits_19_1),
    .io_wgt_rd_0_data_bits_19_2(tensorGemm_io_wgt_rd_0_data_bits_19_2),
    .io_wgt_rd_0_data_bits_19_3(tensorGemm_io_wgt_rd_0_data_bits_19_3),
    .io_wgt_rd_0_data_bits_19_4(tensorGemm_io_wgt_rd_0_data_bits_19_4),
    .io_wgt_rd_0_data_bits_19_5(tensorGemm_io_wgt_rd_0_data_bits_19_5),
    .io_wgt_rd_0_data_bits_19_6(tensorGemm_io_wgt_rd_0_data_bits_19_6),
    .io_wgt_rd_0_data_bits_19_7(tensorGemm_io_wgt_rd_0_data_bits_19_7),
    .io_wgt_rd_0_data_bits_19_8(tensorGemm_io_wgt_rd_0_data_bits_19_8),
    .io_wgt_rd_0_data_bits_19_9(tensorGemm_io_wgt_rd_0_data_bits_19_9),
    .io_wgt_rd_0_data_bits_19_10(tensorGemm_io_wgt_rd_0_data_bits_19_10),
    .io_wgt_rd_0_data_bits_19_11(tensorGemm_io_wgt_rd_0_data_bits_19_11),
    .io_wgt_rd_0_data_bits_19_12(tensorGemm_io_wgt_rd_0_data_bits_19_12),
    .io_wgt_rd_0_data_bits_19_13(tensorGemm_io_wgt_rd_0_data_bits_19_13),
    .io_wgt_rd_0_data_bits_19_14(tensorGemm_io_wgt_rd_0_data_bits_19_14),
    .io_wgt_rd_0_data_bits_19_15(tensorGemm_io_wgt_rd_0_data_bits_19_15),
    .io_wgt_rd_0_data_bits_20_0(tensorGemm_io_wgt_rd_0_data_bits_20_0),
    .io_wgt_rd_0_data_bits_20_1(tensorGemm_io_wgt_rd_0_data_bits_20_1),
    .io_wgt_rd_0_data_bits_20_2(tensorGemm_io_wgt_rd_0_data_bits_20_2),
    .io_wgt_rd_0_data_bits_20_3(tensorGemm_io_wgt_rd_0_data_bits_20_3),
    .io_wgt_rd_0_data_bits_20_4(tensorGemm_io_wgt_rd_0_data_bits_20_4),
    .io_wgt_rd_0_data_bits_20_5(tensorGemm_io_wgt_rd_0_data_bits_20_5),
    .io_wgt_rd_0_data_bits_20_6(tensorGemm_io_wgt_rd_0_data_bits_20_6),
    .io_wgt_rd_0_data_bits_20_7(tensorGemm_io_wgt_rd_0_data_bits_20_7),
    .io_wgt_rd_0_data_bits_20_8(tensorGemm_io_wgt_rd_0_data_bits_20_8),
    .io_wgt_rd_0_data_bits_20_9(tensorGemm_io_wgt_rd_0_data_bits_20_9),
    .io_wgt_rd_0_data_bits_20_10(tensorGemm_io_wgt_rd_0_data_bits_20_10),
    .io_wgt_rd_0_data_bits_20_11(tensorGemm_io_wgt_rd_0_data_bits_20_11),
    .io_wgt_rd_0_data_bits_20_12(tensorGemm_io_wgt_rd_0_data_bits_20_12),
    .io_wgt_rd_0_data_bits_20_13(tensorGemm_io_wgt_rd_0_data_bits_20_13),
    .io_wgt_rd_0_data_bits_20_14(tensorGemm_io_wgt_rd_0_data_bits_20_14),
    .io_wgt_rd_0_data_bits_20_15(tensorGemm_io_wgt_rd_0_data_bits_20_15),
    .io_wgt_rd_0_data_bits_21_0(tensorGemm_io_wgt_rd_0_data_bits_21_0),
    .io_wgt_rd_0_data_bits_21_1(tensorGemm_io_wgt_rd_0_data_bits_21_1),
    .io_wgt_rd_0_data_bits_21_2(tensorGemm_io_wgt_rd_0_data_bits_21_2),
    .io_wgt_rd_0_data_bits_21_3(tensorGemm_io_wgt_rd_0_data_bits_21_3),
    .io_wgt_rd_0_data_bits_21_4(tensorGemm_io_wgt_rd_0_data_bits_21_4),
    .io_wgt_rd_0_data_bits_21_5(tensorGemm_io_wgt_rd_0_data_bits_21_5),
    .io_wgt_rd_0_data_bits_21_6(tensorGemm_io_wgt_rd_0_data_bits_21_6),
    .io_wgt_rd_0_data_bits_21_7(tensorGemm_io_wgt_rd_0_data_bits_21_7),
    .io_wgt_rd_0_data_bits_21_8(tensorGemm_io_wgt_rd_0_data_bits_21_8),
    .io_wgt_rd_0_data_bits_21_9(tensorGemm_io_wgt_rd_0_data_bits_21_9),
    .io_wgt_rd_0_data_bits_21_10(tensorGemm_io_wgt_rd_0_data_bits_21_10),
    .io_wgt_rd_0_data_bits_21_11(tensorGemm_io_wgt_rd_0_data_bits_21_11),
    .io_wgt_rd_0_data_bits_21_12(tensorGemm_io_wgt_rd_0_data_bits_21_12),
    .io_wgt_rd_0_data_bits_21_13(tensorGemm_io_wgt_rd_0_data_bits_21_13),
    .io_wgt_rd_0_data_bits_21_14(tensorGemm_io_wgt_rd_0_data_bits_21_14),
    .io_wgt_rd_0_data_bits_21_15(tensorGemm_io_wgt_rd_0_data_bits_21_15),
    .io_wgt_rd_0_data_bits_22_0(tensorGemm_io_wgt_rd_0_data_bits_22_0),
    .io_wgt_rd_0_data_bits_22_1(tensorGemm_io_wgt_rd_0_data_bits_22_1),
    .io_wgt_rd_0_data_bits_22_2(tensorGemm_io_wgt_rd_0_data_bits_22_2),
    .io_wgt_rd_0_data_bits_22_3(tensorGemm_io_wgt_rd_0_data_bits_22_3),
    .io_wgt_rd_0_data_bits_22_4(tensorGemm_io_wgt_rd_0_data_bits_22_4),
    .io_wgt_rd_0_data_bits_22_5(tensorGemm_io_wgt_rd_0_data_bits_22_5),
    .io_wgt_rd_0_data_bits_22_6(tensorGemm_io_wgt_rd_0_data_bits_22_6),
    .io_wgt_rd_0_data_bits_22_7(tensorGemm_io_wgt_rd_0_data_bits_22_7),
    .io_wgt_rd_0_data_bits_22_8(tensorGemm_io_wgt_rd_0_data_bits_22_8),
    .io_wgt_rd_0_data_bits_22_9(tensorGemm_io_wgt_rd_0_data_bits_22_9),
    .io_wgt_rd_0_data_bits_22_10(tensorGemm_io_wgt_rd_0_data_bits_22_10),
    .io_wgt_rd_0_data_bits_22_11(tensorGemm_io_wgt_rd_0_data_bits_22_11),
    .io_wgt_rd_0_data_bits_22_12(tensorGemm_io_wgt_rd_0_data_bits_22_12),
    .io_wgt_rd_0_data_bits_22_13(tensorGemm_io_wgt_rd_0_data_bits_22_13),
    .io_wgt_rd_0_data_bits_22_14(tensorGemm_io_wgt_rd_0_data_bits_22_14),
    .io_wgt_rd_0_data_bits_22_15(tensorGemm_io_wgt_rd_0_data_bits_22_15),
    .io_wgt_rd_0_data_bits_23_0(tensorGemm_io_wgt_rd_0_data_bits_23_0),
    .io_wgt_rd_0_data_bits_23_1(tensorGemm_io_wgt_rd_0_data_bits_23_1),
    .io_wgt_rd_0_data_bits_23_2(tensorGemm_io_wgt_rd_0_data_bits_23_2),
    .io_wgt_rd_0_data_bits_23_3(tensorGemm_io_wgt_rd_0_data_bits_23_3),
    .io_wgt_rd_0_data_bits_23_4(tensorGemm_io_wgt_rd_0_data_bits_23_4),
    .io_wgt_rd_0_data_bits_23_5(tensorGemm_io_wgt_rd_0_data_bits_23_5),
    .io_wgt_rd_0_data_bits_23_6(tensorGemm_io_wgt_rd_0_data_bits_23_6),
    .io_wgt_rd_0_data_bits_23_7(tensorGemm_io_wgt_rd_0_data_bits_23_7),
    .io_wgt_rd_0_data_bits_23_8(tensorGemm_io_wgt_rd_0_data_bits_23_8),
    .io_wgt_rd_0_data_bits_23_9(tensorGemm_io_wgt_rd_0_data_bits_23_9),
    .io_wgt_rd_0_data_bits_23_10(tensorGemm_io_wgt_rd_0_data_bits_23_10),
    .io_wgt_rd_0_data_bits_23_11(tensorGemm_io_wgt_rd_0_data_bits_23_11),
    .io_wgt_rd_0_data_bits_23_12(tensorGemm_io_wgt_rd_0_data_bits_23_12),
    .io_wgt_rd_0_data_bits_23_13(tensorGemm_io_wgt_rd_0_data_bits_23_13),
    .io_wgt_rd_0_data_bits_23_14(tensorGemm_io_wgt_rd_0_data_bits_23_14),
    .io_wgt_rd_0_data_bits_23_15(tensorGemm_io_wgt_rd_0_data_bits_23_15),
    .io_wgt_rd_0_data_bits_24_0(tensorGemm_io_wgt_rd_0_data_bits_24_0),
    .io_wgt_rd_0_data_bits_24_1(tensorGemm_io_wgt_rd_0_data_bits_24_1),
    .io_wgt_rd_0_data_bits_24_2(tensorGemm_io_wgt_rd_0_data_bits_24_2),
    .io_wgt_rd_0_data_bits_24_3(tensorGemm_io_wgt_rd_0_data_bits_24_3),
    .io_wgt_rd_0_data_bits_24_4(tensorGemm_io_wgt_rd_0_data_bits_24_4),
    .io_wgt_rd_0_data_bits_24_5(tensorGemm_io_wgt_rd_0_data_bits_24_5),
    .io_wgt_rd_0_data_bits_24_6(tensorGemm_io_wgt_rd_0_data_bits_24_6),
    .io_wgt_rd_0_data_bits_24_7(tensorGemm_io_wgt_rd_0_data_bits_24_7),
    .io_wgt_rd_0_data_bits_24_8(tensorGemm_io_wgt_rd_0_data_bits_24_8),
    .io_wgt_rd_0_data_bits_24_9(tensorGemm_io_wgt_rd_0_data_bits_24_9),
    .io_wgt_rd_0_data_bits_24_10(tensorGemm_io_wgt_rd_0_data_bits_24_10),
    .io_wgt_rd_0_data_bits_24_11(tensorGemm_io_wgt_rd_0_data_bits_24_11),
    .io_wgt_rd_0_data_bits_24_12(tensorGemm_io_wgt_rd_0_data_bits_24_12),
    .io_wgt_rd_0_data_bits_24_13(tensorGemm_io_wgt_rd_0_data_bits_24_13),
    .io_wgt_rd_0_data_bits_24_14(tensorGemm_io_wgt_rd_0_data_bits_24_14),
    .io_wgt_rd_0_data_bits_24_15(tensorGemm_io_wgt_rd_0_data_bits_24_15),
    .io_wgt_rd_0_data_bits_25_0(tensorGemm_io_wgt_rd_0_data_bits_25_0),
    .io_wgt_rd_0_data_bits_25_1(tensorGemm_io_wgt_rd_0_data_bits_25_1),
    .io_wgt_rd_0_data_bits_25_2(tensorGemm_io_wgt_rd_0_data_bits_25_2),
    .io_wgt_rd_0_data_bits_25_3(tensorGemm_io_wgt_rd_0_data_bits_25_3),
    .io_wgt_rd_0_data_bits_25_4(tensorGemm_io_wgt_rd_0_data_bits_25_4),
    .io_wgt_rd_0_data_bits_25_5(tensorGemm_io_wgt_rd_0_data_bits_25_5),
    .io_wgt_rd_0_data_bits_25_6(tensorGemm_io_wgt_rd_0_data_bits_25_6),
    .io_wgt_rd_0_data_bits_25_7(tensorGemm_io_wgt_rd_0_data_bits_25_7),
    .io_wgt_rd_0_data_bits_25_8(tensorGemm_io_wgt_rd_0_data_bits_25_8),
    .io_wgt_rd_0_data_bits_25_9(tensorGemm_io_wgt_rd_0_data_bits_25_9),
    .io_wgt_rd_0_data_bits_25_10(tensorGemm_io_wgt_rd_0_data_bits_25_10),
    .io_wgt_rd_0_data_bits_25_11(tensorGemm_io_wgt_rd_0_data_bits_25_11),
    .io_wgt_rd_0_data_bits_25_12(tensorGemm_io_wgt_rd_0_data_bits_25_12),
    .io_wgt_rd_0_data_bits_25_13(tensorGemm_io_wgt_rd_0_data_bits_25_13),
    .io_wgt_rd_0_data_bits_25_14(tensorGemm_io_wgt_rd_0_data_bits_25_14),
    .io_wgt_rd_0_data_bits_25_15(tensorGemm_io_wgt_rd_0_data_bits_25_15),
    .io_wgt_rd_0_data_bits_26_0(tensorGemm_io_wgt_rd_0_data_bits_26_0),
    .io_wgt_rd_0_data_bits_26_1(tensorGemm_io_wgt_rd_0_data_bits_26_1),
    .io_wgt_rd_0_data_bits_26_2(tensorGemm_io_wgt_rd_0_data_bits_26_2),
    .io_wgt_rd_0_data_bits_26_3(tensorGemm_io_wgt_rd_0_data_bits_26_3),
    .io_wgt_rd_0_data_bits_26_4(tensorGemm_io_wgt_rd_0_data_bits_26_4),
    .io_wgt_rd_0_data_bits_26_5(tensorGemm_io_wgt_rd_0_data_bits_26_5),
    .io_wgt_rd_0_data_bits_26_6(tensorGemm_io_wgt_rd_0_data_bits_26_6),
    .io_wgt_rd_0_data_bits_26_7(tensorGemm_io_wgt_rd_0_data_bits_26_7),
    .io_wgt_rd_0_data_bits_26_8(tensorGemm_io_wgt_rd_0_data_bits_26_8),
    .io_wgt_rd_0_data_bits_26_9(tensorGemm_io_wgt_rd_0_data_bits_26_9),
    .io_wgt_rd_0_data_bits_26_10(tensorGemm_io_wgt_rd_0_data_bits_26_10),
    .io_wgt_rd_0_data_bits_26_11(tensorGemm_io_wgt_rd_0_data_bits_26_11),
    .io_wgt_rd_0_data_bits_26_12(tensorGemm_io_wgt_rd_0_data_bits_26_12),
    .io_wgt_rd_0_data_bits_26_13(tensorGemm_io_wgt_rd_0_data_bits_26_13),
    .io_wgt_rd_0_data_bits_26_14(tensorGemm_io_wgt_rd_0_data_bits_26_14),
    .io_wgt_rd_0_data_bits_26_15(tensorGemm_io_wgt_rd_0_data_bits_26_15),
    .io_wgt_rd_0_data_bits_27_0(tensorGemm_io_wgt_rd_0_data_bits_27_0),
    .io_wgt_rd_0_data_bits_27_1(tensorGemm_io_wgt_rd_0_data_bits_27_1),
    .io_wgt_rd_0_data_bits_27_2(tensorGemm_io_wgt_rd_0_data_bits_27_2),
    .io_wgt_rd_0_data_bits_27_3(tensorGemm_io_wgt_rd_0_data_bits_27_3),
    .io_wgt_rd_0_data_bits_27_4(tensorGemm_io_wgt_rd_0_data_bits_27_4),
    .io_wgt_rd_0_data_bits_27_5(tensorGemm_io_wgt_rd_0_data_bits_27_5),
    .io_wgt_rd_0_data_bits_27_6(tensorGemm_io_wgt_rd_0_data_bits_27_6),
    .io_wgt_rd_0_data_bits_27_7(tensorGemm_io_wgt_rd_0_data_bits_27_7),
    .io_wgt_rd_0_data_bits_27_8(tensorGemm_io_wgt_rd_0_data_bits_27_8),
    .io_wgt_rd_0_data_bits_27_9(tensorGemm_io_wgt_rd_0_data_bits_27_9),
    .io_wgt_rd_0_data_bits_27_10(tensorGemm_io_wgt_rd_0_data_bits_27_10),
    .io_wgt_rd_0_data_bits_27_11(tensorGemm_io_wgt_rd_0_data_bits_27_11),
    .io_wgt_rd_0_data_bits_27_12(tensorGemm_io_wgt_rd_0_data_bits_27_12),
    .io_wgt_rd_0_data_bits_27_13(tensorGemm_io_wgt_rd_0_data_bits_27_13),
    .io_wgt_rd_0_data_bits_27_14(tensorGemm_io_wgt_rd_0_data_bits_27_14),
    .io_wgt_rd_0_data_bits_27_15(tensorGemm_io_wgt_rd_0_data_bits_27_15),
    .io_wgt_rd_0_data_bits_28_0(tensorGemm_io_wgt_rd_0_data_bits_28_0),
    .io_wgt_rd_0_data_bits_28_1(tensorGemm_io_wgt_rd_0_data_bits_28_1),
    .io_wgt_rd_0_data_bits_28_2(tensorGemm_io_wgt_rd_0_data_bits_28_2),
    .io_wgt_rd_0_data_bits_28_3(tensorGemm_io_wgt_rd_0_data_bits_28_3),
    .io_wgt_rd_0_data_bits_28_4(tensorGemm_io_wgt_rd_0_data_bits_28_4),
    .io_wgt_rd_0_data_bits_28_5(tensorGemm_io_wgt_rd_0_data_bits_28_5),
    .io_wgt_rd_0_data_bits_28_6(tensorGemm_io_wgt_rd_0_data_bits_28_6),
    .io_wgt_rd_0_data_bits_28_7(tensorGemm_io_wgt_rd_0_data_bits_28_7),
    .io_wgt_rd_0_data_bits_28_8(tensorGemm_io_wgt_rd_0_data_bits_28_8),
    .io_wgt_rd_0_data_bits_28_9(tensorGemm_io_wgt_rd_0_data_bits_28_9),
    .io_wgt_rd_0_data_bits_28_10(tensorGemm_io_wgt_rd_0_data_bits_28_10),
    .io_wgt_rd_0_data_bits_28_11(tensorGemm_io_wgt_rd_0_data_bits_28_11),
    .io_wgt_rd_0_data_bits_28_12(tensorGemm_io_wgt_rd_0_data_bits_28_12),
    .io_wgt_rd_0_data_bits_28_13(tensorGemm_io_wgt_rd_0_data_bits_28_13),
    .io_wgt_rd_0_data_bits_28_14(tensorGemm_io_wgt_rd_0_data_bits_28_14),
    .io_wgt_rd_0_data_bits_28_15(tensorGemm_io_wgt_rd_0_data_bits_28_15),
    .io_wgt_rd_0_data_bits_29_0(tensorGemm_io_wgt_rd_0_data_bits_29_0),
    .io_wgt_rd_0_data_bits_29_1(tensorGemm_io_wgt_rd_0_data_bits_29_1),
    .io_wgt_rd_0_data_bits_29_2(tensorGemm_io_wgt_rd_0_data_bits_29_2),
    .io_wgt_rd_0_data_bits_29_3(tensorGemm_io_wgt_rd_0_data_bits_29_3),
    .io_wgt_rd_0_data_bits_29_4(tensorGemm_io_wgt_rd_0_data_bits_29_4),
    .io_wgt_rd_0_data_bits_29_5(tensorGemm_io_wgt_rd_0_data_bits_29_5),
    .io_wgt_rd_0_data_bits_29_6(tensorGemm_io_wgt_rd_0_data_bits_29_6),
    .io_wgt_rd_0_data_bits_29_7(tensorGemm_io_wgt_rd_0_data_bits_29_7),
    .io_wgt_rd_0_data_bits_29_8(tensorGemm_io_wgt_rd_0_data_bits_29_8),
    .io_wgt_rd_0_data_bits_29_9(tensorGemm_io_wgt_rd_0_data_bits_29_9),
    .io_wgt_rd_0_data_bits_29_10(tensorGemm_io_wgt_rd_0_data_bits_29_10),
    .io_wgt_rd_0_data_bits_29_11(tensorGemm_io_wgt_rd_0_data_bits_29_11),
    .io_wgt_rd_0_data_bits_29_12(tensorGemm_io_wgt_rd_0_data_bits_29_12),
    .io_wgt_rd_0_data_bits_29_13(tensorGemm_io_wgt_rd_0_data_bits_29_13),
    .io_wgt_rd_0_data_bits_29_14(tensorGemm_io_wgt_rd_0_data_bits_29_14),
    .io_wgt_rd_0_data_bits_29_15(tensorGemm_io_wgt_rd_0_data_bits_29_15),
    .io_wgt_rd_0_data_bits_30_0(tensorGemm_io_wgt_rd_0_data_bits_30_0),
    .io_wgt_rd_0_data_bits_30_1(tensorGemm_io_wgt_rd_0_data_bits_30_1),
    .io_wgt_rd_0_data_bits_30_2(tensorGemm_io_wgt_rd_0_data_bits_30_2),
    .io_wgt_rd_0_data_bits_30_3(tensorGemm_io_wgt_rd_0_data_bits_30_3),
    .io_wgt_rd_0_data_bits_30_4(tensorGemm_io_wgt_rd_0_data_bits_30_4),
    .io_wgt_rd_0_data_bits_30_5(tensorGemm_io_wgt_rd_0_data_bits_30_5),
    .io_wgt_rd_0_data_bits_30_6(tensorGemm_io_wgt_rd_0_data_bits_30_6),
    .io_wgt_rd_0_data_bits_30_7(tensorGemm_io_wgt_rd_0_data_bits_30_7),
    .io_wgt_rd_0_data_bits_30_8(tensorGemm_io_wgt_rd_0_data_bits_30_8),
    .io_wgt_rd_0_data_bits_30_9(tensorGemm_io_wgt_rd_0_data_bits_30_9),
    .io_wgt_rd_0_data_bits_30_10(tensorGemm_io_wgt_rd_0_data_bits_30_10),
    .io_wgt_rd_0_data_bits_30_11(tensorGemm_io_wgt_rd_0_data_bits_30_11),
    .io_wgt_rd_0_data_bits_30_12(tensorGemm_io_wgt_rd_0_data_bits_30_12),
    .io_wgt_rd_0_data_bits_30_13(tensorGemm_io_wgt_rd_0_data_bits_30_13),
    .io_wgt_rd_0_data_bits_30_14(tensorGemm_io_wgt_rd_0_data_bits_30_14),
    .io_wgt_rd_0_data_bits_30_15(tensorGemm_io_wgt_rd_0_data_bits_30_15),
    .io_wgt_rd_0_data_bits_31_0(tensorGemm_io_wgt_rd_0_data_bits_31_0),
    .io_wgt_rd_0_data_bits_31_1(tensorGemm_io_wgt_rd_0_data_bits_31_1),
    .io_wgt_rd_0_data_bits_31_2(tensorGemm_io_wgt_rd_0_data_bits_31_2),
    .io_wgt_rd_0_data_bits_31_3(tensorGemm_io_wgt_rd_0_data_bits_31_3),
    .io_wgt_rd_0_data_bits_31_4(tensorGemm_io_wgt_rd_0_data_bits_31_4),
    .io_wgt_rd_0_data_bits_31_5(tensorGemm_io_wgt_rd_0_data_bits_31_5),
    .io_wgt_rd_0_data_bits_31_6(tensorGemm_io_wgt_rd_0_data_bits_31_6),
    .io_wgt_rd_0_data_bits_31_7(tensorGemm_io_wgt_rd_0_data_bits_31_7),
    .io_wgt_rd_0_data_bits_31_8(tensorGemm_io_wgt_rd_0_data_bits_31_8),
    .io_wgt_rd_0_data_bits_31_9(tensorGemm_io_wgt_rd_0_data_bits_31_9),
    .io_wgt_rd_0_data_bits_31_10(tensorGemm_io_wgt_rd_0_data_bits_31_10),
    .io_wgt_rd_0_data_bits_31_11(tensorGemm_io_wgt_rd_0_data_bits_31_11),
    .io_wgt_rd_0_data_bits_31_12(tensorGemm_io_wgt_rd_0_data_bits_31_12),
    .io_wgt_rd_0_data_bits_31_13(tensorGemm_io_wgt_rd_0_data_bits_31_13),
    .io_wgt_rd_0_data_bits_31_14(tensorGemm_io_wgt_rd_0_data_bits_31_14),
    .io_wgt_rd_0_data_bits_31_15(tensorGemm_io_wgt_rd_0_data_bits_31_15),
    .io_acc_rd_0_idx_valid(tensorGemm_io_acc_rd_0_idx_valid),
    .io_acc_rd_0_idx_bits(tensorGemm_io_acc_rd_0_idx_bits),
    .io_acc_rd_0_data_valid(tensorGemm_io_acc_rd_0_data_valid),
    .io_acc_rd_0_data_bits_0_0(tensorGemm_io_acc_rd_0_data_bits_0_0),
    .io_acc_rd_0_data_bits_0_1(tensorGemm_io_acc_rd_0_data_bits_0_1),
    .io_acc_rd_0_data_bits_0_2(tensorGemm_io_acc_rd_0_data_bits_0_2),
    .io_acc_rd_0_data_bits_0_3(tensorGemm_io_acc_rd_0_data_bits_0_3),
    .io_acc_rd_0_data_bits_0_4(tensorGemm_io_acc_rd_0_data_bits_0_4),
    .io_acc_rd_0_data_bits_0_5(tensorGemm_io_acc_rd_0_data_bits_0_5),
    .io_acc_rd_0_data_bits_0_6(tensorGemm_io_acc_rd_0_data_bits_0_6),
    .io_acc_rd_0_data_bits_0_7(tensorGemm_io_acc_rd_0_data_bits_0_7),
    .io_acc_rd_0_data_bits_0_8(tensorGemm_io_acc_rd_0_data_bits_0_8),
    .io_acc_rd_0_data_bits_0_9(tensorGemm_io_acc_rd_0_data_bits_0_9),
    .io_acc_rd_0_data_bits_0_10(tensorGemm_io_acc_rd_0_data_bits_0_10),
    .io_acc_rd_0_data_bits_0_11(tensorGemm_io_acc_rd_0_data_bits_0_11),
    .io_acc_rd_0_data_bits_0_12(tensorGemm_io_acc_rd_0_data_bits_0_12),
    .io_acc_rd_0_data_bits_0_13(tensorGemm_io_acc_rd_0_data_bits_0_13),
    .io_acc_rd_0_data_bits_0_14(tensorGemm_io_acc_rd_0_data_bits_0_14),
    .io_acc_rd_0_data_bits_0_15(tensorGemm_io_acc_rd_0_data_bits_0_15),
    .io_acc_rd_0_data_bits_0_16(tensorGemm_io_acc_rd_0_data_bits_0_16),
    .io_acc_rd_0_data_bits_0_17(tensorGemm_io_acc_rd_0_data_bits_0_17),
    .io_acc_rd_0_data_bits_0_18(tensorGemm_io_acc_rd_0_data_bits_0_18),
    .io_acc_rd_0_data_bits_0_19(tensorGemm_io_acc_rd_0_data_bits_0_19),
    .io_acc_rd_0_data_bits_0_20(tensorGemm_io_acc_rd_0_data_bits_0_20),
    .io_acc_rd_0_data_bits_0_21(tensorGemm_io_acc_rd_0_data_bits_0_21),
    .io_acc_rd_0_data_bits_0_22(tensorGemm_io_acc_rd_0_data_bits_0_22),
    .io_acc_rd_0_data_bits_0_23(tensorGemm_io_acc_rd_0_data_bits_0_23),
    .io_acc_rd_0_data_bits_0_24(tensorGemm_io_acc_rd_0_data_bits_0_24),
    .io_acc_rd_0_data_bits_0_25(tensorGemm_io_acc_rd_0_data_bits_0_25),
    .io_acc_rd_0_data_bits_0_26(tensorGemm_io_acc_rd_0_data_bits_0_26),
    .io_acc_rd_0_data_bits_0_27(tensorGemm_io_acc_rd_0_data_bits_0_27),
    .io_acc_rd_0_data_bits_0_28(tensorGemm_io_acc_rd_0_data_bits_0_28),
    .io_acc_rd_0_data_bits_0_29(tensorGemm_io_acc_rd_0_data_bits_0_29),
    .io_acc_rd_0_data_bits_0_30(tensorGemm_io_acc_rd_0_data_bits_0_30),
    .io_acc_rd_0_data_bits_0_31(tensorGemm_io_acc_rd_0_data_bits_0_31),
    .io_acc_wr_0_valid(tensorGemm_io_acc_wr_0_valid),
    .io_acc_wr_0_bits_idx(tensorGemm_io_acc_wr_0_bits_idx),
    .io_acc_wr_0_bits_data_0_0(tensorGemm_io_acc_wr_0_bits_data_0_0),
    .io_acc_wr_0_bits_data_0_1(tensorGemm_io_acc_wr_0_bits_data_0_1),
    .io_acc_wr_0_bits_data_0_2(tensorGemm_io_acc_wr_0_bits_data_0_2),
    .io_acc_wr_0_bits_data_0_3(tensorGemm_io_acc_wr_0_bits_data_0_3),
    .io_acc_wr_0_bits_data_0_4(tensorGemm_io_acc_wr_0_bits_data_0_4),
    .io_acc_wr_0_bits_data_0_5(tensorGemm_io_acc_wr_0_bits_data_0_5),
    .io_acc_wr_0_bits_data_0_6(tensorGemm_io_acc_wr_0_bits_data_0_6),
    .io_acc_wr_0_bits_data_0_7(tensorGemm_io_acc_wr_0_bits_data_0_7),
    .io_acc_wr_0_bits_data_0_8(tensorGemm_io_acc_wr_0_bits_data_0_8),
    .io_acc_wr_0_bits_data_0_9(tensorGemm_io_acc_wr_0_bits_data_0_9),
    .io_acc_wr_0_bits_data_0_10(tensorGemm_io_acc_wr_0_bits_data_0_10),
    .io_acc_wr_0_bits_data_0_11(tensorGemm_io_acc_wr_0_bits_data_0_11),
    .io_acc_wr_0_bits_data_0_12(tensorGemm_io_acc_wr_0_bits_data_0_12),
    .io_acc_wr_0_bits_data_0_13(tensorGemm_io_acc_wr_0_bits_data_0_13),
    .io_acc_wr_0_bits_data_0_14(tensorGemm_io_acc_wr_0_bits_data_0_14),
    .io_acc_wr_0_bits_data_0_15(tensorGemm_io_acc_wr_0_bits_data_0_15),
    .io_acc_wr_0_bits_data_0_16(tensorGemm_io_acc_wr_0_bits_data_0_16),
    .io_acc_wr_0_bits_data_0_17(tensorGemm_io_acc_wr_0_bits_data_0_17),
    .io_acc_wr_0_bits_data_0_18(tensorGemm_io_acc_wr_0_bits_data_0_18),
    .io_acc_wr_0_bits_data_0_19(tensorGemm_io_acc_wr_0_bits_data_0_19),
    .io_acc_wr_0_bits_data_0_20(tensorGemm_io_acc_wr_0_bits_data_0_20),
    .io_acc_wr_0_bits_data_0_21(tensorGemm_io_acc_wr_0_bits_data_0_21),
    .io_acc_wr_0_bits_data_0_22(tensorGemm_io_acc_wr_0_bits_data_0_22),
    .io_acc_wr_0_bits_data_0_23(tensorGemm_io_acc_wr_0_bits_data_0_23),
    .io_acc_wr_0_bits_data_0_24(tensorGemm_io_acc_wr_0_bits_data_0_24),
    .io_acc_wr_0_bits_data_0_25(tensorGemm_io_acc_wr_0_bits_data_0_25),
    .io_acc_wr_0_bits_data_0_26(tensorGemm_io_acc_wr_0_bits_data_0_26),
    .io_acc_wr_0_bits_data_0_27(tensorGemm_io_acc_wr_0_bits_data_0_27),
    .io_acc_wr_0_bits_data_0_28(tensorGemm_io_acc_wr_0_bits_data_0_28),
    .io_acc_wr_0_bits_data_0_29(tensorGemm_io_acc_wr_0_bits_data_0_29),
    .io_acc_wr_0_bits_data_0_30(tensorGemm_io_acc_wr_0_bits_data_0_30),
    .io_acc_wr_0_bits_data_0_31(tensorGemm_io_acc_wr_0_bits_data_0_31),
    .io_out_rd_0_data_valid(tensorGemm_io_out_rd_0_data_valid),
    .io_out_wr_0_valid(tensorGemm_io_out_wr_0_valid),
    .io_out_wr_0_bits_idx(tensorGemm_io_out_wr_0_bits_idx),
    .io_out_wr_0_bits_data_0_0(tensorGemm_io_out_wr_0_bits_data_0_0),
    .io_out_wr_0_bits_data_0_1(tensorGemm_io_out_wr_0_bits_data_0_1),
    .io_out_wr_0_bits_data_0_2(tensorGemm_io_out_wr_0_bits_data_0_2),
    .io_out_wr_0_bits_data_0_3(tensorGemm_io_out_wr_0_bits_data_0_3),
    .io_out_wr_0_bits_data_0_4(tensorGemm_io_out_wr_0_bits_data_0_4),
    .io_out_wr_0_bits_data_0_5(tensorGemm_io_out_wr_0_bits_data_0_5),
    .io_out_wr_0_bits_data_0_6(tensorGemm_io_out_wr_0_bits_data_0_6),
    .io_out_wr_0_bits_data_0_7(tensorGemm_io_out_wr_0_bits_data_0_7),
    .io_out_wr_0_bits_data_0_8(tensorGemm_io_out_wr_0_bits_data_0_8),
    .io_out_wr_0_bits_data_0_9(tensorGemm_io_out_wr_0_bits_data_0_9),
    .io_out_wr_0_bits_data_0_10(tensorGemm_io_out_wr_0_bits_data_0_10),
    .io_out_wr_0_bits_data_0_11(tensorGemm_io_out_wr_0_bits_data_0_11),
    .io_out_wr_0_bits_data_0_12(tensorGemm_io_out_wr_0_bits_data_0_12),
    .io_out_wr_0_bits_data_0_13(tensorGemm_io_out_wr_0_bits_data_0_13),
    .io_out_wr_0_bits_data_0_14(tensorGemm_io_out_wr_0_bits_data_0_14),
    .io_out_wr_0_bits_data_0_15(tensorGemm_io_out_wr_0_bits_data_0_15),
    .io_out_wr_0_bits_data_0_16(tensorGemm_io_out_wr_0_bits_data_0_16),
    .io_out_wr_0_bits_data_0_17(tensorGemm_io_out_wr_0_bits_data_0_17),
    .io_out_wr_0_bits_data_0_18(tensorGemm_io_out_wr_0_bits_data_0_18),
    .io_out_wr_0_bits_data_0_19(tensorGemm_io_out_wr_0_bits_data_0_19),
    .io_out_wr_0_bits_data_0_20(tensorGemm_io_out_wr_0_bits_data_0_20),
    .io_out_wr_0_bits_data_0_21(tensorGemm_io_out_wr_0_bits_data_0_21),
    .io_out_wr_0_bits_data_0_22(tensorGemm_io_out_wr_0_bits_data_0_22),
    .io_out_wr_0_bits_data_0_23(tensorGemm_io_out_wr_0_bits_data_0_23),
    .io_out_wr_0_bits_data_0_24(tensorGemm_io_out_wr_0_bits_data_0_24),
    .io_out_wr_0_bits_data_0_25(tensorGemm_io_out_wr_0_bits_data_0_25),
    .io_out_wr_0_bits_data_0_26(tensorGemm_io_out_wr_0_bits_data_0_26),
    .io_out_wr_0_bits_data_0_27(tensorGemm_io_out_wr_0_bits_data_0_27),
    .io_out_wr_0_bits_data_0_28(tensorGemm_io_out_wr_0_bits_data_0_28),
    .io_out_wr_0_bits_data_0_29(tensorGemm_io_out_wr_0_bits_data_0_29),
    .io_out_wr_0_bits_data_0_30(tensorGemm_io_out_wr_0_bits_data_0_30),
    .io_out_wr_0_bits_data_0_31(tensorGemm_io_out_wr_0_bits_data_0_31)
  );
  TensorAlu tensorAlu ( // @[Compute.scala 64:25]
    .clock(tensorAlu_clock),
    .reset(tensorAlu_reset),
    .io_start(tensorAlu_io_start),
    .io_done(tensorAlu_io_done),
    .io_dec_alu_imm(tensorAlu_io_dec_alu_imm),
    .io_dec_alu_use_imm(tensorAlu_io_dec_alu_use_imm),
    .io_dec_alu_op(tensorAlu_io_dec_alu_op),
    .io_dec_src_1(tensorAlu_io_dec_src_1),
    .io_dec_src_0(tensorAlu_io_dec_src_0),
    .io_dec_dst_1(tensorAlu_io_dec_dst_1),
    .io_dec_dst_0(tensorAlu_io_dec_dst_0),
    .io_dec_lp_1(tensorAlu_io_dec_lp_1),
    .io_dec_lp_0(tensorAlu_io_dec_lp_0),
    .io_dec_uop_end(tensorAlu_io_dec_uop_end),
    .io_dec_uop_begin(tensorAlu_io_dec_uop_begin),
    .io_uop_idx_valid(tensorAlu_io_uop_idx_valid),
    .io_uop_idx_bits(tensorAlu_io_uop_idx_bits),
    .io_uop_data_bits_u2(tensorAlu_io_uop_data_bits_u2),
    .io_uop_data_bits_u1(tensorAlu_io_uop_data_bits_u1),
    .io_uop_data_bits_u0(tensorAlu_io_uop_data_bits_u0),
    .io_acc_rd_0_idx_valid(tensorAlu_io_acc_rd_0_idx_valid),
    .io_acc_rd_0_idx_bits(tensorAlu_io_acc_rd_0_idx_bits),
    .io_acc_rd_0_data_valid(tensorAlu_io_acc_rd_0_data_valid),
    .io_acc_rd_0_data_bits_0_0(tensorAlu_io_acc_rd_0_data_bits_0_0),
    .io_acc_rd_0_data_bits_0_1(tensorAlu_io_acc_rd_0_data_bits_0_1),
    .io_acc_rd_0_data_bits_0_2(tensorAlu_io_acc_rd_0_data_bits_0_2),
    .io_acc_rd_0_data_bits_0_3(tensorAlu_io_acc_rd_0_data_bits_0_3),
    .io_acc_rd_0_data_bits_0_4(tensorAlu_io_acc_rd_0_data_bits_0_4),
    .io_acc_rd_0_data_bits_0_5(tensorAlu_io_acc_rd_0_data_bits_0_5),
    .io_acc_rd_0_data_bits_0_6(tensorAlu_io_acc_rd_0_data_bits_0_6),
    .io_acc_rd_0_data_bits_0_7(tensorAlu_io_acc_rd_0_data_bits_0_7),
    .io_acc_rd_0_data_bits_0_8(tensorAlu_io_acc_rd_0_data_bits_0_8),
    .io_acc_rd_0_data_bits_0_9(tensorAlu_io_acc_rd_0_data_bits_0_9),
    .io_acc_rd_0_data_bits_0_10(tensorAlu_io_acc_rd_0_data_bits_0_10),
    .io_acc_rd_0_data_bits_0_11(tensorAlu_io_acc_rd_0_data_bits_0_11),
    .io_acc_rd_0_data_bits_0_12(tensorAlu_io_acc_rd_0_data_bits_0_12),
    .io_acc_rd_0_data_bits_0_13(tensorAlu_io_acc_rd_0_data_bits_0_13),
    .io_acc_rd_0_data_bits_0_14(tensorAlu_io_acc_rd_0_data_bits_0_14),
    .io_acc_rd_0_data_bits_0_15(tensorAlu_io_acc_rd_0_data_bits_0_15),
    .io_acc_rd_0_data_bits_0_16(tensorAlu_io_acc_rd_0_data_bits_0_16),
    .io_acc_rd_0_data_bits_0_17(tensorAlu_io_acc_rd_0_data_bits_0_17),
    .io_acc_rd_0_data_bits_0_18(tensorAlu_io_acc_rd_0_data_bits_0_18),
    .io_acc_rd_0_data_bits_0_19(tensorAlu_io_acc_rd_0_data_bits_0_19),
    .io_acc_rd_0_data_bits_0_20(tensorAlu_io_acc_rd_0_data_bits_0_20),
    .io_acc_rd_0_data_bits_0_21(tensorAlu_io_acc_rd_0_data_bits_0_21),
    .io_acc_rd_0_data_bits_0_22(tensorAlu_io_acc_rd_0_data_bits_0_22),
    .io_acc_rd_0_data_bits_0_23(tensorAlu_io_acc_rd_0_data_bits_0_23),
    .io_acc_rd_0_data_bits_0_24(tensorAlu_io_acc_rd_0_data_bits_0_24),
    .io_acc_rd_0_data_bits_0_25(tensorAlu_io_acc_rd_0_data_bits_0_25),
    .io_acc_rd_0_data_bits_0_26(tensorAlu_io_acc_rd_0_data_bits_0_26),
    .io_acc_rd_0_data_bits_0_27(tensorAlu_io_acc_rd_0_data_bits_0_27),
    .io_acc_rd_0_data_bits_0_28(tensorAlu_io_acc_rd_0_data_bits_0_28),
    .io_acc_rd_0_data_bits_0_29(tensorAlu_io_acc_rd_0_data_bits_0_29),
    .io_acc_rd_0_data_bits_0_30(tensorAlu_io_acc_rd_0_data_bits_0_30),
    .io_acc_rd_0_data_bits_0_31(tensorAlu_io_acc_rd_0_data_bits_0_31),
    .io_acc_wr_0_valid(tensorAlu_io_acc_wr_0_valid),
    .io_acc_wr_0_bits_idx(tensorAlu_io_acc_wr_0_bits_idx),
    .io_acc_wr_0_bits_data_0_0(tensorAlu_io_acc_wr_0_bits_data_0_0),
    .io_acc_wr_0_bits_data_0_1(tensorAlu_io_acc_wr_0_bits_data_0_1),
    .io_acc_wr_0_bits_data_0_2(tensorAlu_io_acc_wr_0_bits_data_0_2),
    .io_acc_wr_0_bits_data_0_3(tensorAlu_io_acc_wr_0_bits_data_0_3),
    .io_acc_wr_0_bits_data_0_4(tensorAlu_io_acc_wr_0_bits_data_0_4),
    .io_acc_wr_0_bits_data_0_5(tensorAlu_io_acc_wr_0_bits_data_0_5),
    .io_acc_wr_0_bits_data_0_6(tensorAlu_io_acc_wr_0_bits_data_0_6),
    .io_acc_wr_0_bits_data_0_7(tensorAlu_io_acc_wr_0_bits_data_0_7),
    .io_acc_wr_0_bits_data_0_8(tensorAlu_io_acc_wr_0_bits_data_0_8),
    .io_acc_wr_0_bits_data_0_9(tensorAlu_io_acc_wr_0_bits_data_0_9),
    .io_acc_wr_0_bits_data_0_10(tensorAlu_io_acc_wr_0_bits_data_0_10),
    .io_acc_wr_0_bits_data_0_11(tensorAlu_io_acc_wr_0_bits_data_0_11),
    .io_acc_wr_0_bits_data_0_12(tensorAlu_io_acc_wr_0_bits_data_0_12),
    .io_acc_wr_0_bits_data_0_13(tensorAlu_io_acc_wr_0_bits_data_0_13),
    .io_acc_wr_0_bits_data_0_14(tensorAlu_io_acc_wr_0_bits_data_0_14),
    .io_acc_wr_0_bits_data_0_15(tensorAlu_io_acc_wr_0_bits_data_0_15),
    .io_acc_wr_0_bits_data_0_16(tensorAlu_io_acc_wr_0_bits_data_0_16),
    .io_acc_wr_0_bits_data_0_17(tensorAlu_io_acc_wr_0_bits_data_0_17),
    .io_acc_wr_0_bits_data_0_18(tensorAlu_io_acc_wr_0_bits_data_0_18),
    .io_acc_wr_0_bits_data_0_19(tensorAlu_io_acc_wr_0_bits_data_0_19),
    .io_acc_wr_0_bits_data_0_20(tensorAlu_io_acc_wr_0_bits_data_0_20),
    .io_acc_wr_0_bits_data_0_21(tensorAlu_io_acc_wr_0_bits_data_0_21),
    .io_acc_wr_0_bits_data_0_22(tensorAlu_io_acc_wr_0_bits_data_0_22),
    .io_acc_wr_0_bits_data_0_23(tensorAlu_io_acc_wr_0_bits_data_0_23),
    .io_acc_wr_0_bits_data_0_24(tensorAlu_io_acc_wr_0_bits_data_0_24),
    .io_acc_wr_0_bits_data_0_25(tensorAlu_io_acc_wr_0_bits_data_0_25),
    .io_acc_wr_0_bits_data_0_26(tensorAlu_io_acc_wr_0_bits_data_0_26),
    .io_acc_wr_0_bits_data_0_27(tensorAlu_io_acc_wr_0_bits_data_0_27),
    .io_acc_wr_0_bits_data_0_28(tensorAlu_io_acc_wr_0_bits_data_0_28),
    .io_acc_wr_0_bits_data_0_29(tensorAlu_io_acc_wr_0_bits_data_0_29),
    .io_acc_wr_0_bits_data_0_30(tensorAlu_io_acc_wr_0_bits_data_0_30),
    .io_acc_wr_0_bits_data_0_31(tensorAlu_io_acc_wr_0_bits_data_0_31),
    .io_out_rd_0_data_valid(tensorAlu_io_out_rd_0_data_valid),
    .io_out_wr_0_valid(tensorAlu_io_out_wr_0_valid),
    .io_out_wr_0_bits_idx(tensorAlu_io_out_wr_0_bits_idx),
    .io_out_wr_0_bits_data_0_0(tensorAlu_io_out_wr_0_bits_data_0_0),
    .io_out_wr_0_bits_data_0_1(tensorAlu_io_out_wr_0_bits_data_0_1),
    .io_out_wr_0_bits_data_0_2(tensorAlu_io_out_wr_0_bits_data_0_2),
    .io_out_wr_0_bits_data_0_3(tensorAlu_io_out_wr_0_bits_data_0_3),
    .io_out_wr_0_bits_data_0_4(tensorAlu_io_out_wr_0_bits_data_0_4),
    .io_out_wr_0_bits_data_0_5(tensorAlu_io_out_wr_0_bits_data_0_5),
    .io_out_wr_0_bits_data_0_6(tensorAlu_io_out_wr_0_bits_data_0_6),
    .io_out_wr_0_bits_data_0_7(tensorAlu_io_out_wr_0_bits_data_0_7),
    .io_out_wr_0_bits_data_0_8(tensorAlu_io_out_wr_0_bits_data_0_8),
    .io_out_wr_0_bits_data_0_9(tensorAlu_io_out_wr_0_bits_data_0_9),
    .io_out_wr_0_bits_data_0_10(tensorAlu_io_out_wr_0_bits_data_0_10),
    .io_out_wr_0_bits_data_0_11(tensorAlu_io_out_wr_0_bits_data_0_11),
    .io_out_wr_0_bits_data_0_12(tensorAlu_io_out_wr_0_bits_data_0_12),
    .io_out_wr_0_bits_data_0_13(tensorAlu_io_out_wr_0_bits_data_0_13),
    .io_out_wr_0_bits_data_0_14(tensorAlu_io_out_wr_0_bits_data_0_14),
    .io_out_wr_0_bits_data_0_15(tensorAlu_io_out_wr_0_bits_data_0_15),
    .io_out_wr_0_bits_data_0_16(tensorAlu_io_out_wr_0_bits_data_0_16),
    .io_out_wr_0_bits_data_0_17(tensorAlu_io_out_wr_0_bits_data_0_17),
    .io_out_wr_0_bits_data_0_18(tensorAlu_io_out_wr_0_bits_data_0_18),
    .io_out_wr_0_bits_data_0_19(tensorAlu_io_out_wr_0_bits_data_0_19),
    .io_out_wr_0_bits_data_0_20(tensorAlu_io_out_wr_0_bits_data_0_20),
    .io_out_wr_0_bits_data_0_21(tensorAlu_io_out_wr_0_bits_data_0_21),
    .io_out_wr_0_bits_data_0_22(tensorAlu_io_out_wr_0_bits_data_0_22),
    .io_out_wr_0_bits_data_0_23(tensorAlu_io_out_wr_0_bits_data_0_23),
    .io_out_wr_0_bits_data_0_24(tensorAlu_io_out_wr_0_bits_data_0_24),
    .io_out_wr_0_bits_data_0_25(tensorAlu_io_out_wr_0_bits_data_0_25),
    .io_out_wr_0_bits_data_0_26(tensorAlu_io_out_wr_0_bits_data_0_26),
    .io_out_wr_0_bits_data_0_27(tensorAlu_io_out_wr_0_bits_data_0_27),
    .io_out_wr_0_bits_data_0_28(tensorAlu_io_out_wr_0_bits_data_0_28),
    .io_out_wr_0_bits_data_0_29(tensorAlu_io_out_wr_0_bits_data_0_29),
    .io_out_wr_0_bits_data_0_30(tensorAlu_io_out_wr_0_bits_data_0_30),
    .io_out_wr_0_bits_data_0_31(tensorAlu_io_out_wr_0_bits_data_0_31)
  );
  SyncQueue_1 inst_q ( // @[Compute.scala 69:22]
    .clock(inst_q_clock),
    .reset(inst_q_reset),
    .io_enq_ready(inst_q_io_enq_ready),
    .io_enq_valid(inst_q_io_enq_valid),
    .io_enq_bits(inst_q_io_enq_bits),
    .io_deq_ready(inst_q_io_deq_ready),
    .io_deq_valid(inst_q_io_deq_valid),
    .io_deq_bits(inst_q_io_deq_bits)
  );
  ComputeDecode dec ( // @[Compute.scala 72:19]
    .io_inst(dec_io_inst),
    .io_push_next(dec_io_push_next),
    .io_push_prev(dec_io_push_prev),
    .io_pop_next(dec_io_pop_next),
    .io_pop_prev(dec_io_pop_prev),
    .io_isLoadAcc(dec_io_isLoadAcc),
    .io_isLoadUop(dec_io_isLoadUop),
    .io_isSync(dec_io_isSync),
    .io_isAlu(dec_io_isAlu),
    .io_isGemm(dec_io_isGemm),
    .io_isFinish(dec_io_isFinish)
  );
  assign io_o_post_0 = dec_io_push_prev & _inst_q_io_deq_ready_T_3; // @[Compute.scala 230:36]
  assign io_o_post_1 = dec_io_push_next & _inst_q_io_deq_ready_T_3; // @[Compute.scala 231:36]
  assign io_inst_ready = inst_q_io_enq_ready; // @[Compute.scala 120:17]
  assign io_vme_rd_0_cmd_valid = loadUop_io_vme_rd_cmd_valid; // @[Compute.scala 127:16]
  assign io_vme_rd_0_cmd_bits_addr = loadUop_io_vme_rd_cmd_bits_addr; // @[Compute.scala 127:16]
  assign io_vme_rd_0_cmd_bits_len = loadUop_io_vme_rd_cmd_bits_len; // @[Compute.scala 127:16]
  assign io_vme_rd_0_cmd_bits_tag = loadUop_io_vme_rd_cmd_bits_tag; // @[Compute.scala 127:16]
  assign io_vme_rd_1_cmd_valid = tensorAcc_io_vme_rd_cmd_valid; // @[Compute.scala 158:16]
  assign io_vme_rd_1_cmd_bits_addr = tensorAcc_io_vme_rd_cmd_bits_addr; // @[Compute.scala 158:16]
  assign io_vme_rd_1_cmd_bits_len = tensorAcc_io_vme_rd_cmd_bits_len; // @[Compute.scala 158:16]
  assign io_vme_rd_1_cmd_bits_tag = tensorAcc_io_vme_rd_cmd_bits_tag; // @[Compute.scala 158:16]
  assign io_inp_rd_0_idx_valid = tensorGemm_io_inp_rd_0_idx_valid; // @[Compute.scala 166:21]
  assign io_inp_rd_0_idx_bits = tensorGemm_io_inp_rd_0_idx_bits; // @[Compute.scala 166:21]
  assign io_wgt_rd_0_idx_valid = tensorGemm_io_wgt_rd_0_idx_valid; // @[Compute.scala 167:21]
  assign io_wgt_rd_0_idx_bits = tensorGemm_io_wgt_rd_0_idx_bits; // @[Compute.scala 167:21]
  assign io_out_wr_0_valid = io_out_wr_0_valid_REG ? tensorGemm_io_out_wr_0_valid : tensorAlu_io_out_wr_0_valid; // @[Compute.scala 207:28]
  assign io_out_wr_0_bits_idx = io_out_wr_0_bits_idx_REG ? tensorGemm_io_out_wr_0_bits_idx :
    tensorAlu_io_out_wr_0_bits_idx; // @[Compute.scala 209:31]
  assign io_out_wr_0_bits_data_0_0 = outDataBits_0[7:0]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_1 = outDataBits_0[15:8]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_2 = outDataBits_0[23:16]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_3 = outDataBits_0[31:24]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_4 = outDataBits_0[39:32]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_5 = outDataBits_0[47:40]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_6 = outDataBits_0[55:48]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_7 = outDataBits_0[63:56]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_8 = outDataBits_0[71:64]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_9 = outDataBits_0[79:72]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_10 = outDataBits_0[87:80]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_11 = outDataBits_0[95:88]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_12 = outDataBits_0[103:96]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_13 = outDataBits_0[111:104]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_14 = outDataBits_0[119:112]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_15 = outDataBits_0[127:120]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_16 = outDataBits_0[135:128]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_17 = outDataBits_0[143:136]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_18 = outDataBits_0[151:144]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_19 = outDataBits_0[159:152]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_20 = outDataBits_0[167:160]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_21 = outDataBits_0[175:168]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_22 = outDataBits_0[183:176]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_23 = outDataBits_0[191:184]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_24 = outDataBits_0[199:192]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_25 = outDataBits_0[207:200]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_26 = outDataBits_0[215:208]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_27 = outDataBits_0[223:216]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_28 = outDataBits_0[231:224]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_29 = outDataBits_0[239:232]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_30 = outDataBits_0[247:240]; // @[Compute.scala 214:49]
  assign io_out_wr_0_bits_data_0_31 = outDataBits_0[255:248]; // @[Compute.scala 214:49]
  assign io_finish = _inst_q_io_deq_ready_T_1 & dec_io_isFinish; // @[Compute.scala 234:38]
  assign io_acc_wr_event = tensorAcc_io_tensor_wr_0_valid; // @[Compute.scala 159:19]
  assign s_0_clock = clock;
  assign s_0_reset = reset;
  assign s_0_io_spost = io_i_post_0; // @[Compute.scala 226:17]
  assign s_0_io_swait = dec_io_pop_prev & _loadUop_io_start_T_1; // @[Compute.scala 228:36]
  assign s_1_clock = clock;
  assign s_1_reset = reset;
  assign s_1_io_spost = io_i_post_1; // @[Compute.scala 227:17]
  assign s_1_io_swait = dec_io_pop_next & _loadUop_io_start_T_1; // @[Compute.scala 229:36]
  assign loadUop_clock = clock;
  assign loadUop_reset = reset;
  assign loadUop_io_start = state == 2'h0 & start & dec_io_isLoadUop; // @[Compute.scala 124:47]
  assign loadUop_io_inst = inst_q_io_deq_bits; // @[Compute.scala 125:19]
  assign loadUop_io_baddr = io_uop_baddr; // @[Compute.scala 126:20]
  assign loadUop_io_vme_rd_cmd_ready = io_vme_rd_0_cmd_ready; // @[Compute.scala 127:16]
  assign loadUop_io_vme_rd_data_valid = io_vme_rd_0_data_valid; // @[Compute.scala 127:16]
  assign loadUop_io_vme_rd_data_bits_data = io_vme_rd_0_data_bits_data; // @[Compute.scala 127:16]
  assign loadUop_io_vme_rd_data_bits_tag = io_vme_rd_0_data_bits_tag; // @[Compute.scala 127:16]
  assign loadUop_io_vme_rd_data_bits_last = io_vme_rd_0_data_bits_last; // @[Compute.scala 127:16]
  assign loadUop_io_uop_idx_valid = dec_io_isGemm ? tensorGemm_io_uop_idx_valid : tensorAlu_io_uop_idx_valid; // @[Compute.scala 128:28]
  assign loadUop_io_uop_idx_bits = dec_io_isGemm ? tensorGemm_io_uop_idx_bits : tensorAlu_io_uop_idx_bits; // @[Compute.scala 128:28]
  assign tensorAcc_clock = clock;
  assign tensorAcc_reset = reset;
  assign tensorAcc_io_start = _loadUop_io_start_T_1 & dec_io_isLoadAcc; // @[Compute.scala 132:49]
  assign tensorAcc_io_inst = inst_q_io_deq_bits; // @[Compute.scala 133:21]
  assign tensorAcc_io_baddr = io_acc_baddr; // @[Compute.scala 134:22]
  assign tensorAcc_io_vme_rd_cmd_ready = io_vme_rd_1_cmd_ready; // @[Compute.scala 158:16]
  assign tensorAcc_io_vme_rd_data_valid = io_vme_rd_1_data_valid; // @[Compute.scala 158:16]
  assign tensorAcc_io_vme_rd_data_bits_data = io_vme_rd_1_data_bits_data; // @[Compute.scala 158:16]
  assign tensorAcc_io_vme_rd_data_bits_tag = io_vme_rd_1_data_bits_tag; // @[Compute.scala 158:16]
  assign tensorAcc_io_tensor_rd_0_idx_valid = tensorAcc_io_tensor_rd_0_idx_REG ? tensorGemm_io_acc_rd_0_idx_valid :
    tensorAlu_io_acc_rd_0_idx_valid; // @[Compute.scala 149:43]
  assign tensorAcc_io_tensor_rd_0_idx_bits = tensorAcc_io_tensor_rd_0_idx_REG ? tensorGemm_io_acc_rd_0_idx_bits :
    tensorAlu_io_acc_rd_0_idx_bits; // @[Compute.scala 149:43]
  assign tensorAcc_io_tensor_wr_0_valid = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_valid :
    tensorAlu_io_acc_wr_0_valid; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_idx = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_idx :
    tensorAlu_io_acc_wr_0_bits_idx; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_0 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_0 :
    tensorAlu_io_acc_wr_0_bits_data_0_0; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_1 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_1 :
    tensorAlu_io_acc_wr_0_bits_data_0_1; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_2 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_2 :
    tensorAlu_io_acc_wr_0_bits_data_0_2; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_3 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_3 :
    tensorAlu_io_acc_wr_0_bits_data_0_3; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_4 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_4 :
    tensorAlu_io_acc_wr_0_bits_data_0_4; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_5 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_5 :
    tensorAlu_io_acc_wr_0_bits_data_0_5; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_6 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_6 :
    tensorAlu_io_acc_wr_0_bits_data_0_6; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_7 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_7 :
    tensorAlu_io_acc_wr_0_bits_data_0_7; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_8 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_8 :
    tensorAlu_io_acc_wr_0_bits_data_0_8; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_9 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_9 :
    tensorAlu_io_acc_wr_0_bits_data_0_9; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_10 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_10
     : tensorAlu_io_acc_wr_0_bits_data_0_10; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_11 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_11
     : tensorAlu_io_acc_wr_0_bits_data_0_11; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_12 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_12
     : tensorAlu_io_acc_wr_0_bits_data_0_12; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_13 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_13
     : tensorAlu_io_acc_wr_0_bits_data_0_13; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_14 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_14
     : tensorAlu_io_acc_wr_0_bits_data_0_14; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_15 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_15
     : tensorAlu_io_acc_wr_0_bits_data_0_15; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_16 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_16
     : tensorAlu_io_acc_wr_0_bits_data_0_16; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_17 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_17
     : tensorAlu_io_acc_wr_0_bits_data_0_17; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_18 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_18
     : tensorAlu_io_acc_wr_0_bits_data_0_18; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_19 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_19
     : tensorAlu_io_acc_wr_0_bits_data_0_19; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_20 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_20
     : tensorAlu_io_acc_wr_0_bits_data_0_20; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_21 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_21
     : tensorAlu_io_acc_wr_0_bits_data_0_21; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_22 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_22
     : tensorAlu_io_acc_wr_0_bits_data_0_22; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_23 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_23
     : tensorAlu_io_acc_wr_0_bits_data_0_23; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_24 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_24
     : tensorAlu_io_acc_wr_0_bits_data_0_24; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_25 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_25
     : tensorAlu_io_acc_wr_0_bits_data_0_25; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_26 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_26
     : tensorAlu_io_acc_wr_0_bits_data_0_26; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_27 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_27
     : tensorAlu_io_acc_wr_0_bits_data_0_27; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_28 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_28
     : tensorAlu_io_acc_wr_0_bits_data_0_28; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_29 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_29
     : tensorAlu_io_acc_wr_0_bits_data_0_29; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_30 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_30
     : tensorAlu_io_acc_wr_0_bits_data_0_30; // @[Compute.scala 153:39]
  assign tensorAcc_io_tensor_wr_0_bits_data_0_31 = tensorAcc_io_tensor_wr_0_REG ? tensorGemm_io_acc_wr_0_bits_data_0_31
     : tensorAlu_io_acc_wr_0_bits_data_0_31; // @[Compute.scala 153:39]
  assign tensorGemm_clock = clock;
  assign tensorGemm_reset = reset;
  assign tensorGemm_io_start = tensorGemm_io_start_REG; // @[Compute.scala 162:23]
  assign tensorGemm_io_dec_wgt_1 = _tensorGemm_io_dec_WIRE_1[127:118]; // @[Compute.scala 163:51]
  assign tensorGemm_io_dec_wgt_0 = _tensorGemm_io_dec_WIRE_1[117:108]; // @[Compute.scala 163:51]
  assign tensorGemm_io_dec_inp_1 = _tensorGemm_io_dec_WIRE_1[107:97]; // @[Compute.scala 163:51]
  assign tensorGemm_io_dec_inp_0 = _tensorGemm_io_dec_WIRE_1[96:86]; // @[Compute.scala 163:51]
  assign tensorGemm_io_dec_acc_1 = _tensorGemm_io_dec_WIRE_1[85:75]; // @[Compute.scala 163:51]
  assign tensorGemm_io_dec_acc_0 = _tensorGemm_io_dec_WIRE_1[74:64]; // @[Compute.scala 163:51]
  assign tensorGemm_io_dec_empty_0 = _tensorGemm_io_dec_WIRE_1[63]; // @[Compute.scala 163:51]
  assign tensorGemm_io_dec_lp_1 = _tensorGemm_io_dec_WIRE_1[62:49]; // @[Compute.scala 163:51]
  assign tensorGemm_io_dec_lp_0 = _tensorGemm_io_dec_WIRE_1[48:35]; // @[Compute.scala 163:51]
  assign tensorGemm_io_dec_uop_end = _tensorGemm_io_dec_WIRE_1[34:21]; // @[Compute.scala 163:51]
  assign tensorGemm_io_dec_uop_begin = _tensorGemm_io_dec_WIRE_1[20:8]; // @[Compute.scala 163:51]
  assign tensorGemm_io_dec_reset = _tensorGemm_io_dec_WIRE_1[7]; // @[Compute.scala 163:51]
  assign tensorGemm_io_dec_push_next = _tensorGemm_io_dec_WIRE_1[6]; // @[Compute.scala 163:51]
  assign tensorGemm_io_dec_push_prev = _tensorGemm_io_dec_WIRE_1[5]; // @[Compute.scala 163:51]
  assign tensorGemm_io_dec_pop_next = _tensorGemm_io_dec_WIRE_1[4]; // @[Compute.scala 163:51]
  assign tensorGemm_io_dec_pop_prev = _tensorGemm_io_dec_WIRE_1[3]; // @[Compute.scala 163:51]
  assign tensorGemm_io_dec_op = _tensorGemm_io_dec_WIRE_1[2:0]; // @[Compute.scala 163:51]
  assign tensorGemm_io_uop_data_valid = loadUop_io_uop_data_valid & dec_io_isGemm; // @[Compute.scala 164:61]
  assign tensorGemm_io_uop_data_bits_u2 = loadUop_io_uop_data_bits_u2; // @[Compute.scala 165:31]
  assign tensorGemm_io_uop_data_bits_u1 = loadUop_io_uop_data_bits_u1; // @[Compute.scala 165:31]
  assign tensorGemm_io_uop_data_bits_u0 = loadUop_io_uop_data_bits_u0; // @[Compute.scala 165:31]
  assign tensorGemm_io_inp_rd_0_data_valid = io_inp_rd_0_data_valid; // @[Compute.scala 166:21]
  assign tensorGemm_io_inp_rd_0_data_bits_0_0 = io_inp_rd_0_data_bits_0_0; // @[Compute.scala 166:21]
  assign tensorGemm_io_inp_rd_0_data_bits_0_1 = io_inp_rd_0_data_bits_0_1; // @[Compute.scala 166:21]
  assign tensorGemm_io_inp_rd_0_data_bits_0_2 = io_inp_rd_0_data_bits_0_2; // @[Compute.scala 166:21]
  assign tensorGemm_io_inp_rd_0_data_bits_0_3 = io_inp_rd_0_data_bits_0_3; // @[Compute.scala 166:21]
  assign tensorGemm_io_inp_rd_0_data_bits_0_4 = io_inp_rd_0_data_bits_0_4; // @[Compute.scala 166:21]
  assign tensorGemm_io_inp_rd_0_data_bits_0_5 = io_inp_rd_0_data_bits_0_5; // @[Compute.scala 166:21]
  assign tensorGemm_io_inp_rd_0_data_bits_0_6 = io_inp_rd_0_data_bits_0_6; // @[Compute.scala 166:21]
  assign tensorGemm_io_inp_rd_0_data_bits_0_7 = io_inp_rd_0_data_bits_0_7; // @[Compute.scala 166:21]
  assign tensorGemm_io_inp_rd_0_data_bits_0_8 = io_inp_rd_0_data_bits_0_8; // @[Compute.scala 166:21]
  assign tensorGemm_io_inp_rd_0_data_bits_0_9 = io_inp_rd_0_data_bits_0_9; // @[Compute.scala 166:21]
  assign tensorGemm_io_inp_rd_0_data_bits_0_10 = io_inp_rd_0_data_bits_0_10; // @[Compute.scala 166:21]
  assign tensorGemm_io_inp_rd_0_data_bits_0_11 = io_inp_rd_0_data_bits_0_11; // @[Compute.scala 166:21]
  assign tensorGemm_io_inp_rd_0_data_bits_0_12 = io_inp_rd_0_data_bits_0_12; // @[Compute.scala 166:21]
  assign tensorGemm_io_inp_rd_0_data_bits_0_13 = io_inp_rd_0_data_bits_0_13; // @[Compute.scala 166:21]
  assign tensorGemm_io_inp_rd_0_data_bits_0_14 = io_inp_rd_0_data_bits_0_14; // @[Compute.scala 166:21]
  assign tensorGemm_io_inp_rd_0_data_bits_0_15 = io_inp_rd_0_data_bits_0_15; // @[Compute.scala 166:21]
  assign tensorGemm_io_wgt_rd_0_data_valid = io_wgt_rd_0_data_valid; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_0_0 = io_wgt_rd_0_data_bits_0_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_0_1 = io_wgt_rd_0_data_bits_0_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_0_2 = io_wgt_rd_0_data_bits_0_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_0_3 = io_wgt_rd_0_data_bits_0_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_0_4 = io_wgt_rd_0_data_bits_0_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_0_5 = io_wgt_rd_0_data_bits_0_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_0_6 = io_wgt_rd_0_data_bits_0_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_0_7 = io_wgt_rd_0_data_bits_0_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_0_8 = io_wgt_rd_0_data_bits_0_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_0_9 = io_wgt_rd_0_data_bits_0_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_0_10 = io_wgt_rd_0_data_bits_0_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_0_11 = io_wgt_rd_0_data_bits_0_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_0_12 = io_wgt_rd_0_data_bits_0_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_0_13 = io_wgt_rd_0_data_bits_0_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_0_14 = io_wgt_rd_0_data_bits_0_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_0_15 = io_wgt_rd_0_data_bits_0_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_1_0 = io_wgt_rd_0_data_bits_1_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_1_1 = io_wgt_rd_0_data_bits_1_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_1_2 = io_wgt_rd_0_data_bits_1_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_1_3 = io_wgt_rd_0_data_bits_1_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_1_4 = io_wgt_rd_0_data_bits_1_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_1_5 = io_wgt_rd_0_data_bits_1_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_1_6 = io_wgt_rd_0_data_bits_1_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_1_7 = io_wgt_rd_0_data_bits_1_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_1_8 = io_wgt_rd_0_data_bits_1_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_1_9 = io_wgt_rd_0_data_bits_1_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_1_10 = io_wgt_rd_0_data_bits_1_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_1_11 = io_wgt_rd_0_data_bits_1_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_1_12 = io_wgt_rd_0_data_bits_1_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_1_13 = io_wgt_rd_0_data_bits_1_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_1_14 = io_wgt_rd_0_data_bits_1_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_1_15 = io_wgt_rd_0_data_bits_1_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_2_0 = io_wgt_rd_0_data_bits_2_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_2_1 = io_wgt_rd_0_data_bits_2_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_2_2 = io_wgt_rd_0_data_bits_2_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_2_3 = io_wgt_rd_0_data_bits_2_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_2_4 = io_wgt_rd_0_data_bits_2_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_2_5 = io_wgt_rd_0_data_bits_2_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_2_6 = io_wgt_rd_0_data_bits_2_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_2_7 = io_wgt_rd_0_data_bits_2_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_2_8 = io_wgt_rd_0_data_bits_2_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_2_9 = io_wgt_rd_0_data_bits_2_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_2_10 = io_wgt_rd_0_data_bits_2_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_2_11 = io_wgt_rd_0_data_bits_2_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_2_12 = io_wgt_rd_0_data_bits_2_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_2_13 = io_wgt_rd_0_data_bits_2_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_2_14 = io_wgt_rd_0_data_bits_2_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_2_15 = io_wgt_rd_0_data_bits_2_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_3_0 = io_wgt_rd_0_data_bits_3_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_3_1 = io_wgt_rd_0_data_bits_3_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_3_2 = io_wgt_rd_0_data_bits_3_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_3_3 = io_wgt_rd_0_data_bits_3_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_3_4 = io_wgt_rd_0_data_bits_3_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_3_5 = io_wgt_rd_0_data_bits_3_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_3_6 = io_wgt_rd_0_data_bits_3_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_3_7 = io_wgt_rd_0_data_bits_3_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_3_8 = io_wgt_rd_0_data_bits_3_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_3_9 = io_wgt_rd_0_data_bits_3_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_3_10 = io_wgt_rd_0_data_bits_3_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_3_11 = io_wgt_rd_0_data_bits_3_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_3_12 = io_wgt_rd_0_data_bits_3_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_3_13 = io_wgt_rd_0_data_bits_3_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_3_14 = io_wgt_rd_0_data_bits_3_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_3_15 = io_wgt_rd_0_data_bits_3_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_4_0 = io_wgt_rd_0_data_bits_4_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_4_1 = io_wgt_rd_0_data_bits_4_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_4_2 = io_wgt_rd_0_data_bits_4_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_4_3 = io_wgt_rd_0_data_bits_4_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_4_4 = io_wgt_rd_0_data_bits_4_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_4_5 = io_wgt_rd_0_data_bits_4_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_4_6 = io_wgt_rd_0_data_bits_4_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_4_7 = io_wgt_rd_0_data_bits_4_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_4_8 = io_wgt_rd_0_data_bits_4_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_4_9 = io_wgt_rd_0_data_bits_4_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_4_10 = io_wgt_rd_0_data_bits_4_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_4_11 = io_wgt_rd_0_data_bits_4_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_4_12 = io_wgt_rd_0_data_bits_4_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_4_13 = io_wgt_rd_0_data_bits_4_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_4_14 = io_wgt_rd_0_data_bits_4_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_4_15 = io_wgt_rd_0_data_bits_4_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_5_0 = io_wgt_rd_0_data_bits_5_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_5_1 = io_wgt_rd_0_data_bits_5_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_5_2 = io_wgt_rd_0_data_bits_5_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_5_3 = io_wgt_rd_0_data_bits_5_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_5_4 = io_wgt_rd_0_data_bits_5_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_5_5 = io_wgt_rd_0_data_bits_5_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_5_6 = io_wgt_rd_0_data_bits_5_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_5_7 = io_wgt_rd_0_data_bits_5_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_5_8 = io_wgt_rd_0_data_bits_5_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_5_9 = io_wgt_rd_0_data_bits_5_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_5_10 = io_wgt_rd_0_data_bits_5_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_5_11 = io_wgt_rd_0_data_bits_5_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_5_12 = io_wgt_rd_0_data_bits_5_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_5_13 = io_wgt_rd_0_data_bits_5_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_5_14 = io_wgt_rd_0_data_bits_5_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_5_15 = io_wgt_rd_0_data_bits_5_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_6_0 = io_wgt_rd_0_data_bits_6_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_6_1 = io_wgt_rd_0_data_bits_6_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_6_2 = io_wgt_rd_0_data_bits_6_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_6_3 = io_wgt_rd_0_data_bits_6_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_6_4 = io_wgt_rd_0_data_bits_6_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_6_5 = io_wgt_rd_0_data_bits_6_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_6_6 = io_wgt_rd_0_data_bits_6_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_6_7 = io_wgt_rd_0_data_bits_6_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_6_8 = io_wgt_rd_0_data_bits_6_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_6_9 = io_wgt_rd_0_data_bits_6_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_6_10 = io_wgt_rd_0_data_bits_6_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_6_11 = io_wgt_rd_0_data_bits_6_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_6_12 = io_wgt_rd_0_data_bits_6_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_6_13 = io_wgt_rd_0_data_bits_6_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_6_14 = io_wgt_rd_0_data_bits_6_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_6_15 = io_wgt_rd_0_data_bits_6_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_7_0 = io_wgt_rd_0_data_bits_7_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_7_1 = io_wgt_rd_0_data_bits_7_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_7_2 = io_wgt_rd_0_data_bits_7_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_7_3 = io_wgt_rd_0_data_bits_7_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_7_4 = io_wgt_rd_0_data_bits_7_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_7_5 = io_wgt_rd_0_data_bits_7_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_7_6 = io_wgt_rd_0_data_bits_7_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_7_7 = io_wgt_rd_0_data_bits_7_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_7_8 = io_wgt_rd_0_data_bits_7_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_7_9 = io_wgt_rd_0_data_bits_7_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_7_10 = io_wgt_rd_0_data_bits_7_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_7_11 = io_wgt_rd_0_data_bits_7_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_7_12 = io_wgt_rd_0_data_bits_7_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_7_13 = io_wgt_rd_0_data_bits_7_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_7_14 = io_wgt_rd_0_data_bits_7_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_7_15 = io_wgt_rd_0_data_bits_7_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_8_0 = io_wgt_rd_0_data_bits_8_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_8_1 = io_wgt_rd_0_data_bits_8_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_8_2 = io_wgt_rd_0_data_bits_8_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_8_3 = io_wgt_rd_0_data_bits_8_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_8_4 = io_wgt_rd_0_data_bits_8_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_8_5 = io_wgt_rd_0_data_bits_8_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_8_6 = io_wgt_rd_0_data_bits_8_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_8_7 = io_wgt_rd_0_data_bits_8_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_8_8 = io_wgt_rd_0_data_bits_8_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_8_9 = io_wgt_rd_0_data_bits_8_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_8_10 = io_wgt_rd_0_data_bits_8_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_8_11 = io_wgt_rd_0_data_bits_8_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_8_12 = io_wgt_rd_0_data_bits_8_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_8_13 = io_wgt_rd_0_data_bits_8_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_8_14 = io_wgt_rd_0_data_bits_8_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_8_15 = io_wgt_rd_0_data_bits_8_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_9_0 = io_wgt_rd_0_data_bits_9_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_9_1 = io_wgt_rd_0_data_bits_9_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_9_2 = io_wgt_rd_0_data_bits_9_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_9_3 = io_wgt_rd_0_data_bits_9_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_9_4 = io_wgt_rd_0_data_bits_9_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_9_5 = io_wgt_rd_0_data_bits_9_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_9_6 = io_wgt_rd_0_data_bits_9_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_9_7 = io_wgt_rd_0_data_bits_9_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_9_8 = io_wgt_rd_0_data_bits_9_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_9_9 = io_wgt_rd_0_data_bits_9_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_9_10 = io_wgt_rd_0_data_bits_9_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_9_11 = io_wgt_rd_0_data_bits_9_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_9_12 = io_wgt_rd_0_data_bits_9_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_9_13 = io_wgt_rd_0_data_bits_9_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_9_14 = io_wgt_rd_0_data_bits_9_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_9_15 = io_wgt_rd_0_data_bits_9_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_10_0 = io_wgt_rd_0_data_bits_10_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_10_1 = io_wgt_rd_0_data_bits_10_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_10_2 = io_wgt_rd_0_data_bits_10_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_10_3 = io_wgt_rd_0_data_bits_10_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_10_4 = io_wgt_rd_0_data_bits_10_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_10_5 = io_wgt_rd_0_data_bits_10_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_10_6 = io_wgt_rd_0_data_bits_10_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_10_7 = io_wgt_rd_0_data_bits_10_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_10_8 = io_wgt_rd_0_data_bits_10_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_10_9 = io_wgt_rd_0_data_bits_10_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_10_10 = io_wgt_rd_0_data_bits_10_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_10_11 = io_wgt_rd_0_data_bits_10_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_10_12 = io_wgt_rd_0_data_bits_10_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_10_13 = io_wgt_rd_0_data_bits_10_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_10_14 = io_wgt_rd_0_data_bits_10_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_10_15 = io_wgt_rd_0_data_bits_10_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_11_0 = io_wgt_rd_0_data_bits_11_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_11_1 = io_wgt_rd_0_data_bits_11_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_11_2 = io_wgt_rd_0_data_bits_11_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_11_3 = io_wgt_rd_0_data_bits_11_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_11_4 = io_wgt_rd_0_data_bits_11_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_11_5 = io_wgt_rd_0_data_bits_11_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_11_6 = io_wgt_rd_0_data_bits_11_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_11_7 = io_wgt_rd_0_data_bits_11_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_11_8 = io_wgt_rd_0_data_bits_11_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_11_9 = io_wgt_rd_0_data_bits_11_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_11_10 = io_wgt_rd_0_data_bits_11_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_11_11 = io_wgt_rd_0_data_bits_11_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_11_12 = io_wgt_rd_0_data_bits_11_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_11_13 = io_wgt_rd_0_data_bits_11_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_11_14 = io_wgt_rd_0_data_bits_11_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_11_15 = io_wgt_rd_0_data_bits_11_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_12_0 = io_wgt_rd_0_data_bits_12_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_12_1 = io_wgt_rd_0_data_bits_12_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_12_2 = io_wgt_rd_0_data_bits_12_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_12_3 = io_wgt_rd_0_data_bits_12_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_12_4 = io_wgt_rd_0_data_bits_12_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_12_5 = io_wgt_rd_0_data_bits_12_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_12_6 = io_wgt_rd_0_data_bits_12_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_12_7 = io_wgt_rd_0_data_bits_12_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_12_8 = io_wgt_rd_0_data_bits_12_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_12_9 = io_wgt_rd_0_data_bits_12_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_12_10 = io_wgt_rd_0_data_bits_12_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_12_11 = io_wgt_rd_0_data_bits_12_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_12_12 = io_wgt_rd_0_data_bits_12_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_12_13 = io_wgt_rd_0_data_bits_12_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_12_14 = io_wgt_rd_0_data_bits_12_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_12_15 = io_wgt_rd_0_data_bits_12_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_13_0 = io_wgt_rd_0_data_bits_13_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_13_1 = io_wgt_rd_0_data_bits_13_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_13_2 = io_wgt_rd_0_data_bits_13_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_13_3 = io_wgt_rd_0_data_bits_13_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_13_4 = io_wgt_rd_0_data_bits_13_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_13_5 = io_wgt_rd_0_data_bits_13_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_13_6 = io_wgt_rd_0_data_bits_13_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_13_7 = io_wgt_rd_0_data_bits_13_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_13_8 = io_wgt_rd_0_data_bits_13_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_13_9 = io_wgt_rd_0_data_bits_13_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_13_10 = io_wgt_rd_0_data_bits_13_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_13_11 = io_wgt_rd_0_data_bits_13_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_13_12 = io_wgt_rd_0_data_bits_13_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_13_13 = io_wgt_rd_0_data_bits_13_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_13_14 = io_wgt_rd_0_data_bits_13_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_13_15 = io_wgt_rd_0_data_bits_13_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_14_0 = io_wgt_rd_0_data_bits_14_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_14_1 = io_wgt_rd_0_data_bits_14_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_14_2 = io_wgt_rd_0_data_bits_14_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_14_3 = io_wgt_rd_0_data_bits_14_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_14_4 = io_wgt_rd_0_data_bits_14_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_14_5 = io_wgt_rd_0_data_bits_14_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_14_6 = io_wgt_rd_0_data_bits_14_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_14_7 = io_wgt_rd_0_data_bits_14_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_14_8 = io_wgt_rd_0_data_bits_14_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_14_9 = io_wgt_rd_0_data_bits_14_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_14_10 = io_wgt_rd_0_data_bits_14_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_14_11 = io_wgt_rd_0_data_bits_14_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_14_12 = io_wgt_rd_0_data_bits_14_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_14_13 = io_wgt_rd_0_data_bits_14_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_14_14 = io_wgt_rd_0_data_bits_14_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_14_15 = io_wgt_rd_0_data_bits_14_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_15_0 = io_wgt_rd_0_data_bits_15_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_15_1 = io_wgt_rd_0_data_bits_15_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_15_2 = io_wgt_rd_0_data_bits_15_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_15_3 = io_wgt_rd_0_data_bits_15_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_15_4 = io_wgt_rd_0_data_bits_15_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_15_5 = io_wgt_rd_0_data_bits_15_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_15_6 = io_wgt_rd_0_data_bits_15_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_15_7 = io_wgt_rd_0_data_bits_15_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_15_8 = io_wgt_rd_0_data_bits_15_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_15_9 = io_wgt_rd_0_data_bits_15_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_15_10 = io_wgt_rd_0_data_bits_15_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_15_11 = io_wgt_rd_0_data_bits_15_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_15_12 = io_wgt_rd_0_data_bits_15_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_15_13 = io_wgt_rd_0_data_bits_15_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_15_14 = io_wgt_rd_0_data_bits_15_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_15_15 = io_wgt_rd_0_data_bits_15_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_16_0 = io_wgt_rd_0_data_bits_16_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_16_1 = io_wgt_rd_0_data_bits_16_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_16_2 = io_wgt_rd_0_data_bits_16_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_16_3 = io_wgt_rd_0_data_bits_16_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_16_4 = io_wgt_rd_0_data_bits_16_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_16_5 = io_wgt_rd_0_data_bits_16_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_16_6 = io_wgt_rd_0_data_bits_16_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_16_7 = io_wgt_rd_0_data_bits_16_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_16_8 = io_wgt_rd_0_data_bits_16_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_16_9 = io_wgt_rd_0_data_bits_16_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_16_10 = io_wgt_rd_0_data_bits_16_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_16_11 = io_wgt_rd_0_data_bits_16_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_16_12 = io_wgt_rd_0_data_bits_16_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_16_13 = io_wgt_rd_0_data_bits_16_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_16_14 = io_wgt_rd_0_data_bits_16_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_16_15 = io_wgt_rd_0_data_bits_16_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_17_0 = io_wgt_rd_0_data_bits_17_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_17_1 = io_wgt_rd_0_data_bits_17_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_17_2 = io_wgt_rd_0_data_bits_17_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_17_3 = io_wgt_rd_0_data_bits_17_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_17_4 = io_wgt_rd_0_data_bits_17_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_17_5 = io_wgt_rd_0_data_bits_17_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_17_6 = io_wgt_rd_0_data_bits_17_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_17_7 = io_wgt_rd_0_data_bits_17_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_17_8 = io_wgt_rd_0_data_bits_17_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_17_9 = io_wgt_rd_0_data_bits_17_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_17_10 = io_wgt_rd_0_data_bits_17_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_17_11 = io_wgt_rd_0_data_bits_17_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_17_12 = io_wgt_rd_0_data_bits_17_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_17_13 = io_wgt_rd_0_data_bits_17_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_17_14 = io_wgt_rd_0_data_bits_17_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_17_15 = io_wgt_rd_0_data_bits_17_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_18_0 = io_wgt_rd_0_data_bits_18_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_18_1 = io_wgt_rd_0_data_bits_18_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_18_2 = io_wgt_rd_0_data_bits_18_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_18_3 = io_wgt_rd_0_data_bits_18_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_18_4 = io_wgt_rd_0_data_bits_18_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_18_5 = io_wgt_rd_0_data_bits_18_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_18_6 = io_wgt_rd_0_data_bits_18_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_18_7 = io_wgt_rd_0_data_bits_18_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_18_8 = io_wgt_rd_0_data_bits_18_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_18_9 = io_wgt_rd_0_data_bits_18_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_18_10 = io_wgt_rd_0_data_bits_18_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_18_11 = io_wgt_rd_0_data_bits_18_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_18_12 = io_wgt_rd_0_data_bits_18_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_18_13 = io_wgt_rd_0_data_bits_18_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_18_14 = io_wgt_rd_0_data_bits_18_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_18_15 = io_wgt_rd_0_data_bits_18_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_19_0 = io_wgt_rd_0_data_bits_19_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_19_1 = io_wgt_rd_0_data_bits_19_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_19_2 = io_wgt_rd_0_data_bits_19_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_19_3 = io_wgt_rd_0_data_bits_19_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_19_4 = io_wgt_rd_0_data_bits_19_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_19_5 = io_wgt_rd_0_data_bits_19_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_19_6 = io_wgt_rd_0_data_bits_19_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_19_7 = io_wgt_rd_0_data_bits_19_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_19_8 = io_wgt_rd_0_data_bits_19_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_19_9 = io_wgt_rd_0_data_bits_19_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_19_10 = io_wgt_rd_0_data_bits_19_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_19_11 = io_wgt_rd_0_data_bits_19_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_19_12 = io_wgt_rd_0_data_bits_19_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_19_13 = io_wgt_rd_0_data_bits_19_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_19_14 = io_wgt_rd_0_data_bits_19_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_19_15 = io_wgt_rd_0_data_bits_19_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_20_0 = io_wgt_rd_0_data_bits_20_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_20_1 = io_wgt_rd_0_data_bits_20_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_20_2 = io_wgt_rd_0_data_bits_20_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_20_3 = io_wgt_rd_0_data_bits_20_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_20_4 = io_wgt_rd_0_data_bits_20_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_20_5 = io_wgt_rd_0_data_bits_20_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_20_6 = io_wgt_rd_0_data_bits_20_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_20_7 = io_wgt_rd_0_data_bits_20_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_20_8 = io_wgt_rd_0_data_bits_20_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_20_9 = io_wgt_rd_0_data_bits_20_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_20_10 = io_wgt_rd_0_data_bits_20_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_20_11 = io_wgt_rd_0_data_bits_20_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_20_12 = io_wgt_rd_0_data_bits_20_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_20_13 = io_wgt_rd_0_data_bits_20_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_20_14 = io_wgt_rd_0_data_bits_20_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_20_15 = io_wgt_rd_0_data_bits_20_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_21_0 = io_wgt_rd_0_data_bits_21_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_21_1 = io_wgt_rd_0_data_bits_21_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_21_2 = io_wgt_rd_0_data_bits_21_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_21_3 = io_wgt_rd_0_data_bits_21_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_21_4 = io_wgt_rd_0_data_bits_21_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_21_5 = io_wgt_rd_0_data_bits_21_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_21_6 = io_wgt_rd_0_data_bits_21_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_21_7 = io_wgt_rd_0_data_bits_21_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_21_8 = io_wgt_rd_0_data_bits_21_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_21_9 = io_wgt_rd_0_data_bits_21_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_21_10 = io_wgt_rd_0_data_bits_21_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_21_11 = io_wgt_rd_0_data_bits_21_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_21_12 = io_wgt_rd_0_data_bits_21_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_21_13 = io_wgt_rd_0_data_bits_21_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_21_14 = io_wgt_rd_0_data_bits_21_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_21_15 = io_wgt_rd_0_data_bits_21_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_22_0 = io_wgt_rd_0_data_bits_22_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_22_1 = io_wgt_rd_0_data_bits_22_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_22_2 = io_wgt_rd_0_data_bits_22_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_22_3 = io_wgt_rd_0_data_bits_22_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_22_4 = io_wgt_rd_0_data_bits_22_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_22_5 = io_wgt_rd_0_data_bits_22_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_22_6 = io_wgt_rd_0_data_bits_22_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_22_7 = io_wgt_rd_0_data_bits_22_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_22_8 = io_wgt_rd_0_data_bits_22_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_22_9 = io_wgt_rd_0_data_bits_22_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_22_10 = io_wgt_rd_0_data_bits_22_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_22_11 = io_wgt_rd_0_data_bits_22_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_22_12 = io_wgt_rd_0_data_bits_22_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_22_13 = io_wgt_rd_0_data_bits_22_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_22_14 = io_wgt_rd_0_data_bits_22_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_22_15 = io_wgt_rd_0_data_bits_22_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_23_0 = io_wgt_rd_0_data_bits_23_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_23_1 = io_wgt_rd_0_data_bits_23_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_23_2 = io_wgt_rd_0_data_bits_23_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_23_3 = io_wgt_rd_0_data_bits_23_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_23_4 = io_wgt_rd_0_data_bits_23_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_23_5 = io_wgt_rd_0_data_bits_23_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_23_6 = io_wgt_rd_0_data_bits_23_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_23_7 = io_wgt_rd_0_data_bits_23_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_23_8 = io_wgt_rd_0_data_bits_23_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_23_9 = io_wgt_rd_0_data_bits_23_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_23_10 = io_wgt_rd_0_data_bits_23_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_23_11 = io_wgt_rd_0_data_bits_23_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_23_12 = io_wgt_rd_0_data_bits_23_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_23_13 = io_wgt_rd_0_data_bits_23_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_23_14 = io_wgt_rd_0_data_bits_23_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_23_15 = io_wgt_rd_0_data_bits_23_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_24_0 = io_wgt_rd_0_data_bits_24_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_24_1 = io_wgt_rd_0_data_bits_24_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_24_2 = io_wgt_rd_0_data_bits_24_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_24_3 = io_wgt_rd_0_data_bits_24_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_24_4 = io_wgt_rd_0_data_bits_24_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_24_5 = io_wgt_rd_0_data_bits_24_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_24_6 = io_wgt_rd_0_data_bits_24_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_24_7 = io_wgt_rd_0_data_bits_24_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_24_8 = io_wgt_rd_0_data_bits_24_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_24_9 = io_wgt_rd_0_data_bits_24_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_24_10 = io_wgt_rd_0_data_bits_24_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_24_11 = io_wgt_rd_0_data_bits_24_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_24_12 = io_wgt_rd_0_data_bits_24_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_24_13 = io_wgt_rd_0_data_bits_24_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_24_14 = io_wgt_rd_0_data_bits_24_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_24_15 = io_wgt_rd_0_data_bits_24_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_25_0 = io_wgt_rd_0_data_bits_25_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_25_1 = io_wgt_rd_0_data_bits_25_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_25_2 = io_wgt_rd_0_data_bits_25_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_25_3 = io_wgt_rd_0_data_bits_25_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_25_4 = io_wgt_rd_0_data_bits_25_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_25_5 = io_wgt_rd_0_data_bits_25_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_25_6 = io_wgt_rd_0_data_bits_25_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_25_7 = io_wgt_rd_0_data_bits_25_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_25_8 = io_wgt_rd_0_data_bits_25_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_25_9 = io_wgt_rd_0_data_bits_25_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_25_10 = io_wgt_rd_0_data_bits_25_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_25_11 = io_wgt_rd_0_data_bits_25_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_25_12 = io_wgt_rd_0_data_bits_25_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_25_13 = io_wgt_rd_0_data_bits_25_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_25_14 = io_wgt_rd_0_data_bits_25_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_25_15 = io_wgt_rd_0_data_bits_25_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_26_0 = io_wgt_rd_0_data_bits_26_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_26_1 = io_wgt_rd_0_data_bits_26_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_26_2 = io_wgt_rd_0_data_bits_26_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_26_3 = io_wgt_rd_0_data_bits_26_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_26_4 = io_wgt_rd_0_data_bits_26_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_26_5 = io_wgt_rd_0_data_bits_26_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_26_6 = io_wgt_rd_0_data_bits_26_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_26_7 = io_wgt_rd_0_data_bits_26_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_26_8 = io_wgt_rd_0_data_bits_26_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_26_9 = io_wgt_rd_0_data_bits_26_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_26_10 = io_wgt_rd_0_data_bits_26_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_26_11 = io_wgt_rd_0_data_bits_26_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_26_12 = io_wgt_rd_0_data_bits_26_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_26_13 = io_wgt_rd_0_data_bits_26_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_26_14 = io_wgt_rd_0_data_bits_26_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_26_15 = io_wgt_rd_0_data_bits_26_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_27_0 = io_wgt_rd_0_data_bits_27_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_27_1 = io_wgt_rd_0_data_bits_27_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_27_2 = io_wgt_rd_0_data_bits_27_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_27_3 = io_wgt_rd_0_data_bits_27_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_27_4 = io_wgt_rd_0_data_bits_27_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_27_5 = io_wgt_rd_0_data_bits_27_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_27_6 = io_wgt_rd_0_data_bits_27_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_27_7 = io_wgt_rd_0_data_bits_27_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_27_8 = io_wgt_rd_0_data_bits_27_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_27_9 = io_wgt_rd_0_data_bits_27_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_27_10 = io_wgt_rd_0_data_bits_27_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_27_11 = io_wgt_rd_0_data_bits_27_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_27_12 = io_wgt_rd_0_data_bits_27_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_27_13 = io_wgt_rd_0_data_bits_27_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_27_14 = io_wgt_rd_0_data_bits_27_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_27_15 = io_wgt_rd_0_data_bits_27_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_28_0 = io_wgt_rd_0_data_bits_28_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_28_1 = io_wgt_rd_0_data_bits_28_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_28_2 = io_wgt_rd_0_data_bits_28_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_28_3 = io_wgt_rd_0_data_bits_28_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_28_4 = io_wgt_rd_0_data_bits_28_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_28_5 = io_wgt_rd_0_data_bits_28_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_28_6 = io_wgt_rd_0_data_bits_28_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_28_7 = io_wgt_rd_0_data_bits_28_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_28_8 = io_wgt_rd_0_data_bits_28_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_28_9 = io_wgt_rd_0_data_bits_28_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_28_10 = io_wgt_rd_0_data_bits_28_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_28_11 = io_wgt_rd_0_data_bits_28_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_28_12 = io_wgt_rd_0_data_bits_28_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_28_13 = io_wgt_rd_0_data_bits_28_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_28_14 = io_wgt_rd_0_data_bits_28_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_28_15 = io_wgt_rd_0_data_bits_28_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_29_0 = io_wgt_rd_0_data_bits_29_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_29_1 = io_wgt_rd_0_data_bits_29_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_29_2 = io_wgt_rd_0_data_bits_29_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_29_3 = io_wgt_rd_0_data_bits_29_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_29_4 = io_wgt_rd_0_data_bits_29_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_29_5 = io_wgt_rd_0_data_bits_29_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_29_6 = io_wgt_rd_0_data_bits_29_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_29_7 = io_wgt_rd_0_data_bits_29_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_29_8 = io_wgt_rd_0_data_bits_29_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_29_9 = io_wgt_rd_0_data_bits_29_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_29_10 = io_wgt_rd_0_data_bits_29_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_29_11 = io_wgt_rd_0_data_bits_29_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_29_12 = io_wgt_rd_0_data_bits_29_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_29_13 = io_wgt_rd_0_data_bits_29_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_29_14 = io_wgt_rd_0_data_bits_29_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_29_15 = io_wgt_rd_0_data_bits_29_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_30_0 = io_wgt_rd_0_data_bits_30_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_30_1 = io_wgt_rd_0_data_bits_30_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_30_2 = io_wgt_rd_0_data_bits_30_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_30_3 = io_wgt_rd_0_data_bits_30_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_30_4 = io_wgt_rd_0_data_bits_30_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_30_5 = io_wgt_rd_0_data_bits_30_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_30_6 = io_wgt_rd_0_data_bits_30_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_30_7 = io_wgt_rd_0_data_bits_30_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_30_8 = io_wgt_rd_0_data_bits_30_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_30_9 = io_wgt_rd_0_data_bits_30_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_30_10 = io_wgt_rd_0_data_bits_30_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_30_11 = io_wgt_rd_0_data_bits_30_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_30_12 = io_wgt_rd_0_data_bits_30_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_30_13 = io_wgt_rd_0_data_bits_30_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_30_14 = io_wgt_rd_0_data_bits_30_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_30_15 = io_wgt_rd_0_data_bits_30_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_31_0 = io_wgt_rd_0_data_bits_31_0; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_31_1 = io_wgt_rd_0_data_bits_31_1; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_31_2 = io_wgt_rd_0_data_bits_31_2; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_31_3 = io_wgt_rd_0_data_bits_31_3; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_31_4 = io_wgt_rd_0_data_bits_31_4; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_31_5 = io_wgt_rd_0_data_bits_31_5; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_31_6 = io_wgt_rd_0_data_bits_31_6; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_31_7 = io_wgt_rd_0_data_bits_31_7; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_31_8 = io_wgt_rd_0_data_bits_31_8; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_31_9 = io_wgt_rd_0_data_bits_31_9; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_31_10 = io_wgt_rd_0_data_bits_31_10; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_31_11 = io_wgt_rd_0_data_bits_31_11; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_31_12 = io_wgt_rd_0_data_bits_31_12; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_31_13 = io_wgt_rd_0_data_bits_31_13; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_31_14 = io_wgt_rd_0_data_bits_31_14; // @[Compute.scala 167:21]
  assign tensorGemm_io_wgt_rd_0_data_bits_31_15 = io_wgt_rd_0_data_bits_31_15; // @[Compute.scala 167:21]
  assign tensorGemm_io_acc_rd_0_data_valid = tensorAcc_io_tensor_rd_0_data_valid & tensorGemm_io_acc_rd_0_data_valid_REG
    ; // @[Compute.scala 170:46]
  assign tensorGemm_io_acc_rd_0_data_bits_0_0 = tensorAcc_io_tensor_rd_0_data_bits_0_0; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_1 = tensorAcc_io_tensor_rd_0_data_bits_0_1; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_2 = tensorAcc_io_tensor_rd_0_data_bits_0_2; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_3 = tensorAcc_io_tensor_rd_0_data_bits_0_3; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_4 = tensorAcc_io_tensor_rd_0_data_bits_0_4; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_5 = tensorAcc_io_tensor_rd_0_data_bits_0_5; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_6 = tensorAcc_io_tensor_rd_0_data_bits_0_6; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_7 = tensorAcc_io_tensor_rd_0_data_bits_0_7; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_8 = tensorAcc_io_tensor_rd_0_data_bits_0_8; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_9 = tensorAcc_io_tensor_rd_0_data_bits_0_9; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_10 = tensorAcc_io_tensor_rd_0_data_bits_0_10; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_11 = tensorAcc_io_tensor_rd_0_data_bits_0_11; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_12 = tensorAcc_io_tensor_rd_0_data_bits_0_12; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_13 = tensorAcc_io_tensor_rd_0_data_bits_0_13; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_14 = tensorAcc_io_tensor_rd_0_data_bits_0_14; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_15 = tensorAcc_io_tensor_rd_0_data_bits_0_15; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_16 = tensorAcc_io_tensor_rd_0_data_bits_0_16; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_17 = tensorAcc_io_tensor_rd_0_data_bits_0_17; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_18 = tensorAcc_io_tensor_rd_0_data_bits_0_18; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_19 = tensorAcc_io_tensor_rd_0_data_bits_0_19; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_20 = tensorAcc_io_tensor_rd_0_data_bits_0_20; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_21 = tensorAcc_io_tensor_rd_0_data_bits_0_21; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_22 = tensorAcc_io_tensor_rd_0_data_bits_0_22; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_23 = tensorAcc_io_tensor_rd_0_data_bits_0_23; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_24 = tensorAcc_io_tensor_rd_0_data_bits_0_24; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_25 = tensorAcc_io_tensor_rd_0_data_bits_0_25; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_26 = tensorAcc_io_tensor_rd_0_data_bits_0_26; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_27 = tensorAcc_io_tensor_rd_0_data_bits_0_27; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_28 = tensorAcc_io_tensor_rd_0_data_bits_0_28; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_29 = tensorAcc_io_tensor_rd_0_data_bits_0_29; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_30 = tensorAcc_io_tensor_rd_0_data_bits_0_30; // @[Compute.scala 171:41]
  assign tensorGemm_io_acc_rd_0_data_bits_0_31 = tensorAcc_io_tensor_rd_0_data_bits_0_31; // @[Compute.scala 171:41]
  assign tensorGemm_io_out_rd_0_data_valid = 1'h0; // @[Compute.scala 175:33]
  assign tensorAlu_clock = clock;
  assign tensorAlu_reset = reset;
  assign tensorAlu_io_start = tensorAlu_io_start_REG; // @[Compute.scala 180:22]
  assign tensorAlu_io_dec_alu_imm = _tensorGemm_io_dec_WIRE_1[127:112]; // @[Compute.scala 181:50]
  assign tensorAlu_io_dec_alu_use_imm = _tensorGemm_io_dec_WIRE_1[111]; // @[Compute.scala 181:50]
  assign tensorAlu_io_dec_alu_op = _tensorGemm_io_dec_WIRE_1[110:108]; // @[Compute.scala 181:50]
  assign tensorAlu_io_dec_src_1 = _tensorGemm_io_dec_WIRE_1[107:97]; // @[Compute.scala 181:50]
  assign tensorAlu_io_dec_src_0 = _tensorGemm_io_dec_WIRE_1[96:86]; // @[Compute.scala 181:50]
  assign tensorAlu_io_dec_dst_1 = _tensorGemm_io_dec_WIRE_1[85:75]; // @[Compute.scala 181:50]
  assign tensorAlu_io_dec_dst_0 = _tensorGemm_io_dec_WIRE_1[74:64]; // @[Compute.scala 181:50]
  assign tensorAlu_io_dec_lp_1 = _tensorGemm_io_dec_WIRE_1[62:49]; // @[Compute.scala 181:50]
  assign tensorAlu_io_dec_lp_0 = _tensorGemm_io_dec_WIRE_1[48:35]; // @[Compute.scala 181:50]
  assign tensorAlu_io_dec_uop_end = _tensorGemm_io_dec_WIRE_1[34:21]; // @[Compute.scala 181:50]
  assign tensorAlu_io_dec_uop_begin = _tensorGemm_io_dec_WIRE_1[20:8]; // @[Compute.scala 181:50]
  assign tensorAlu_io_uop_data_bits_u2 = loadUop_io_uop_data_bits_u2; // @[Compute.scala 183:30]
  assign tensorAlu_io_uop_data_bits_u1 = loadUop_io_uop_data_bits_u1; // @[Compute.scala 183:30]
  assign tensorAlu_io_uop_data_bits_u0 = loadUop_io_uop_data_bits_u0; // @[Compute.scala 183:30]
  assign tensorAlu_io_acc_rd_0_data_valid = tensorAcc_io_tensor_rd_0_data_valid & tensorAlu_io_acc_rd_0_data_valid_REG; // @[Compute.scala 186:46]
  assign tensorAlu_io_acc_rd_0_data_bits_0_0 = tensorAcc_io_tensor_rd_0_data_bits_0_0; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_1 = tensorAcc_io_tensor_rd_0_data_bits_0_1; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_2 = tensorAcc_io_tensor_rd_0_data_bits_0_2; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_3 = tensorAcc_io_tensor_rd_0_data_bits_0_3; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_4 = tensorAcc_io_tensor_rd_0_data_bits_0_4; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_5 = tensorAcc_io_tensor_rd_0_data_bits_0_5; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_6 = tensorAcc_io_tensor_rd_0_data_bits_0_6; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_7 = tensorAcc_io_tensor_rd_0_data_bits_0_7; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_8 = tensorAcc_io_tensor_rd_0_data_bits_0_8; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_9 = tensorAcc_io_tensor_rd_0_data_bits_0_9; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_10 = tensorAcc_io_tensor_rd_0_data_bits_0_10; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_11 = tensorAcc_io_tensor_rd_0_data_bits_0_11; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_12 = tensorAcc_io_tensor_rd_0_data_bits_0_12; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_13 = tensorAcc_io_tensor_rd_0_data_bits_0_13; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_14 = tensorAcc_io_tensor_rd_0_data_bits_0_14; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_15 = tensorAcc_io_tensor_rd_0_data_bits_0_15; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_16 = tensorAcc_io_tensor_rd_0_data_bits_0_16; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_17 = tensorAcc_io_tensor_rd_0_data_bits_0_17; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_18 = tensorAcc_io_tensor_rd_0_data_bits_0_18; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_19 = tensorAcc_io_tensor_rd_0_data_bits_0_19; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_20 = tensorAcc_io_tensor_rd_0_data_bits_0_20; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_21 = tensorAcc_io_tensor_rd_0_data_bits_0_21; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_22 = tensorAcc_io_tensor_rd_0_data_bits_0_22; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_23 = tensorAcc_io_tensor_rd_0_data_bits_0_23; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_24 = tensorAcc_io_tensor_rd_0_data_bits_0_24; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_25 = tensorAcc_io_tensor_rd_0_data_bits_0_25; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_26 = tensorAcc_io_tensor_rd_0_data_bits_0_26; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_27 = tensorAcc_io_tensor_rd_0_data_bits_0_27; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_28 = tensorAcc_io_tensor_rd_0_data_bits_0_28; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_29 = tensorAcc_io_tensor_rd_0_data_bits_0_29; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_30 = tensorAcc_io_tensor_rd_0_data_bits_0_30; // @[Compute.scala 187:40]
  assign tensorAlu_io_acc_rd_0_data_bits_0_31 = tensorAcc_io_tensor_rd_0_data_bits_0_31; // @[Compute.scala 187:40]
  assign tensorAlu_io_out_rd_0_data_valid = 1'h0; // @[Compute.scala 191:33]
  assign inst_q_clock = clock;
  assign inst_q_reset = reset;
  assign inst_q_io_enq_valid = io_inst_valid; // @[Compute.scala 120:17]
  assign inst_q_io_enq_bits = io_inst_bits; // @[Compute.scala 120:17]
  assign inst_q_io_deq_ready = state == 2'h2 & done | state == 2'h1; // @[Compute.scala 121:50]
  assign dec_io_inst = inst_q_io_deq_bits; // @[Compute.scala 73:15]
  always @(posedge clock) begin
    if (reset) begin // @[Compute.scala 55:22]
      state <= 2'h0; // @[Compute.scala 55:22]
    end else if (2'h0 == state) begin // @[Compute.scala 99:17]
      if (start) begin // @[Compute.scala 101:19]
        if (dec_io_isSync) begin // @[Compute.scala 102:29]
          state <= 2'h1; // @[Compute.scala 103:17]
        end else begin
          state <= _GEN_0;
        end
      end
    end else if (2'h1 == state) begin // @[Compute.scala 99:17]
      state <= 2'h0; // @[Compute.scala 110:13]
    end else if (2'h2 == state) begin // @[Compute.scala 99:17]
      state <= _GEN_3;
    end
    if (reset) begin // @[Compute.scala 150:14]
      tensorAcc_io_tensor_rd_0_idx_REG <= 1'h0; // @[Compute.scala 150:14]
    end else begin
      tensorAcc_io_tensor_rd_0_idx_REG <= dec_io_isGemm; // @[Compute.scala 150:14]
    end
    if (reset) begin // @[Compute.scala 154:14]
      tensorAcc_io_tensor_wr_0_REG <= 1'h0; // @[Compute.scala 154:14]
    end else begin
      tensorAcc_io_tensor_wr_0_REG <= dec_io_isGemm; // @[Compute.scala 154:14]
    end
    if (reset) begin // @[Compute.scala 162:33]
      tensorGemm_io_start_REG <= 1'h0; // @[Compute.scala 162:33]
    end else begin
      tensorGemm_io_start_REG <= _loadUop_io_start_T_1 & dec_io_isGemm; // @[Compute.scala 162:33]
    end
    if (reset) begin // @[Compute.scala 170:55]
      tensorGemm_io_acc_rd_0_data_valid_REG <= 1'h0; // @[Compute.scala 170:55]
    end else begin
      tensorGemm_io_acc_rd_0_data_valid_REG <= dec_io_isGemm; // @[Compute.scala 170:55]
    end
    if (reset) begin // @[Compute.scala 180:32]
      tensorAlu_io_start_REG <= 1'h0; // @[Compute.scala 180:32]
    end else begin
      tensorAlu_io_start_REG <= _loadUop_io_start_T_1 & dec_io_isAlu; // @[Compute.scala 180:32]
    end
    if (reset) begin // @[Compute.scala 186:55]
      tensorAlu_io_acc_rd_0_data_valid_REG <= 1'h0; // @[Compute.scala 186:55]
    end else begin
      tensorAlu_io_acc_rd_0_data_valid_REG <= dec_io_isAlu; // @[Compute.scala 186:55]
    end
    if (reset) begin // @[Compute.scala 208:12]
      io_out_wr_0_valid_REG <= 1'h0; // @[Compute.scala 208:12]
    end else begin
      io_out_wr_0_valid_REG <= dec_io_isGemm; // @[Compute.scala 208:12]
    end
    if (reset) begin // @[Compute.scala 210:12]
      io_out_wr_0_bits_idx_REG <= 1'h0; // @[Compute.scala 210:12]
    end else begin
      io_out_wr_0_bits_idx_REG <= dec_io_isGemm; // @[Compute.scala 210:12]
    end
    if (reset) begin // @[Compute.scala 221:14]
      outDataBits_0_REG <= 1'h0; // @[Compute.scala 221:14]
    end else begin
      outDataBits_0_REG <= dec_io_isGemm; // @[Compute.scala 221:14]
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~reset & ~(~tensorGemm_io_uop_idx_valid | ~tensorAlu_io_uop_idx_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Compute.scala:129 assert(!tensorGemm.io.uop.idx.valid || !tensorAlu.io.uop.idx.valid)\n"
            ); // @[Compute.scala 129:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(~tensorGemm_io_out_rd_0_data_valid | ~tensorAlu_io_out_rd_0_data_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Compute.scala:201 assert(!tensorGemm.io.out.rd(idx).data.valid || !tensorAlu.io.out.rd(idx).data.valid)\n"
            ); // @[Compute.scala 201:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_8 & ~(~tensorGemm_io_out_wr_0_valid | ~tensorAlu_io_out_wr_0_valid)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at Compute.scala:203 assert(!tensorGemm.io.out.wr(idx).valid || !tensorAlu.io.out.wr(idx).valid)\n"
            ); // @[Compute.scala 203:11]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  tensorAcc_io_tensor_rd_0_idx_REG = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  tensorAcc_io_tensor_wr_0_REG = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  tensorGemm_io_start_REG = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  tensorGemm_io_acc_rd_0_data_valid_REG = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  tensorAlu_io_start_REG = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  tensorAlu_io_acc_rd_0_data_valid_REG = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  io_out_wr_0_valid_REG = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  io_out_wr_0_bits_idx_REG = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  outDataBits_0_REG = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (~reset) begin
      assert(~tensorGemm_io_uop_idx_valid | ~tensorAlu_io_uop_idx_valid); // @[Compute.scala 129:9]
    end
    //
    if (_T_8) begin
      assert(1'h1); // @[Compute.scala 200:11]
    end
    //
    if (_T_8) begin
      assert(~tensorGemm_io_out_rd_0_data_valid | ~tensorAlu_io_out_rd_0_data_valid); // @[Compute.scala 201:11]
    end
    //
    if (_T_8) begin
      assert(~tensorGemm_io_out_wr_0_valid | ~tensorAlu_io_out_wr_0_valid); // @[Compute.scala 203:11]
    end
  end
endmodule
module StoreDecode(
  input  [127:0] io_inst,
  output         io_push_prev,
  output         io_pop_prev,
  output         io_isStore,
  output         io_isSync
);
  wire [15:0] dec_xsize = io_inst[95:80]; // @[Decode.scala 224:29]
  wire [127:0] _io_isStore_T = io_inst & 128'h7; // @[Decode.scala 227:25]
  wire  _io_isStore_T_1 = 128'h1 == _io_isStore_T; // @[Decode.scala 227:25]
  assign io_push_prev = io_inst[5]; // @[Decode.scala 224:29]
  assign io_pop_prev = io_inst[3]; // @[Decode.scala 224:29]
  assign io_isStore = 128'h1 == _io_isStore_T & dec_xsize != 16'h0; // @[Decode.scala 227:34]
  assign io_isSync = _io_isStore_T_1 & dec_xsize == 16'h0; // @[Decode.scala 228:33]
endmodule
module TensorStoreNarrowVME(
  input          clock,
  input          reset,
  input          io_start,
  output         io_done,
  input  [127:0] io_inst,
  input  [31:0]  io_baddr,
  input          io_vme_wr_cmd_ready,
  output         io_vme_wr_cmd_valid,
  output [31:0]  io_vme_wr_cmd_bits_addr,
  output [3:0]   io_vme_wr_cmd_bits_len,
  input          io_vme_wr_data_ready,
  output         io_vme_wr_data_valid,
  output [63:0]  io_vme_wr_data_bits_data,
  input          io_vme_wr_ack,
  input          io_tensor_wr_0_valid,
  input  [6:0]   io_tensor_wr_0_bits_idx,
  input  [7:0]   io_tensor_wr_0_bits_data_0_0,
  input  [7:0]   io_tensor_wr_0_bits_data_0_1,
  input  [7:0]   io_tensor_wr_0_bits_data_0_2,
  input  [7:0]   io_tensor_wr_0_bits_data_0_3,
  input  [7:0]   io_tensor_wr_0_bits_data_0_4,
  input  [7:0]   io_tensor_wr_0_bits_data_0_5,
  input  [7:0]   io_tensor_wr_0_bits_data_0_6,
  input  [7:0]   io_tensor_wr_0_bits_data_0_7,
  input  [7:0]   io_tensor_wr_0_bits_data_0_8,
  input  [7:0]   io_tensor_wr_0_bits_data_0_9,
  input  [7:0]   io_tensor_wr_0_bits_data_0_10,
  input  [7:0]   io_tensor_wr_0_bits_data_0_11,
  input  [7:0]   io_tensor_wr_0_bits_data_0_12,
  input  [7:0]   io_tensor_wr_0_bits_data_0_13,
  input  [7:0]   io_tensor_wr_0_bits_data_0_14,
  input  [7:0]   io_tensor_wr_0_bits_data_0_15,
  input  [7:0]   io_tensor_wr_0_bits_data_0_16,
  input  [7:0]   io_tensor_wr_0_bits_data_0_17,
  input  [7:0]   io_tensor_wr_0_bits_data_0_18,
  input  [7:0]   io_tensor_wr_0_bits_data_0_19,
  input  [7:0]   io_tensor_wr_0_bits_data_0_20,
  input  [7:0]   io_tensor_wr_0_bits_data_0_21,
  input  [7:0]   io_tensor_wr_0_bits_data_0_22,
  input  [7:0]   io_tensor_wr_0_bits_data_0_23,
  input  [7:0]   io_tensor_wr_0_bits_data_0_24,
  input  [7:0]   io_tensor_wr_0_bits_data_0_25,
  input  [7:0]   io_tensor_wr_0_bits_data_0_26,
  input  [7:0]   io_tensor_wr_0_bits_data_0_27,
  input  [7:0]   io_tensor_wr_0_bits_data_0_28,
  input  [7:0]   io_tensor_wr_0_bits_data_0_29,
  input  [7:0]   io_tensor_wr_0_bits_data_0_30,
  input  [7:0]   io_tensor_wr_0_bits_data_0_31
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] tensorFile_0_0 [0:127]; // @[TensorStoreNarrowVME.scala 167:16]
  wire  tensorFile_0_0_MPORT_1_en; // @[TensorStoreNarrowVME.scala 167:16]
  wire [6:0] tensorFile_0_0_MPORT_1_addr; // @[TensorStoreNarrowVME.scala 167:16]
  wire [63:0] tensorFile_0_0_MPORT_1_data; // @[TensorStoreNarrowVME.scala 167:16]
  wire [63:0] tensorFile_0_0_MPORT_data; // @[TensorStoreNarrowVME.scala 167:16]
  wire [6:0] tensorFile_0_0_MPORT_addr; // @[TensorStoreNarrowVME.scala 167:16]
  wire  tensorFile_0_0_MPORT_mask; // @[TensorStoreNarrowVME.scala 167:16]
  wire  tensorFile_0_0_MPORT_en; // @[TensorStoreNarrowVME.scala 167:16]
  reg  tensorFile_0_0_MPORT_1_en_pipe_0;
  reg [6:0] tensorFile_0_0_MPORT_1_addr_pipe_0;
  reg [63:0] tensorFile_0_1 [0:127]; // @[TensorStoreNarrowVME.scala 167:16]
  wire  tensorFile_0_1_MPORT_1_en; // @[TensorStoreNarrowVME.scala 167:16]
  wire [6:0] tensorFile_0_1_MPORT_1_addr; // @[TensorStoreNarrowVME.scala 167:16]
  wire [63:0] tensorFile_0_1_MPORT_1_data; // @[TensorStoreNarrowVME.scala 167:16]
  wire [63:0] tensorFile_0_1_MPORT_data; // @[TensorStoreNarrowVME.scala 167:16]
  wire [6:0] tensorFile_0_1_MPORT_addr; // @[TensorStoreNarrowVME.scala 167:16]
  wire  tensorFile_0_1_MPORT_mask; // @[TensorStoreNarrowVME.scala 167:16]
  wire  tensorFile_0_1_MPORT_en; // @[TensorStoreNarrowVME.scala 167:16]
  reg  tensorFile_0_1_MPORT_1_en_pipe_0;
  reg [6:0] tensorFile_0_1_MPORT_1_addr_pipe_0;
  reg [63:0] tensorFile_0_2 [0:127]; // @[TensorStoreNarrowVME.scala 167:16]
  wire  tensorFile_0_2_MPORT_1_en; // @[TensorStoreNarrowVME.scala 167:16]
  wire [6:0] tensorFile_0_2_MPORT_1_addr; // @[TensorStoreNarrowVME.scala 167:16]
  wire [63:0] tensorFile_0_2_MPORT_1_data; // @[TensorStoreNarrowVME.scala 167:16]
  wire [63:0] tensorFile_0_2_MPORT_data; // @[TensorStoreNarrowVME.scala 167:16]
  wire [6:0] tensorFile_0_2_MPORT_addr; // @[TensorStoreNarrowVME.scala 167:16]
  wire  tensorFile_0_2_MPORT_mask; // @[TensorStoreNarrowVME.scala 167:16]
  wire  tensorFile_0_2_MPORT_en; // @[TensorStoreNarrowVME.scala 167:16]
  reg  tensorFile_0_2_MPORT_1_en_pipe_0;
  reg [6:0] tensorFile_0_2_MPORT_1_addr_pipe_0;
  reg [63:0] tensorFile_0_3 [0:127]; // @[TensorStoreNarrowVME.scala 167:16]
  wire  tensorFile_0_3_MPORT_1_en; // @[TensorStoreNarrowVME.scala 167:16]
  wire [6:0] tensorFile_0_3_MPORT_1_addr; // @[TensorStoreNarrowVME.scala 167:16]
  wire [63:0] tensorFile_0_3_MPORT_1_data; // @[TensorStoreNarrowVME.scala 167:16]
  wire [63:0] tensorFile_0_3_MPORT_data; // @[TensorStoreNarrowVME.scala 167:16]
  wire [6:0] tensorFile_0_3_MPORT_addr; // @[TensorStoreNarrowVME.scala 167:16]
  wire  tensorFile_0_3_MPORT_mask; // @[TensorStoreNarrowVME.scala 167:16]
  wire  tensorFile_0_3_MPORT_en; // @[TensorStoreNarrowVME.scala 167:16]
  reg  tensorFile_0_3_MPORT_1_en_pipe_0;
  reg [6:0] tensorFile_0_3_MPORT_1_addr_pipe_0;
  wire [15:0] dec_sram_offset = io_inst[25:10]; // @[TensorStoreNarrowVME.scala 60:29]
  wire [31:0] dec_dram_offset = io_inst[57:26]; // @[TensorStoreNarrowVME.scala 60:29]
  wire [15:0] dec_ysize = io_inst[79:64]; // @[TensorStoreNarrowVME.scala 60:29]
  wire [15:0] dec_xsize = io_inst[95:80]; // @[TensorStoreNarrowVME.scala 60:29]
  wire [15:0] dec_xstride = io_inst[111:96]; // @[TensorStoreNarrowVME.scala 60:29]
  reg [31:0] waddr_cur; // @[TensorStoreNarrowVME.scala 61:22]
  reg [31:0] waddr_nxt; // @[TensorStoreNarrowVME.scala 62:22]
  reg [3:0] xcnt; // @[TensorStoreNarrowVME.scala 63:17]
  reg [3:0] xlen; // @[TensorStoreNarrowVME.scala 64:17]
  reg [15:0] xrem; // @[TensorStoreNarrowVME.scala 65:17]
  wire [17:0] xsize = {dec_xsize, 2'h0}; // @[TensorStoreNarrowVME.scala 66:26]
  reg [15:0] ycnt; // @[TensorStoreNarrowVME.scala 69:17]
  reg [7:0] tag; // @[TensorStoreNarrowVME.scala 71:16]
  reg [7:0] set; // @[TensorStoreNarrowVME.scala 72:16]
  reg [31:0] xfer_bytes; // @[TensorStoreNarrowVME.scala 74:23]
  wire [20:0] xstride_bytes = {dec_xstride, 5'h0}; // @[TensorStoreNarrowVME.scala 75:35]
  wire [36:0] _xfer_init_addr_T = {dec_dram_offset, 5'h0}; // @[TensorStoreNarrowVME.scala 80:66]
  wire [36:0] _xfer_init_addr_T_1 = 37'hffffffff & _xfer_init_addr_T; // @[TensorStoreNarrowVME.scala 80:47]
  wire [36:0] _GEN_94 = {{5'd0}, io_baddr}; // @[TensorStoreNarrowVME.scala 80:33]
  wire [36:0] xfer_init_addr = _GEN_94 | _xfer_init_addr_T_1; // @[TensorStoreNarrowVME.scala 80:33]
  wire [31:0] xfer_split_addr = waddr_cur + xfer_bytes; // @[TensorStoreNarrowVME.scala 81:35]
  wire [31:0] _GEN_95 = {{11'd0}, xstride_bytes}; // @[TensorStoreNarrowVME.scala 82:36]
  wire [31:0] xfer_stride_addr = waddr_nxt + _GEN_95; // @[TensorStoreNarrowVME.scala 82:36]
  wire [36:0] _GEN_2 = xfer_init_addr % 37'h80; // @[TensorStoreNarrowVME.scala 84:55]
  wire [7:0] _xfer_init_bytes_T = _GEN_2[7:0]; // @[TensorStoreNarrowVME.scala 84:55]
  wire [7:0] xfer_init_bytes = 8'h80 - _xfer_init_bytes_T; // @[TensorStoreNarrowVME.scala 84:38]
  wire [4:0] xfer_init_pulses = xfer_init_bytes[7:3]; // @[TensorStoreNarrowVME.scala 85:43]
  wire [31:0] _GEN_5 = xfer_split_addr % 32'h80; // @[TensorStoreNarrowVME.scala 86:56]
  wire [7:0] _xfer_split_bytes_T = _GEN_5[7:0]; // @[TensorStoreNarrowVME.scala 86:56]
  wire [7:0] xfer_split_bytes = 8'h80 - _xfer_split_bytes_T; // @[TensorStoreNarrowVME.scala 86:38]
  wire [4:0] xfer_split_pulses = xfer_split_bytes[7:3]; // @[TensorStoreNarrowVME.scala 87:44]
  wire [31:0] _GEN_15 = xfer_stride_addr % 32'h80; // @[TensorStoreNarrowVME.scala 88:57]
  wire [7:0] _xfer_stride_bytes_T = _GEN_15[7:0]; // @[TensorStoreNarrowVME.scala 88:57]
  wire [7:0] xfer_stride_bytes = 8'h80 - _xfer_stride_bytes_T; // @[TensorStoreNarrowVME.scala 88:38]
  wire [4:0] xfer_stride_pulses = xfer_stride_bytes[7:3]; // @[TensorStoreNarrowVME.scala 89:45]
  reg [2:0] state; // @[TensorStoreNarrowVME.scala 92:22]
  wire  _T = 3'h0 == state; // @[TensorStoreNarrowVME.scala 95:17]
  wire [17:0] _GEN_96 = {{13'd0}, xfer_init_pulses}; // @[TensorStoreNarrowVME.scala 100:21]
  wire  _T_1 = xsize < _GEN_96; // @[TensorStoreNarrowVME.scala 100:21]
  wire  _T_2 = xsize > 18'h0; // @[TensorStoreNarrowVME.scala 101:24]
  wire  _T_4 = ~reset; // @[TensorStoreNarrowVME.scala 101:17]
  wire  _T_5 = ~(xsize > 18'h0); // @[TensorStoreNarrowVME.scala 101:17]
  wire [17:0] _xlen_T_1 = xsize - 18'h1; // @[TensorStoreNarrowVME.scala 102:25]
  wire [4:0] _xlen_T_3 = xfer_init_pulses - 5'h1; // @[TensorStoreNarrowVME.scala 105:36]
  wire [17:0] _xrem_T_1 = xsize - _GEN_96; // @[TensorStoreNarrowVME.scala 107:25]
  wire [17:0] _GEN_0 = xsize < _GEN_96 ? _xlen_T_1 : {{13'd0}, _xlen_T_3}; // @[TensorStoreNarrowVME.scala 100:41 102:16 105:16]
  wire [17:0] _GEN_1 = xsize < _GEN_96 ? 18'h0 : _xrem_T_1; // @[TensorStoreNarrowVME.scala 100:41 103:16 107:16]
  wire [17:0] _GEN_3 = io_start ? _GEN_0 : {{14'd0}, xlen}; // @[TensorStoreNarrowVME.scala 64:17 98:25]
  wire [17:0] _GEN_4 = io_start ? _GEN_1 : {{2'd0}, xrem}; // @[TensorStoreNarrowVME.scala 65:17 98:25]
  wire  _T_10 = 3'h1 == state; // @[TensorStoreNarrowVME.scala 95:17]
  wire  _T_11 = 3'h2 == state; // @[TensorStoreNarrowVME.scala 95:17]
  wire  _T_13 = tag == 8'h3; // @[TensorStoreNarrowVME.scala 120:24]
  wire [2:0] _GEN_6 = tag == 8'h3 ? 3'h3 : state; // @[TensorStoreNarrowVME.scala 120:49 121:17 92:22]
  wire [2:0] _GEN_7 = xcnt == xlen ? 3'h4 : _GEN_6; // @[TensorStoreNarrowVME.scala 118:29 119:17]
  wire [2:0] _GEN_8 = io_vme_wr_data_ready ? _GEN_7 : state; // @[TensorStoreNarrowVME.scala 117:34 92:22]
  wire  _T_14 = 3'h3 == state; // @[TensorStoreNarrowVME.scala 95:17]
  wire  _T_15 = 3'h4 == state; // @[TensorStoreNarrowVME.scala 95:17]
  wire  _T_16 = xrem == 16'h0; // @[TensorStoreNarrowVME.scala 130:19]
  wire [15:0] _T_18 = dec_ysize - 16'h1; // @[TensorStoreNarrowVME.scala 131:31]
  wire  _T_19 = ycnt == _T_18; // @[TensorStoreNarrowVME.scala 131:21]
  wire [17:0] _GEN_99 = {{13'd0}, xfer_stride_pulses}; // @[TensorStoreNarrowVME.scala 136:24]
  wire  _T_20 = xsize < _GEN_99; // @[TensorStoreNarrowVME.scala 136:24]
  wire [4:0] _xlen_T_7 = xfer_stride_pulses - 5'h1; // @[TensorStoreNarrowVME.scala 141:42]
  wire [17:0] _xrem_T_3 = xsize - _GEN_99; // @[TensorStoreNarrowVME.scala 143:29]
  wire [17:0] _GEN_9 = xsize < _GEN_99 ? _xlen_T_1 : {{13'd0}, _xlen_T_7}; // @[TensorStoreNarrowVME.scala 136:46 138:20 141:20]
  wire [17:0] _GEN_10 = xsize < _GEN_99 ? 18'h0 : _xrem_T_3; // @[TensorStoreNarrowVME.scala 136:46 139:20 143:20]
  wire [2:0] _GEN_11 = ycnt == _T_18 ? 3'h0 : 3'h1; // @[TensorStoreNarrowVME.scala 131:38 132:19 134:19]
  wire [31:0] _GEN_12 = ycnt == _T_18 ? xfer_bytes : {{24'd0}, xfer_stride_bytes}; // @[TensorStoreNarrowVME.scala 131:38 74:23 135:24]
  wire [17:0] _GEN_13 = ycnt == _T_18 ? {{14'd0}, xlen} : _GEN_9; // @[TensorStoreNarrowVME.scala 131:38 64:17]
  wire [17:0] _GEN_14 = ycnt == _T_18 ? {{2'd0}, xrem} : _GEN_10; // @[TensorStoreNarrowVME.scala 131:38 65:17]
  wire [15:0] _GEN_102 = {{11'd0}, xfer_split_pulses}; // @[TensorStoreNarrowVME.scala 147:24]
  wire  _T_29 = xrem < _GEN_102; // @[TensorStoreNarrowVME.scala 147:24]
  wire [15:0] _xlen_T_9 = xrem - 16'h1; // @[TensorStoreNarrowVME.scala 151:24]
  wire [4:0] _xlen_T_11 = xfer_split_pulses - 5'h1; // @[TensorStoreNarrowVME.scala 157:37]
  wire [15:0] _xrem_T_5 = xrem - _GEN_102; // @[TensorStoreNarrowVME.scala 159:24]
  wire [15:0] _GEN_17 = xrem < _GEN_102 ? _xlen_T_9 : {{11'd0}, _xlen_T_11}; // @[TensorStoreNarrowVME.scala 147:45 151:16 157:16]
  wire [15:0] _GEN_18 = xrem < _GEN_102 ? 16'h0 : _xrem_T_5; // @[TensorStoreNarrowVME.scala 147:45 152:16 159:16]
  wire [2:0] _GEN_19 = xrem == 16'h0 ? _GEN_11 : 3'h1; // @[TensorStoreNarrowVME.scala 130:28]
  wire [31:0] _GEN_20 = xrem == 16'h0 ? _GEN_12 : {{24'd0}, xfer_split_bytes}; // @[TensorStoreNarrowVME.scala 130:28]
  wire [17:0] _GEN_21 = xrem == 16'h0 ? _GEN_13 : {{2'd0}, _GEN_17}; // @[TensorStoreNarrowVME.scala 130:28]
  wire [17:0] _GEN_22 = xrem == 16'h0 ? _GEN_14 : {{2'd0}, _GEN_18}; // @[TensorStoreNarrowVME.scala 130:28]
  wire [2:0] _GEN_23 = io_vme_wr_ack ? _GEN_19 : state; // @[TensorStoreNarrowVME.scala 129:27 92:22]
  wire [31:0] _GEN_24 = io_vme_wr_ack ? _GEN_20 : xfer_bytes; // @[TensorStoreNarrowVME.scala 129:27 74:23]
  wire [17:0] _GEN_25 = io_vme_wr_ack ? _GEN_21 : {{14'd0}, xlen}; // @[TensorStoreNarrowVME.scala 129:27 64:17]
  wire [17:0] _GEN_26 = io_vme_wr_ack ? _GEN_22 : {{2'd0}, xrem}; // @[TensorStoreNarrowVME.scala 129:27 65:17]
  wire [2:0] _GEN_27 = 3'h4 == state ? _GEN_23 : state; // @[TensorStoreNarrowVME.scala 95:17 92:22]
  wire [31:0] _GEN_28 = 3'h4 == state ? _GEN_24 : xfer_bytes; // @[TensorStoreNarrowVME.scala 95:17 74:23]
  wire [17:0] _GEN_29 = 3'h4 == state ? _GEN_25 : {{14'd0}, xlen}; // @[TensorStoreNarrowVME.scala 64:17 95:17]
  wire [17:0] _GEN_30 = 3'h4 == state ? _GEN_26 : {{2'd0}, xrem}; // @[TensorStoreNarrowVME.scala 65:17 95:17]
  wire [2:0] _GEN_31 = 3'h3 == state ? 3'h2 : _GEN_27; // @[TensorStoreNarrowVME.scala 126:13 95:17]
  wire [17:0] _GEN_33 = 3'h3 == state ? {{14'd0}, xlen} : _GEN_29; // @[TensorStoreNarrowVME.scala 64:17 95:17]
  wire [17:0] _GEN_34 = 3'h3 == state ? {{2'd0}, xrem} : _GEN_30; // @[TensorStoreNarrowVME.scala 65:17 95:17]
  wire [17:0] _GEN_37 = 3'h2 == state ? {{14'd0}, xlen} : _GEN_33; // @[TensorStoreNarrowVME.scala 64:17 95:17]
  wire [17:0] _GEN_38 = 3'h2 == state ? {{2'd0}, xrem} : _GEN_34; // @[TensorStoreNarrowVME.scala 65:17 95:17]
  wire [17:0] _GEN_41 = 3'h1 == state ? {{14'd0}, xlen} : _GEN_37; // @[TensorStoreNarrowVME.scala 64:17 95:17]
  wire [17:0] _GEN_42 = 3'h1 == state ? {{2'd0}, xrem} : _GEN_38; // @[TensorStoreNarrowVME.scala 65:17 95:17]
  wire [17:0] _GEN_45 = 3'h0 == state ? _GEN_3 : _GEN_41; // @[TensorStoreNarrowVME.scala 95:17]
  wire [17:0] _GEN_46 = 3'h0 == state ? _GEN_4 : _GEN_42; // @[TensorStoreNarrowVME.scala 95:17]
  wire [63:0] inWrData_lo_lo = {io_tensor_wr_0_bits_data_0_7,io_tensor_wr_0_bits_data_0_6,io_tensor_wr_0_bits_data_0_5,
    io_tensor_wr_0_bits_data_0_4,io_tensor_wr_0_bits_data_0_3,io_tensor_wr_0_bits_data_0_2,io_tensor_wr_0_bits_data_0_1,
    io_tensor_wr_0_bits_data_0_0}; // @[TensorStoreNarrowVME.scala 178:49]
  wire [127:0] inWrData_lo = {io_tensor_wr_0_bits_data_0_15,io_tensor_wr_0_bits_data_0_14,io_tensor_wr_0_bits_data_0_13,
    io_tensor_wr_0_bits_data_0_12,io_tensor_wr_0_bits_data_0_11,io_tensor_wr_0_bits_data_0_10,
    io_tensor_wr_0_bits_data_0_9,io_tensor_wr_0_bits_data_0_8,inWrData_lo_lo}; // @[TensorStoreNarrowVME.scala 178:49]
  wire [63:0] inWrData_hi_lo = {io_tensor_wr_0_bits_data_0_23,io_tensor_wr_0_bits_data_0_22,
    io_tensor_wr_0_bits_data_0_21,io_tensor_wr_0_bits_data_0_20,io_tensor_wr_0_bits_data_0_19,
    io_tensor_wr_0_bits_data_0_18,io_tensor_wr_0_bits_data_0_17,io_tensor_wr_0_bits_data_0_16}; // @[TensorStoreNarrowVME.scala 178:49]
  wire [255:0] _inWrData_T = {io_tensor_wr_0_bits_data_0_31,io_tensor_wr_0_bits_data_0_30,io_tensor_wr_0_bits_data_0_29,
    io_tensor_wr_0_bits_data_0_28,io_tensor_wr_0_bits_data_0_27,io_tensor_wr_0_bits_data_0_26,
    io_tensor_wr_0_bits_data_0_25,io_tensor_wr_0_bits_data_0_24,inWrData_hi_lo,inWrData_lo}; // @[TensorStoreNarrowVME.scala 178:49]
  wire  _stride_T_1 = state == 3'h4 & io_vme_wr_ack; // @[TensorStoreNarrowVME.scala 186:36]
  wire [3:0] _stride_T_3 = xlen + 4'h1; // @[TensorStoreNarrowVME.scala 188:19]
  wire  _stride_T_4 = xcnt == _stride_T_3; // @[TensorStoreNarrowVME.scala 188:10]
  wire  _stride_T_5 = _stride_T_1 & _stride_T_4; // @[TensorStoreNarrowVME.scala 187:19]
  wire  _stride_T_7 = _stride_T_5 & _T_16; // @[TensorStoreNarrowVME.scala 188:25]
  wire  _stride_T_10 = ycnt != _T_18; // @[TensorStoreNarrowVME.scala 190:10]
  wire  stride = _stride_T_7 & _stride_T_10; // @[TensorStoreNarrowVME.scala 189:18]
  wire  _T_38 = state == 3'h0; // @[TensorStoreNarrowVME.scala 192:14]
  wire [15:0] _ycnt_T_1 = ycnt + 16'h1; // @[TensorStoreNarrowVME.scala 195:18]
  wire  _T_39 = state == 3'h1; // @[TensorStoreNarrowVME.scala 198:14]
  wire  _T_42 = io_vme_wr_data_ready & io_vme_wr_data_valid; // @[Decoupled.scala 50:35]
  wire [7:0] _tag_T_1 = tag + 8'h1; // @[TensorStoreNarrowVME.scala 201:16]
  wire  _T_45 = set == 8'h0; // @[TensorStoreNarrowVME.scala 205:55]
  wire [7:0] _set_T_1 = set + 8'h1; // @[TensorStoreNarrowVME.scala 208:16]
  reg [6:0] raddr_cur; // @[TensorStoreNarrowVME.scala 211:22]
  reg [6:0] raddr_nxt; // @[TensorStoreNarrowVME.scala 212:22]
  wire [6:0] _raddr_cur_T_1 = raddr_cur + 7'h1; // @[TensorStoreNarrowVME.scala 217:28]
  wire [15:0] _GEN_105 = {{9'd0}, raddr_nxt}; // @[TensorStoreNarrowVME.scala 219:28]
  wire [15:0] _raddr_cur_T_3 = _GEN_105 + dec_xsize; // @[TensorStoreNarrowVME.scala 219:28]
  wire [15:0] _GEN_72 = stride ? _raddr_cur_T_3 : {{9'd0}, raddr_cur}; // @[TensorStoreNarrowVME.scala 218:22 219:15 211:22]
  wire [15:0] _GEN_73 = stride ? _raddr_cur_T_3 : {{9'd0}, raddr_nxt}; // @[TensorStoreNarrowVME.scala 218:22 220:15 212:22]
  wire [15:0] _GEN_74 = _T_42 & _T_45 & _T_13 ? {{9'd0}, _raddr_cur_T_1} : _GEN_72; // @[TensorStoreNarrowVME.scala 216:98 217:15]
  wire [15:0] _GEN_75 = _T_42 & _T_45 & _T_13 ? {{9'd0}, raddr_nxt} : _GEN_73; // @[TensorStoreNarrowVME.scala 212:22 216:98]
  wire [15:0] _GEN_76 = _T_38 ? dec_sram_offset : _GEN_74; // @[TensorStoreNarrowVME.scala 213:25 214:15]
  wire [15:0] _GEN_77 = _T_38 ? dec_sram_offset : _GEN_75; // @[TensorStoreNarrowVME.scala 213:25 215:15]
  wire  _T_60 = state == 3'h3; // @[TensorStoreNarrowVME.scala 225:65]
  wire [63:0] mdata_0 = 8'h0 == set ? tensorFile_0_0_MPORT_1_data : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] mdata_1 = 8'h0 == set ? tensorFile_0_1_MPORT_1_data : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] mdata_2 = 8'h0 == set ? tensorFile_0_2_MPORT_1_data : 64'h0; // @[Mux.scala 81:58]
  wire [63:0] mdata_3 = 8'h0 == set ? tensorFile_0_3_MPORT_1_data : 64'h0; // @[Mux.scala 81:58]
  wire [31:0] _GEN_82 = stride ? xfer_stride_addr : waddr_cur; // @[TensorStoreNarrowVME.scala 235:22 236:15 61:22]
  wire [31:0] _GEN_83 = stride ? xfer_stride_addr : waddr_nxt; // @[TensorStoreNarrowVME.scala 235:22 237:15 62:22]
  wire [31:0] _GEN_84 = _stride_T_1 & xrem != 16'h0 ? xfer_split_addr : _GEN_82; // @[TensorStoreNarrowVME.scala 233:68 234:15]
  wire [31:0] _GEN_85 = _stride_T_1 & xrem != 16'h0 ? waddr_nxt : _GEN_83; // @[TensorStoreNarrowVME.scala 233:68 62:22]
  wire [36:0] _GEN_86 = _T_38 ? xfer_init_addr : {{5'd0}, _GEN_84}; // @[TensorStoreNarrowVME.scala 230:25 231:15]
  wire [36:0] _GEN_87 = _T_38 ? xfer_init_addr : {{5'd0}, _GEN_85}; // @[TensorStoreNarrowVME.scala 230:25 232:15]
  wire [63:0] _GEN_89 = 2'h1 == tag[1:0] ? mdata_1 : mdata_0; // @[TensorStoreNarrowVME.scala 246:{28,28}]
  wire [63:0] _GEN_90 = 2'h2 == tag[1:0] ? mdata_2 : _GEN_89; // @[TensorStoreNarrowVME.scala 246:{28,28}]
  wire [3:0] _xcnt_T_1 = xcnt + 4'h1; // @[TensorStoreNarrowVME.scala 252:18]
  wire  _GEN_107 = _T & io_start; // @[TensorStoreNarrowVME.scala 101:17]
  wire  _GEN_127 = ~_T & ~_T_10 & ~_T_11 & ~_T_14 & _T_15 & io_vme_wr_ack; // @[TensorStoreNarrowVME.scala 137:21]
  wire  _GEN_130 = ~_T & ~_T_10 & ~_T_11 & ~_T_14 & _T_15 & io_vme_wr_ack & _T_16 & ~_T_19; // @[TensorStoreNarrowVME.scala 137:21]
  wire  _GEN_185 = _GEN_127 & ~_T_16; // @[TensorStoreNarrowVME.scala 150:17]
  assign tensorFile_0_0_MPORT_1_en = tensorFile_0_0_MPORT_1_en_pipe_0;
  assign tensorFile_0_0_MPORT_1_addr = tensorFile_0_0_MPORT_1_addr_pipe_0;
  assign tensorFile_0_0_MPORT_1_data = tensorFile_0_0[tensorFile_0_0_MPORT_1_addr]; // @[TensorStoreNarrowVME.scala 167:16]
  assign tensorFile_0_0_MPORT_data = _inWrData_T[63:0];
  assign tensorFile_0_0_MPORT_addr = io_tensor_wr_0_bits_idx;
  assign tensorFile_0_0_MPORT_mask = 1'h1;
  assign tensorFile_0_0_MPORT_en = io_tensor_wr_0_valid;
  assign tensorFile_0_1_MPORT_1_en = tensorFile_0_1_MPORT_1_en_pipe_0;
  assign tensorFile_0_1_MPORT_1_addr = tensorFile_0_1_MPORT_1_addr_pipe_0;
  assign tensorFile_0_1_MPORT_1_data = tensorFile_0_1[tensorFile_0_1_MPORT_1_addr]; // @[TensorStoreNarrowVME.scala 167:16]
  assign tensorFile_0_1_MPORT_data = _inWrData_T[127:64];
  assign tensorFile_0_1_MPORT_addr = io_tensor_wr_0_bits_idx;
  assign tensorFile_0_1_MPORT_mask = 1'h1;
  assign tensorFile_0_1_MPORT_en = io_tensor_wr_0_valid;
  assign tensorFile_0_2_MPORT_1_en = tensorFile_0_2_MPORT_1_en_pipe_0;
  assign tensorFile_0_2_MPORT_1_addr = tensorFile_0_2_MPORT_1_addr_pipe_0;
  assign tensorFile_0_2_MPORT_1_data = tensorFile_0_2[tensorFile_0_2_MPORT_1_addr]; // @[TensorStoreNarrowVME.scala 167:16]
  assign tensorFile_0_2_MPORT_data = _inWrData_T[191:128];
  assign tensorFile_0_2_MPORT_addr = io_tensor_wr_0_bits_idx;
  assign tensorFile_0_2_MPORT_mask = 1'h1;
  assign tensorFile_0_2_MPORT_en = io_tensor_wr_0_valid;
  assign tensorFile_0_3_MPORT_1_en = tensorFile_0_3_MPORT_1_en_pipe_0;
  assign tensorFile_0_3_MPORT_1_addr = tensorFile_0_3_MPORT_1_addr_pipe_0;
  assign tensorFile_0_3_MPORT_1_data = tensorFile_0_3[tensorFile_0_3_MPORT_1_addr]; // @[TensorStoreNarrowVME.scala 167:16]
  assign tensorFile_0_3_MPORT_data = _inWrData_T[255:192];
  assign tensorFile_0_3_MPORT_addr = io_tensor_wr_0_bits_idx;
  assign tensorFile_0_3_MPORT_mask = 1'h1;
  assign tensorFile_0_3_MPORT_en = io_tensor_wr_0_valid;
  assign io_done = _stride_T_1 & _T_16 & _T_19; // @[TensorStoreNarrowVME.scala 259:65]
  assign io_vme_wr_cmd_valid = state == 3'h1; // @[TensorStoreNarrowVME.scala 240:32]
  assign io_vme_wr_cmd_bits_addr = waddr_cur; // @[TensorStoreNarrowVME.scala 241:27]
  assign io_vme_wr_cmd_bits_len = xlen; // @[TensorStoreNarrowVME.scala 242:26]
  assign io_vme_wr_data_valid = state == 3'h2; // @[TensorStoreNarrowVME.scala 245:33]
  assign io_vme_wr_data_bits_data = 2'h3 == tag[1:0] ? mdata_3 : _GEN_90; // @[TensorStoreNarrowVME.scala 246:{28,28}]
  always @(posedge clock) begin
    if (tensorFile_0_0_MPORT_en & tensorFile_0_0_MPORT_mask) begin
      tensorFile_0_0[tensorFile_0_0_MPORT_addr] <= tensorFile_0_0_MPORT_data; // @[TensorStoreNarrowVME.scala 167:16]
    end
    tensorFile_0_0_MPORT_1_en_pipe_0 <= _T_39 | _T_60;
    if (_T_39 | _T_60) begin
      tensorFile_0_0_MPORT_1_addr_pipe_0 <= raddr_cur;
    end
    if (tensorFile_0_1_MPORT_en & tensorFile_0_1_MPORT_mask) begin
      tensorFile_0_1[tensorFile_0_1_MPORT_addr] <= tensorFile_0_1_MPORT_data; // @[TensorStoreNarrowVME.scala 167:16]
    end
    tensorFile_0_1_MPORT_1_en_pipe_0 <= _T_39 | _T_60;
    if (_T_39 | _T_60) begin
      tensorFile_0_1_MPORT_1_addr_pipe_0 <= raddr_cur;
    end
    if (tensorFile_0_2_MPORT_en & tensorFile_0_2_MPORT_mask) begin
      tensorFile_0_2[tensorFile_0_2_MPORT_addr] <= tensorFile_0_2_MPORT_data; // @[TensorStoreNarrowVME.scala 167:16]
    end
    tensorFile_0_2_MPORT_1_en_pipe_0 <= _T_39 | _T_60;
    if (_T_39 | _T_60) begin
      tensorFile_0_2_MPORT_1_addr_pipe_0 <= raddr_cur;
    end
    if (tensorFile_0_3_MPORT_en & tensorFile_0_3_MPORT_mask) begin
      tensorFile_0_3[tensorFile_0_3_MPORT_addr] <= tensorFile_0_3_MPORT_data; // @[TensorStoreNarrowVME.scala 167:16]
    end
    tensorFile_0_3_MPORT_1_en_pipe_0 <= _T_39 | _T_60;
    if (_T_39 | _T_60) begin
      tensorFile_0_3_MPORT_1_addr_pipe_0 <= raddr_cur;
    end
    waddr_cur <= _GEN_86[31:0];
    waddr_nxt <= _GEN_87[31:0];
    if (_T_39) begin // @[TensorStoreNarrowVME.scala 249:29]
      xcnt <= 4'h0; // @[TensorStoreNarrowVME.scala 250:10]
    end else if (_T_42) begin // @[TensorStoreNarrowVME.scala 251:35]
      xcnt <= _xcnt_T_1; // @[TensorStoreNarrowVME.scala 252:10]
    end
    xlen <= _GEN_45[3:0];
    xrem <= _GEN_46[15:0];
    if (state == 3'h0) begin // @[TensorStoreNarrowVME.scala 192:25]
      ycnt <= 16'h0; // @[TensorStoreNarrowVME.scala 193:10]
    end else if (stride) begin // @[TensorStoreNarrowVME.scala 194:22]
      ycnt <= _ycnt_T_1; // @[TensorStoreNarrowVME.scala 195:10]
    end
    if (state == 3'h1 | _T_13) begin // @[TensorStoreNarrowVME.scala 198:60]
      tag <= 8'h0; // @[TensorStoreNarrowVME.scala 199:9]
    end else if (_T_42) begin // @[TensorStoreNarrowVME.scala 200:35]
      tag <= _tag_T_1; // @[TensorStoreNarrowVME.scala 201:9]
    end
    if (_T_39 | state != 3'h3 & set == 8'h0 & _T_13) begin // @[TensorStoreNarrowVME.scala 205:113]
      set <= 8'h0; // @[TensorStoreNarrowVME.scala 206:9]
    end else if (_T_42 & _T_13) begin // @[TensorStoreNarrowVME.scala 207:66]
      set <= _set_T_1; // @[TensorStoreNarrowVME.scala 208:9]
    end
    if (3'h0 == state) begin // @[TensorStoreNarrowVME.scala 95:17]
      xfer_bytes <= {{24'd0}, xfer_init_bytes}; // @[TensorStoreNarrowVME.scala 97:18]
    end else if (!(3'h1 == state)) begin // @[TensorStoreNarrowVME.scala 95:17]
      if (!(3'h2 == state)) begin // @[TensorStoreNarrowVME.scala 95:17]
        if (!(3'h3 == state)) begin // @[TensorStoreNarrowVME.scala 95:17]
          xfer_bytes <= _GEN_28;
        end
      end
    end
    if (reset) begin // @[TensorStoreNarrowVME.scala 92:22]
      state <= 3'h0; // @[TensorStoreNarrowVME.scala 92:22]
    end else if (3'h0 == state) begin // @[TensorStoreNarrowVME.scala 95:17]
      if (io_start) begin // @[TensorStoreNarrowVME.scala 98:25]
        state <= 3'h1; // @[TensorStoreNarrowVME.scala 99:15]
      end
    end else if (3'h1 == state) begin // @[TensorStoreNarrowVME.scala 95:17]
      if (io_vme_wr_cmd_ready) begin // @[TensorStoreNarrowVME.scala 112:33]
        state <= 3'h2; // @[TensorStoreNarrowVME.scala 113:15]
      end
    end else if (3'h2 == state) begin // @[TensorStoreNarrowVME.scala 95:17]
      state <= _GEN_8;
    end else begin
      state <= _GEN_31;
    end
    raddr_cur <= _GEN_76[6:0];
    raddr_nxt <= _GEN_77[6:0];
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T & io_start & _T_1 & ~reset & ~(xsize > 18'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TensorStoreNarrowVME.scala:101 assert(xsize > 0.U)\n"); // @[TensorStoreNarrowVME.scala 101:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_107 & ~_T_1 & _T_4 & ~(xsize >= _GEN_96)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorStoreNarrowVME.scala:106 assert(xsize >= xfer_init_pulses)\n"); // @[TensorStoreNarrowVME.scala 106:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (~_T & ~_T_10 & ~_T_11 & ~_T_14 & _T_15 & io_vme_wr_ack & _T_16 & ~_T_19 & _T_20 & _T_4 & _T_5) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TensorStoreNarrowVME.scala:137 assert(xsize > 0.U)\n"); // @[TensorStoreNarrowVME.scala 137:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_130 & ~_T_20 & _T_4 & ~(xsize >= _GEN_99)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorStoreNarrowVME.scala:142 assert(xsize >= xfer_stride_pulses)\n"); // @[TensorStoreNarrowVME.scala 142:21]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_127 & ~_T_16 & _T_29 & _T_4 & ~(xrem > 16'h0)) begin
          $fwrite(32'h80000002,"Assertion failed\n    at TensorStoreNarrowVME.scala:150 assert(xrem > 0.U)\n"); // @[TensorStoreNarrowVME.scala 150:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_185 & ~_T_29 & _T_4 & ~(xrem >= _GEN_102)) begin
          $fwrite(32'h80000002,
            "Assertion failed\n    at TensorStoreNarrowVME.scala:158 assert(xrem >= xfer_split_pulses)\n"); // @[TensorStoreNarrowVME.scala 158:17]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_0_0[initvar] = _RAND_0[63:0];
  _RAND_3 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_0_1[initvar] = _RAND_3[63:0];
  _RAND_6 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_0_2[initvar] = _RAND_6[63:0];
  _RAND_9 = {2{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tensorFile_0_3[initvar] = _RAND_9[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  tensorFile_0_0_MPORT_1_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  tensorFile_0_0_MPORT_1_addr_pipe_0 = _RAND_2[6:0];
  _RAND_4 = {1{`RANDOM}};
  tensorFile_0_1_MPORT_1_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  tensorFile_0_1_MPORT_1_addr_pipe_0 = _RAND_5[6:0];
  _RAND_7 = {1{`RANDOM}};
  tensorFile_0_2_MPORT_1_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  tensorFile_0_2_MPORT_1_addr_pipe_0 = _RAND_8[6:0];
  _RAND_10 = {1{`RANDOM}};
  tensorFile_0_3_MPORT_1_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  tensorFile_0_3_MPORT_1_addr_pipe_0 = _RAND_11[6:0];
  _RAND_12 = {1{`RANDOM}};
  waddr_cur = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  waddr_nxt = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  xcnt = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  xlen = _RAND_15[3:0];
  _RAND_16 = {1{`RANDOM}};
  xrem = _RAND_16[15:0];
  _RAND_17 = {1{`RANDOM}};
  ycnt = _RAND_17[15:0];
  _RAND_18 = {1{`RANDOM}};
  tag = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  set = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  xfer_bytes = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  state = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  raddr_cur = _RAND_22[6:0];
  _RAND_23 = {1{`RANDOM}};
  raddr_nxt = _RAND_23[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    //
    if (_T & io_start & _T_1 & ~reset) begin
      assert(xsize > 18'h0); // @[TensorStoreNarrowVME.scala 101:17]
    end
    //
    if (_GEN_107 & ~_T_1 & _T_4) begin
      assert(xsize >= _GEN_96); // @[TensorStoreNarrowVME.scala 106:17]
    end
    //
    if (~_T & ~_T_10 & ~_T_11 & ~_T_14 & _T_15 & io_vme_wr_ack & _T_16 & ~_T_19 & _T_20 & _T_4) begin
      assert(_T_2); // @[TensorStoreNarrowVME.scala 137:21]
    end
    //
    if (_GEN_130 & ~_T_20 & _T_4) begin
      assert(xsize >= _GEN_99); // @[TensorStoreNarrowVME.scala 142:21]
    end
    //
    if (_GEN_127 & ~_T_16 & _T_29 & _T_4) begin
      assert(xrem > 16'h0); // @[TensorStoreNarrowVME.scala 150:17]
    end
    //
    if (_GEN_185 & ~_T_29 & _T_4) begin
      assert(xrem >= _GEN_102); // @[TensorStoreNarrowVME.scala 158:17]
    end
  end
endmodule
module TensorStoreOut(
  input          clock,
  input          reset,
  input          io_start,
  output         io_done,
  input  [127:0] io_inst,
  input  [31:0]  io_baddr,
  input          io_vme_wr_cmd_ready,
  output         io_vme_wr_cmd_valid,
  output [31:0]  io_vme_wr_cmd_bits_addr,
  output [3:0]   io_vme_wr_cmd_bits_len,
  input          io_vme_wr_data_ready,
  output         io_vme_wr_data_valid,
  output [63:0]  io_vme_wr_data_bits_data,
  input          io_vme_wr_ack,
  input          io_tensor_wr_0_valid,
  input  [6:0]   io_tensor_wr_0_bits_idx,
  input  [7:0]   io_tensor_wr_0_bits_data_0_0,
  input  [7:0]   io_tensor_wr_0_bits_data_0_1,
  input  [7:0]   io_tensor_wr_0_bits_data_0_2,
  input  [7:0]   io_tensor_wr_0_bits_data_0_3,
  input  [7:0]   io_tensor_wr_0_bits_data_0_4,
  input  [7:0]   io_tensor_wr_0_bits_data_0_5,
  input  [7:0]   io_tensor_wr_0_bits_data_0_6,
  input  [7:0]   io_tensor_wr_0_bits_data_0_7,
  input  [7:0]   io_tensor_wr_0_bits_data_0_8,
  input  [7:0]   io_tensor_wr_0_bits_data_0_9,
  input  [7:0]   io_tensor_wr_0_bits_data_0_10,
  input  [7:0]   io_tensor_wr_0_bits_data_0_11,
  input  [7:0]   io_tensor_wr_0_bits_data_0_12,
  input  [7:0]   io_tensor_wr_0_bits_data_0_13,
  input  [7:0]   io_tensor_wr_0_bits_data_0_14,
  input  [7:0]   io_tensor_wr_0_bits_data_0_15,
  input  [7:0]   io_tensor_wr_0_bits_data_0_16,
  input  [7:0]   io_tensor_wr_0_bits_data_0_17,
  input  [7:0]   io_tensor_wr_0_bits_data_0_18,
  input  [7:0]   io_tensor_wr_0_bits_data_0_19,
  input  [7:0]   io_tensor_wr_0_bits_data_0_20,
  input  [7:0]   io_tensor_wr_0_bits_data_0_21,
  input  [7:0]   io_tensor_wr_0_bits_data_0_22,
  input  [7:0]   io_tensor_wr_0_bits_data_0_23,
  input  [7:0]   io_tensor_wr_0_bits_data_0_24,
  input  [7:0]   io_tensor_wr_0_bits_data_0_25,
  input  [7:0]   io_tensor_wr_0_bits_data_0_26,
  input  [7:0]   io_tensor_wr_0_bits_data_0_27,
  input  [7:0]   io_tensor_wr_0_bits_data_0_28,
  input  [7:0]   io_tensor_wr_0_bits_data_0_29,
  input  [7:0]   io_tensor_wr_0_bits_data_0_30,
  input  [7:0]   io_tensor_wr_0_bits_data_0_31
);
  wire  tensorStore_clock; // @[TensorStore.scala 59:29]
  wire  tensorStore_reset; // @[TensorStore.scala 59:29]
  wire  tensorStore_io_start; // @[TensorStore.scala 59:29]
  wire  tensorStore_io_done; // @[TensorStore.scala 59:29]
  wire [127:0] tensorStore_io_inst; // @[TensorStore.scala 59:29]
  wire [31:0] tensorStore_io_baddr; // @[TensorStore.scala 59:29]
  wire  tensorStore_io_vme_wr_cmd_ready; // @[TensorStore.scala 59:29]
  wire  tensorStore_io_vme_wr_cmd_valid; // @[TensorStore.scala 59:29]
  wire [31:0] tensorStore_io_vme_wr_cmd_bits_addr; // @[TensorStore.scala 59:29]
  wire [3:0] tensorStore_io_vme_wr_cmd_bits_len; // @[TensorStore.scala 59:29]
  wire  tensorStore_io_vme_wr_data_ready; // @[TensorStore.scala 59:29]
  wire  tensorStore_io_vme_wr_data_valid; // @[TensorStore.scala 59:29]
  wire [63:0] tensorStore_io_vme_wr_data_bits_data; // @[TensorStore.scala 59:29]
  wire  tensorStore_io_vme_wr_ack; // @[TensorStore.scala 59:29]
  wire  tensorStore_io_tensor_wr_0_valid; // @[TensorStore.scala 59:29]
  wire [6:0] tensorStore_io_tensor_wr_0_bits_idx; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_0; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_1; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_2; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_3; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_4; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_5; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_6; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_7; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_8; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_9; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_10; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_11; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_12; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_13; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_14; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_15; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_16; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_17; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_18; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_19; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_20; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_21; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_22; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_23; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_24; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_25; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_26; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_27; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_28; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_29; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_30; // @[TensorStore.scala 59:29]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_31; // @[TensorStore.scala 59:29]
  TensorStoreNarrowVME tensorStore ( // @[TensorStore.scala 59:29]
    .clock(tensorStore_clock),
    .reset(tensorStore_reset),
    .io_start(tensorStore_io_start),
    .io_done(tensorStore_io_done),
    .io_inst(tensorStore_io_inst),
    .io_baddr(tensorStore_io_baddr),
    .io_vme_wr_cmd_ready(tensorStore_io_vme_wr_cmd_ready),
    .io_vme_wr_cmd_valid(tensorStore_io_vme_wr_cmd_valid),
    .io_vme_wr_cmd_bits_addr(tensorStore_io_vme_wr_cmd_bits_addr),
    .io_vme_wr_cmd_bits_len(tensorStore_io_vme_wr_cmd_bits_len),
    .io_vme_wr_data_ready(tensorStore_io_vme_wr_data_ready),
    .io_vme_wr_data_valid(tensorStore_io_vme_wr_data_valid),
    .io_vme_wr_data_bits_data(tensorStore_io_vme_wr_data_bits_data),
    .io_vme_wr_ack(tensorStore_io_vme_wr_ack),
    .io_tensor_wr_0_valid(tensorStore_io_tensor_wr_0_valid),
    .io_tensor_wr_0_bits_idx(tensorStore_io_tensor_wr_0_bits_idx),
    .io_tensor_wr_0_bits_data_0_0(tensorStore_io_tensor_wr_0_bits_data_0_0),
    .io_tensor_wr_0_bits_data_0_1(tensorStore_io_tensor_wr_0_bits_data_0_1),
    .io_tensor_wr_0_bits_data_0_2(tensorStore_io_tensor_wr_0_bits_data_0_2),
    .io_tensor_wr_0_bits_data_0_3(tensorStore_io_tensor_wr_0_bits_data_0_3),
    .io_tensor_wr_0_bits_data_0_4(tensorStore_io_tensor_wr_0_bits_data_0_4),
    .io_tensor_wr_0_bits_data_0_5(tensorStore_io_tensor_wr_0_bits_data_0_5),
    .io_tensor_wr_0_bits_data_0_6(tensorStore_io_tensor_wr_0_bits_data_0_6),
    .io_tensor_wr_0_bits_data_0_7(tensorStore_io_tensor_wr_0_bits_data_0_7),
    .io_tensor_wr_0_bits_data_0_8(tensorStore_io_tensor_wr_0_bits_data_0_8),
    .io_tensor_wr_0_bits_data_0_9(tensorStore_io_tensor_wr_0_bits_data_0_9),
    .io_tensor_wr_0_bits_data_0_10(tensorStore_io_tensor_wr_0_bits_data_0_10),
    .io_tensor_wr_0_bits_data_0_11(tensorStore_io_tensor_wr_0_bits_data_0_11),
    .io_tensor_wr_0_bits_data_0_12(tensorStore_io_tensor_wr_0_bits_data_0_12),
    .io_tensor_wr_0_bits_data_0_13(tensorStore_io_tensor_wr_0_bits_data_0_13),
    .io_tensor_wr_0_bits_data_0_14(tensorStore_io_tensor_wr_0_bits_data_0_14),
    .io_tensor_wr_0_bits_data_0_15(tensorStore_io_tensor_wr_0_bits_data_0_15),
    .io_tensor_wr_0_bits_data_0_16(tensorStore_io_tensor_wr_0_bits_data_0_16),
    .io_tensor_wr_0_bits_data_0_17(tensorStore_io_tensor_wr_0_bits_data_0_17),
    .io_tensor_wr_0_bits_data_0_18(tensorStore_io_tensor_wr_0_bits_data_0_18),
    .io_tensor_wr_0_bits_data_0_19(tensorStore_io_tensor_wr_0_bits_data_0_19),
    .io_tensor_wr_0_bits_data_0_20(tensorStore_io_tensor_wr_0_bits_data_0_20),
    .io_tensor_wr_0_bits_data_0_21(tensorStore_io_tensor_wr_0_bits_data_0_21),
    .io_tensor_wr_0_bits_data_0_22(tensorStore_io_tensor_wr_0_bits_data_0_22),
    .io_tensor_wr_0_bits_data_0_23(tensorStore_io_tensor_wr_0_bits_data_0_23),
    .io_tensor_wr_0_bits_data_0_24(tensorStore_io_tensor_wr_0_bits_data_0_24),
    .io_tensor_wr_0_bits_data_0_25(tensorStore_io_tensor_wr_0_bits_data_0_25),
    .io_tensor_wr_0_bits_data_0_26(tensorStore_io_tensor_wr_0_bits_data_0_26),
    .io_tensor_wr_0_bits_data_0_27(tensorStore_io_tensor_wr_0_bits_data_0_27),
    .io_tensor_wr_0_bits_data_0_28(tensorStore_io_tensor_wr_0_bits_data_0_28),
    .io_tensor_wr_0_bits_data_0_29(tensorStore_io_tensor_wr_0_bits_data_0_29),
    .io_tensor_wr_0_bits_data_0_30(tensorStore_io_tensor_wr_0_bits_data_0_30),
    .io_tensor_wr_0_bits_data_0_31(tensorStore_io_tensor_wr_0_bits_data_0_31)
  );
  assign io_done = tensorStore_io_done; // @[TensorStore.scala 60:8]
  assign io_vme_wr_cmd_valid = tensorStore_io_vme_wr_cmd_valid; // @[TensorStore.scala 60:8]
  assign io_vme_wr_cmd_bits_addr = tensorStore_io_vme_wr_cmd_bits_addr; // @[TensorStore.scala 60:8]
  assign io_vme_wr_cmd_bits_len = tensorStore_io_vme_wr_cmd_bits_len; // @[TensorStore.scala 60:8]
  assign io_vme_wr_data_valid = tensorStore_io_vme_wr_data_valid; // @[TensorStore.scala 60:8]
  assign io_vme_wr_data_bits_data = tensorStore_io_vme_wr_data_bits_data; // @[TensorStore.scala 60:8]
  assign tensorStore_clock = clock;
  assign tensorStore_reset = reset;
  assign tensorStore_io_start = io_start; // @[TensorStore.scala 60:8]
  assign tensorStore_io_inst = io_inst; // @[TensorStore.scala 60:8]
  assign tensorStore_io_baddr = io_baddr; // @[TensorStore.scala 60:8]
  assign tensorStore_io_vme_wr_cmd_ready = io_vme_wr_cmd_ready; // @[TensorStore.scala 60:8]
  assign tensorStore_io_vme_wr_data_ready = io_vme_wr_data_ready; // @[TensorStore.scala 60:8]
  assign tensorStore_io_vme_wr_ack = io_vme_wr_ack; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_valid = io_tensor_wr_0_valid; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_idx = io_tensor_wr_0_bits_idx; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_0 = io_tensor_wr_0_bits_data_0_0; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_1 = io_tensor_wr_0_bits_data_0_1; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_2 = io_tensor_wr_0_bits_data_0_2; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_3 = io_tensor_wr_0_bits_data_0_3; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_4 = io_tensor_wr_0_bits_data_0_4; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_5 = io_tensor_wr_0_bits_data_0_5; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_6 = io_tensor_wr_0_bits_data_0_6; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_7 = io_tensor_wr_0_bits_data_0_7; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_8 = io_tensor_wr_0_bits_data_0_8; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_9 = io_tensor_wr_0_bits_data_0_9; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_10 = io_tensor_wr_0_bits_data_0_10; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_11 = io_tensor_wr_0_bits_data_0_11; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_12 = io_tensor_wr_0_bits_data_0_12; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_13 = io_tensor_wr_0_bits_data_0_13; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_14 = io_tensor_wr_0_bits_data_0_14; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_15 = io_tensor_wr_0_bits_data_0_15; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_16 = io_tensor_wr_0_bits_data_0_16; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_17 = io_tensor_wr_0_bits_data_0_17; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_18 = io_tensor_wr_0_bits_data_0_18; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_19 = io_tensor_wr_0_bits_data_0_19; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_20 = io_tensor_wr_0_bits_data_0_20; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_21 = io_tensor_wr_0_bits_data_0_21; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_22 = io_tensor_wr_0_bits_data_0_22; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_23 = io_tensor_wr_0_bits_data_0_23; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_24 = io_tensor_wr_0_bits_data_0_24; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_25 = io_tensor_wr_0_bits_data_0_25; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_26 = io_tensor_wr_0_bits_data_0_26; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_27 = io_tensor_wr_0_bits_data_0_27; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_28 = io_tensor_wr_0_bits_data_0_28; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_29 = io_tensor_wr_0_bits_data_0_29; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_30 = io_tensor_wr_0_bits_data_0_30; // @[TensorStore.scala 60:8]
  assign tensorStore_io_tensor_wr_0_bits_data_0_31 = io_tensor_wr_0_bits_data_0_31; // @[TensorStore.scala 60:8]
endmodule
module Store(
  input          clock,
  input          reset,
  input          io_i_post,
  output         io_o_post,
  output         io_inst_ready,
  input          io_inst_valid,
  input  [127:0] io_inst_bits,
  input  [31:0]  io_out_baddr,
  input          io_vme_wr_cmd_ready,
  output         io_vme_wr_cmd_valid,
  output [31:0]  io_vme_wr_cmd_bits_addr,
  output [3:0]   io_vme_wr_cmd_bits_len,
  input          io_vme_wr_data_ready,
  output         io_vme_wr_data_valid,
  output [63:0]  io_vme_wr_data_bits_data,
  input          io_vme_wr_ack,
  input          io_out_wr_0_valid,
  input  [6:0]   io_out_wr_0_bits_idx,
  input  [7:0]   io_out_wr_0_bits_data_0_0,
  input  [7:0]   io_out_wr_0_bits_data_0_1,
  input  [7:0]   io_out_wr_0_bits_data_0_2,
  input  [7:0]   io_out_wr_0_bits_data_0_3,
  input  [7:0]   io_out_wr_0_bits_data_0_4,
  input  [7:0]   io_out_wr_0_bits_data_0_5,
  input  [7:0]   io_out_wr_0_bits_data_0_6,
  input  [7:0]   io_out_wr_0_bits_data_0_7,
  input  [7:0]   io_out_wr_0_bits_data_0_8,
  input  [7:0]   io_out_wr_0_bits_data_0_9,
  input  [7:0]   io_out_wr_0_bits_data_0_10,
  input  [7:0]   io_out_wr_0_bits_data_0_11,
  input  [7:0]   io_out_wr_0_bits_data_0_12,
  input  [7:0]   io_out_wr_0_bits_data_0_13,
  input  [7:0]   io_out_wr_0_bits_data_0_14,
  input  [7:0]   io_out_wr_0_bits_data_0_15,
  input  [7:0]   io_out_wr_0_bits_data_0_16,
  input  [7:0]   io_out_wr_0_bits_data_0_17,
  input  [7:0]   io_out_wr_0_bits_data_0_18,
  input  [7:0]   io_out_wr_0_bits_data_0_19,
  input  [7:0]   io_out_wr_0_bits_data_0_20,
  input  [7:0]   io_out_wr_0_bits_data_0_21,
  input  [7:0]   io_out_wr_0_bits_data_0_22,
  input  [7:0]   io_out_wr_0_bits_data_0_23,
  input  [7:0]   io_out_wr_0_bits_data_0_24,
  input  [7:0]   io_out_wr_0_bits_data_0_25,
  input  [7:0]   io_out_wr_0_bits_data_0_26,
  input  [7:0]   io_out_wr_0_bits_data_0_27,
  input  [7:0]   io_out_wr_0_bits_data_0_28,
  input  [7:0]   io_out_wr_0_bits_data_0_29,
  input  [7:0]   io_out_wr_0_bits_data_0_30,
  input  [7:0]   io_out_wr_0_bits_data_0_31
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  s_clock; // @[Store.scala 46:17]
  wire  s_reset; // @[Store.scala 46:17]
  wire  s_io_spost; // @[Store.scala 46:17]
  wire  s_io_swait; // @[Store.scala 46:17]
  wire  s_io_sready; // @[Store.scala 46:17]
  wire  inst_q_clock; // @[Store.scala 47:22]
  wire  inst_q_reset; // @[Store.scala 47:22]
  wire  inst_q_io_enq_ready; // @[Store.scala 47:22]
  wire  inst_q_io_enq_valid; // @[Store.scala 47:22]
  wire [127:0] inst_q_io_enq_bits; // @[Store.scala 47:22]
  wire  inst_q_io_deq_ready; // @[Store.scala 47:22]
  wire  inst_q_io_deq_valid; // @[Store.scala 47:22]
  wire [127:0] inst_q_io_deq_bits; // @[Store.scala 47:22]
  wire [127:0] dec_io_inst; // @[Store.scala 49:19]
  wire  dec_io_push_prev; // @[Store.scala 49:19]
  wire  dec_io_pop_prev; // @[Store.scala 49:19]
  wire  dec_io_isStore; // @[Store.scala 49:19]
  wire  dec_io_isSync; // @[Store.scala 49:19]
  wire  tensorStore_clock; // @[Store.scala 52:27]
  wire  tensorStore_reset; // @[Store.scala 52:27]
  wire  tensorStore_io_start; // @[Store.scala 52:27]
  wire  tensorStore_io_done; // @[Store.scala 52:27]
  wire [127:0] tensorStore_io_inst; // @[Store.scala 52:27]
  wire [31:0] tensorStore_io_baddr; // @[Store.scala 52:27]
  wire  tensorStore_io_vme_wr_cmd_ready; // @[Store.scala 52:27]
  wire  tensorStore_io_vme_wr_cmd_valid; // @[Store.scala 52:27]
  wire [31:0] tensorStore_io_vme_wr_cmd_bits_addr; // @[Store.scala 52:27]
  wire [3:0] tensorStore_io_vme_wr_cmd_bits_len; // @[Store.scala 52:27]
  wire  tensorStore_io_vme_wr_data_ready; // @[Store.scala 52:27]
  wire  tensorStore_io_vme_wr_data_valid; // @[Store.scala 52:27]
  wire [63:0] tensorStore_io_vme_wr_data_bits_data; // @[Store.scala 52:27]
  wire  tensorStore_io_vme_wr_ack; // @[Store.scala 52:27]
  wire  tensorStore_io_tensor_wr_0_valid; // @[Store.scala 52:27]
  wire [6:0] tensorStore_io_tensor_wr_0_bits_idx; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_0; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_1; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_2; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_3; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_4; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_5; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_6; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_7; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_8; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_9; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_10; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_11; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_12; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_13; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_14; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_15; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_16; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_17; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_18; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_19; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_20; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_21; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_22; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_23; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_24; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_25; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_26; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_27; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_28; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_29; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_30; // @[Store.scala 52:27]
  wire [7:0] tensorStore_io_tensor_wr_0_bits_data_0_31; // @[Store.scala 52:27]
  reg [1:0] state; // @[Store.scala 44:22]
  wire  _start_T = dec_io_pop_prev ? s_io_sready : 1'h1; // @[Store.scala 54:40]
  wire  start = inst_q_io_deq_valid & _start_T; // @[Store.scala 54:35]
  wire [1:0] _GEN_0 = dec_io_isStore ? 2'h2 : state; // @[Store.scala 63:36 64:17 44:22]
  wire [1:0] _GEN_3 = tensorStore_io_done ? 2'h0 : state; // @[Store.scala 72:18 73:15 44:22]
  wire  _inst_q_io_deq_ready_T_3 = state == 2'h2 & tensorStore_io_done | state == 2'h1; // @[Store.scala 80:50]
  wire  _tensorStore_io_start_T_1 = state == 2'h0 & start; // @[Store.scala 83:43]
  Semaphore s ( // @[Store.scala 46:17]
    .clock(s_clock),
    .reset(s_reset),
    .io_spost(s_io_spost),
    .io_swait(s_io_swait),
    .io_sready(s_io_sready)
  );
  Queue_6 inst_q ( // @[Store.scala 47:22]
    .clock(inst_q_clock),
    .reset(inst_q_reset),
    .io_enq_ready(inst_q_io_enq_ready),
    .io_enq_valid(inst_q_io_enq_valid),
    .io_enq_bits(inst_q_io_enq_bits),
    .io_deq_ready(inst_q_io_deq_ready),
    .io_deq_valid(inst_q_io_deq_valid),
    .io_deq_bits(inst_q_io_deq_bits)
  );
  StoreDecode dec ( // @[Store.scala 49:19]
    .io_inst(dec_io_inst),
    .io_push_prev(dec_io_push_prev),
    .io_pop_prev(dec_io_pop_prev),
    .io_isStore(dec_io_isStore),
    .io_isSync(dec_io_isSync)
  );
  TensorStoreOut tensorStore ( // @[Store.scala 52:27]
    .clock(tensorStore_clock),
    .reset(tensorStore_reset),
    .io_start(tensorStore_io_start),
    .io_done(tensorStore_io_done),
    .io_inst(tensorStore_io_inst),
    .io_baddr(tensorStore_io_baddr),
    .io_vme_wr_cmd_ready(tensorStore_io_vme_wr_cmd_ready),
    .io_vme_wr_cmd_valid(tensorStore_io_vme_wr_cmd_valid),
    .io_vme_wr_cmd_bits_addr(tensorStore_io_vme_wr_cmd_bits_addr),
    .io_vme_wr_cmd_bits_len(tensorStore_io_vme_wr_cmd_bits_len),
    .io_vme_wr_data_ready(tensorStore_io_vme_wr_data_ready),
    .io_vme_wr_data_valid(tensorStore_io_vme_wr_data_valid),
    .io_vme_wr_data_bits_data(tensorStore_io_vme_wr_data_bits_data),
    .io_vme_wr_ack(tensorStore_io_vme_wr_ack),
    .io_tensor_wr_0_valid(tensorStore_io_tensor_wr_0_valid),
    .io_tensor_wr_0_bits_idx(tensorStore_io_tensor_wr_0_bits_idx),
    .io_tensor_wr_0_bits_data_0_0(tensorStore_io_tensor_wr_0_bits_data_0_0),
    .io_tensor_wr_0_bits_data_0_1(tensorStore_io_tensor_wr_0_bits_data_0_1),
    .io_tensor_wr_0_bits_data_0_2(tensorStore_io_tensor_wr_0_bits_data_0_2),
    .io_tensor_wr_0_bits_data_0_3(tensorStore_io_tensor_wr_0_bits_data_0_3),
    .io_tensor_wr_0_bits_data_0_4(tensorStore_io_tensor_wr_0_bits_data_0_4),
    .io_tensor_wr_0_bits_data_0_5(tensorStore_io_tensor_wr_0_bits_data_0_5),
    .io_tensor_wr_0_bits_data_0_6(tensorStore_io_tensor_wr_0_bits_data_0_6),
    .io_tensor_wr_0_bits_data_0_7(tensorStore_io_tensor_wr_0_bits_data_0_7),
    .io_tensor_wr_0_bits_data_0_8(tensorStore_io_tensor_wr_0_bits_data_0_8),
    .io_tensor_wr_0_bits_data_0_9(tensorStore_io_tensor_wr_0_bits_data_0_9),
    .io_tensor_wr_0_bits_data_0_10(tensorStore_io_tensor_wr_0_bits_data_0_10),
    .io_tensor_wr_0_bits_data_0_11(tensorStore_io_tensor_wr_0_bits_data_0_11),
    .io_tensor_wr_0_bits_data_0_12(tensorStore_io_tensor_wr_0_bits_data_0_12),
    .io_tensor_wr_0_bits_data_0_13(tensorStore_io_tensor_wr_0_bits_data_0_13),
    .io_tensor_wr_0_bits_data_0_14(tensorStore_io_tensor_wr_0_bits_data_0_14),
    .io_tensor_wr_0_bits_data_0_15(tensorStore_io_tensor_wr_0_bits_data_0_15),
    .io_tensor_wr_0_bits_data_0_16(tensorStore_io_tensor_wr_0_bits_data_0_16),
    .io_tensor_wr_0_bits_data_0_17(tensorStore_io_tensor_wr_0_bits_data_0_17),
    .io_tensor_wr_0_bits_data_0_18(tensorStore_io_tensor_wr_0_bits_data_0_18),
    .io_tensor_wr_0_bits_data_0_19(tensorStore_io_tensor_wr_0_bits_data_0_19),
    .io_tensor_wr_0_bits_data_0_20(tensorStore_io_tensor_wr_0_bits_data_0_20),
    .io_tensor_wr_0_bits_data_0_21(tensorStore_io_tensor_wr_0_bits_data_0_21),
    .io_tensor_wr_0_bits_data_0_22(tensorStore_io_tensor_wr_0_bits_data_0_22),
    .io_tensor_wr_0_bits_data_0_23(tensorStore_io_tensor_wr_0_bits_data_0_23),
    .io_tensor_wr_0_bits_data_0_24(tensorStore_io_tensor_wr_0_bits_data_0_24),
    .io_tensor_wr_0_bits_data_0_25(tensorStore_io_tensor_wr_0_bits_data_0_25),
    .io_tensor_wr_0_bits_data_0_26(tensorStore_io_tensor_wr_0_bits_data_0_26),
    .io_tensor_wr_0_bits_data_0_27(tensorStore_io_tensor_wr_0_bits_data_0_27),
    .io_tensor_wr_0_bits_data_0_28(tensorStore_io_tensor_wr_0_bits_data_0_28),
    .io_tensor_wr_0_bits_data_0_29(tensorStore_io_tensor_wr_0_bits_data_0_29),
    .io_tensor_wr_0_bits_data_0_30(tensorStore_io_tensor_wr_0_bits_data_0_30),
    .io_tensor_wr_0_bits_data_0_31(tensorStore_io_tensor_wr_0_bits_data_0_31)
  );
  assign io_o_post = dec_io_push_prev & _inst_q_io_deq_ready_T_3; // @[Store.scala 92:33]
  assign io_inst_ready = inst_q_io_enq_ready; // @[Store.scala 79:17]
  assign io_vme_wr_cmd_valid = tensorStore_io_vme_wr_cmd_valid; // @[Store.scala 86:13]
  assign io_vme_wr_cmd_bits_addr = tensorStore_io_vme_wr_cmd_bits_addr; // @[Store.scala 86:13]
  assign io_vme_wr_cmd_bits_len = tensorStore_io_vme_wr_cmd_bits_len; // @[Store.scala 86:13]
  assign io_vme_wr_data_valid = tensorStore_io_vme_wr_data_valid; // @[Store.scala 86:13]
  assign io_vme_wr_data_bits_data = tensorStore_io_vme_wr_data_bits_data; // @[Store.scala 86:13]
  assign s_clock = clock;
  assign s_reset = reset;
  assign s_io_spost = io_i_post; // @[Store.scala 90:14]
  assign s_io_swait = dec_io_pop_prev & _tensorStore_io_start_T_1; // @[Store.scala 91:33]
  assign inst_q_clock = clock;
  assign inst_q_reset = reset;
  assign inst_q_io_enq_valid = io_inst_valid; // @[Store.scala 79:17]
  assign inst_q_io_enq_bits = io_inst_bits; // @[Store.scala 79:17]
  assign inst_q_io_deq_ready = state == 2'h2 & tensorStore_io_done | state == 2'h1; // @[Store.scala 80:50]
  assign dec_io_inst = inst_q_io_deq_bits; // @[Store.scala 50:15]
  assign tensorStore_clock = clock;
  assign tensorStore_reset = reset;
  assign tensorStore_io_start = state == 2'h0 & start & dec_io_isStore; // @[Store.scala 83:51]
  assign tensorStore_io_inst = inst_q_io_deq_bits; // @[Store.scala 84:23]
  assign tensorStore_io_baddr = io_out_baddr; // @[Store.scala 85:24]
  assign tensorStore_io_vme_wr_cmd_ready = io_vme_wr_cmd_ready; // @[Store.scala 86:13]
  assign tensorStore_io_vme_wr_data_ready = io_vme_wr_data_ready; // @[Store.scala 86:13]
  assign tensorStore_io_vme_wr_ack = io_vme_wr_ack; // @[Store.scala 86:13]
  assign tensorStore_io_tensor_wr_0_valid = io_out_wr_0_valid; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_idx = io_out_wr_0_bits_idx; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_0 = io_out_wr_0_bits_data_0_0; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_1 = io_out_wr_0_bits_data_0_1; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_2 = io_out_wr_0_bits_data_0_2; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_3 = io_out_wr_0_bits_data_0_3; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_4 = io_out_wr_0_bits_data_0_4; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_5 = io_out_wr_0_bits_data_0_5; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_6 = io_out_wr_0_bits_data_0_6; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_7 = io_out_wr_0_bits_data_0_7; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_8 = io_out_wr_0_bits_data_0_8; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_9 = io_out_wr_0_bits_data_0_9; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_10 = io_out_wr_0_bits_data_0_10; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_11 = io_out_wr_0_bits_data_0_11; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_12 = io_out_wr_0_bits_data_0_12; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_13 = io_out_wr_0_bits_data_0_13; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_14 = io_out_wr_0_bits_data_0_14; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_15 = io_out_wr_0_bits_data_0_15; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_16 = io_out_wr_0_bits_data_0_16; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_17 = io_out_wr_0_bits_data_0_17; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_18 = io_out_wr_0_bits_data_0_18; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_19 = io_out_wr_0_bits_data_0_19; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_20 = io_out_wr_0_bits_data_0_20; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_21 = io_out_wr_0_bits_data_0_21; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_22 = io_out_wr_0_bits_data_0_22; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_23 = io_out_wr_0_bits_data_0_23; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_24 = io_out_wr_0_bits_data_0_24; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_25 = io_out_wr_0_bits_data_0_25; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_26 = io_out_wr_0_bits_data_0_26; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_27 = io_out_wr_0_bits_data_0_27; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_28 = io_out_wr_0_bits_data_0_28; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_29 = io_out_wr_0_bits_data_0_29; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_30 = io_out_wr_0_bits_data_0_30; // @[Store.scala 87:25]
  assign tensorStore_io_tensor_wr_0_bits_data_0_31 = io_out_wr_0_bits_data_0_31; // @[Store.scala 87:25]
  always @(posedge clock) begin
    if (reset) begin // @[Store.scala 44:22]
      state <= 2'h0; // @[Store.scala 44:22]
    end else if (2'h0 == state) begin // @[Store.scala 58:17]
      if (start) begin // @[Store.scala 60:19]
        if (dec_io_isSync) begin // @[Store.scala 61:29]
          state <= 2'h1; // @[Store.scala 62:17]
        end else begin
          state <= _GEN_0;
        end
      end
    end else if (2'h1 == state) begin // @[Store.scala 58:17]
      state <= 2'h0; // @[Store.scala 69:13]
    end else if (2'h2 == state) begin // @[Store.scala 58:17]
      state <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module EventCounters(
  input         clock,
  input         reset,
  input         io_launch,
  input         io_finish,
  output        io_ecnt_0_valid,
  output [31:0] io_ecnt_0_bits,
  output        io_ucnt_0_valid,
  output [31:0] io_ucnt_0_bits,
  input         io_acc_wr_event
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] cycle_cnt; // @[EventCounters.scala 50:26]
  wire [31:0] _cycle_cnt_T_1 = cycle_cnt + 32'h1; // @[EventCounters.scala 52:28]
  reg [31:0] acc_wr_count; // @[EventCounters.scala 59:25]
  wire [31:0] _acc_wr_count_T_1 = acc_wr_count + 32'h1; // @[EventCounters.scala 63:34]
  assign io_ecnt_0_valid = io_finish; // @[EventCounters.scala 56:20]
  assign io_ecnt_0_bits = cycle_cnt; // @[EventCounters.scala 57:19]
  assign io_ucnt_0_valid = io_finish; // @[EventCounters.scala 65:20]
  assign io_ucnt_0_bits = acc_wr_count; // @[EventCounters.scala 66:19]
  always @(posedge clock) begin
    if (reset) begin // @[EventCounters.scala 50:26]
      cycle_cnt <= 32'h0; // @[EventCounters.scala 50:26]
    end else if (io_launch & ~io_finish) begin // @[EventCounters.scala 51:33]
      cycle_cnt <= _cycle_cnt_T_1; // @[EventCounters.scala 52:15]
    end else begin
      cycle_cnt <= 32'h0; // @[EventCounters.scala 54:15]
    end
    if (~io_launch | io_finish) begin // @[EventCounters.scala 60:34]
      acc_wr_count <= 32'h0; // @[EventCounters.scala 61:18]
    end else if (io_acc_wr_event) begin // @[EventCounters.scala 62:32]
      acc_wr_count <= _acc_wr_count_T_1; // @[EventCounters.scala 63:18]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cycle_cnt = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  acc_wr_count = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Core(
  input         clock,
  input         reset,
  input         io_vcr_launch,
  output        io_vcr_finish,
  output        io_vcr_ecnt_0_valid,
  output [31:0] io_vcr_ecnt_0_bits,
  input  [31:0] io_vcr_vals_0,
  input  [31:0] io_vcr_ptrs_0,
  input  [31:0] io_vcr_ptrs_1,
  input  [31:0] io_vcr_ptrs_2,
  input  [31:0] io_vcr_ptrs_3,
  input  [31:0] io_vcr_ptrs_4,
  input  [31:0] io_vcr_ptrs_5,
  output        io_vcr_ucnt_0_valid,
  output [31:0] io_vcr_ucnt_0_bits,
  input         io_vme_rd_0_cmd_ready,
  output        io_vme_rd_0_cmd_valid,
  output [31:0] io_vme_rd_0_cmd_bits_addr,
  output [3:0]  io_vme_rd_0_cmd_bits_len,
  output        io_vme_rd_0_data_ready,
  input         io_vme_rd_0_data_valid,
  input  [63:0] io_vme_rd_0_data_bits_data,
  input         io_vme_rd_1_cmd_ready,
  output        io_vme_rd_1_cmd_valid,
  output [31:0] io_vme_rd_1_cmd_bits_addr,
  output [3:0]  io_vme_rd_1_cmd_bits_len,
  output [20:0] io_vme_rd_1_cmd_bits_tag,
  input         io_vme_rd_1_data_valid,
  input  [63:0] io_vme_rd_1_data_bits_data,
  input  [20:0] io_vme_rd_1_data_bits_tag,
  input         io_vme_rd_1_data_bits_last,
  input         io_vme_rd_2_cmd_ready,
  output        io_vme_rd_2_cmd_valid,
  output [31:0] io_vme_rd_2_cmd_bits_addr,
  output [3:0]  io_vme_rd_2_cmd_bits_len,
  output [20:0] io_vme_rd_2_cmd_bits_tag,
  input         io_vme_rd_2_data_valid,
  input  [63:0] io_vme_rd_2_data_bits_data,
  input  [20:0] io_vme_rd_2_data_bits_tag,
  input         io_vme_rd_3_cmd_ready,
  output        io_vme_rd_3_cmd_valid,
  output [31:0] io_vme_rd_3_cmd_bits_addr,
  output [3:0]  io_vme_rd_3_cmd_bits_len,
  output [20:0] io_vme_rd_3_cmd_bits_tag,
  input         io_vme_rd_3_data_valid,
  input  [63:0] io_vme_rd_3_data_bits_data,
  input  [20:0] io_vme_rd_3_data_bits_tag,
  input         io_vme_rd_4_cmd_ready,
  output        io_vme_rd_4_cmd_valid,
  output [31:0] io_vme_rd_4_cmd_bits_addr,
  output [3:0]  io_vme_rd_4_cmd_bits_len,
  output [20:0] io_vme_rd_4_cmd_bits_tag,
  input         io_vme_rd_4_data_valid,
  input  [63:0] io_vme_rd_4_data_bits_data,
  input  [20:0] io_vme_rd_4_data_bits_tag,
  input         io_vme_wr_0_cmd_ready,
  output        io_vme_wr_0_cmd_valid,
  output [31:0] io_vme_wr_0_cmd_bits_addr,
  output [3:0]  io_vme_wr_0_cmd_bits_len,
  input         io_vme_wr_0_data_ready,
  output        io_vme_wr_0_data_valid,
  output [63:0] io_vme_wr_0_data_bits_data,
  input         io_vme_wr_0_ack
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  fetch_clock; // @[Core.scala 67:21]
  wire  fetch_reset; // @[Core.scala 67:21]
  wire  fetch_io_launch; // @[Core.scala 67:21]
  wire [31:0] fetch_io_ins_baddr; // @[Core.scala 67:21]
  wire [31:0] fetch_io_ins_count; // @[Core.scala 67:21]
  wire  fetch_io_vme_rd_cmd_ready; // @[Core.scala 67:21]
  wire  fetch_io_vme_rd_cmd_valid; // @[Core.scala 67:21]
  wire [31:0] fetch_io_vme_rd_cmd_bits_addr; // @[Core.scala 67:21]
  wire [3:0] fetch_io_vme_rd_cmd_bits_len; // @[Core.scala 67:21]
  wire  fetch_io_vme_rd_data_ready; // @[Core.scala 67:21]
  wire  fetch_io_vme_rd_data_valid; // @[Core.scala 67:21]
  wire [63:0] fetch_io_vme_rd_data_bits_data; // @[Core.scala 67:21]
  wire  fetch_io_inst_ld_ready; // @[Core.scala 67:21]
  wire  fetch_io_inst_ld_valid; // @[Core.scala 67:21]
  wire [127:0] fetch_io_inst_ld_bits; // @[Core.scala 67:21]
  wire  fetch_io_inst_co_ready; // @[Core.scala 67:21]
  wire  fetch_io_inst_co_valid; // @[Core.scala 67:21]
  wire [127:0] fetch_io_inst_co_bits; // @[Core.scala 67:21]
  wire  fetch_io_inst_st_ready; // @[Core.scala 67:21]
  wire  fetch_io_inst_st_valid; // @[Core.scala 67:21]
  wire [127:0] fetch_io_inst_st_bits; // @[Core.scala 67:21]
  wire  load_clock; // @[Core.scala 68:20]
  wire  load_reset; // @[Core.scala 68:20]
  wire  load_io_i_post; // @[Core.scala 68:20]
  wire  load_io_o_post; // @[Core.scala 68:20]
  wire  load_io_inst_ready; // @[Core.scala 68:20]
  wire  load_io_inst_valid; // @[Core.scala 68:20]
  wire [127:0] load_io_inst_bits; // @[Core.scala 68:20]
  wire [31:0] load_io_inp_baddr; // @[Core.scala 68:20]
  wire [31:0] load_io_wgt_baddr; // @[Core.scala 68:20]
  wire  load_io_vme_rd_0_cmd_ready; // @[Core.scala 68:20]
  wire  load_io_vme_rd_0_cmd_valid; // @[Core.scala 68:20]
  wire [31:0] load_io_vme_rd_0_cmd_bits_addr; // @[Core.scala 68:20]
  wire [3:0] load_io_vme_rd_0_cmd_bits_len; // @[Core.scala 68:20]
  wire [20:0] load_io_vme_rd_0_cmd_bits_tag; // @[Core.scala 68:20]
  wire  load_io_vme_rd_0_data_valid; // @[Core.scala 68:20]
  wire [63:0] load_io_vme_rd_0_data_bits_data; // @[Core.scala 68:20]
  wire [20:0] load_io_vme_rd_0_data_bits_tag; // @[Core.scala 68:20]
  wire  load_io_vme_rd_1_cmd_ready; // @[Core.scala 68:20]
  wire  load_io_vme_rd_1_cmd_valid; // @[Core.scala 68:20]
  wire [31:0] load_io_vme_rd_1_cmd_bits_addr; // @[Core.scala 68:20]
  wire [3:0] load_io_vme_rd_1_cmd_bits_len; // @[Core.scala 68:20]
  wire [20:0] load_io_vme_rd_1_cmd_bits_tag; // @[Core.scala 68:20]
  wire  load_io_vme_rd_1_data_valid; // @[Core.scala 68:20]
  wire [63:0] load_io_vme_rd_1_data_bits_data; // @[Core.scala 68:20]
  wire [20:0] load_io_vme_rd_1_data_bits_tag; // @[Core.scala 68:20]
  wire  load_io_inp_rd_0_idx_valid; // @[Core.scala 68:20]
  wire [6:0] load_io_inp_rd_0_idx_bits; // @[Core.scala 68:20]
  wire  load_io_inp_rd_0_data_valid; // @[Core.scala 68:20]
  wire [7:0] load_io_inp_rd_0_data_bits_0_0; // @[Core.scala 68:20]
  wire [7:0] load_io_inp_rd_0_data_bits_0_1; // @[Core.scala 68:20]
  wire [7:0] load_io_inp_rd_0_data_bits_0_2; // @[Core.scala 68:20]
  wire [7:0] load_io_inp_rd_0_data_bits_0_3; // @[Core.scala 68:20]
  wire [7:0] load_io_inp_rd_0_data_bits_0_4; // @[Core.scala 68:20]
  wire [7:0] load_io_inp_rd_0_data_bits_0_5; // @[Core.scala 68:20]
  wire [7:0] load_io_inp_rd_0_data_bits_0_6; // @[Core.scala 68:20]
  wire [7:0] load_io_inp_rd_0_data_bits_0_7; // @[Core.scala 68:20]
  wire [7:0] load_io_inp_rd_0_data_bits_0_8; // @[Core.scala 68:20]
  wire [7:0] load_io_inp_rd_0_data_bits_0_9; // @[Core.scala 68:20]
  wire [7:0] load_io_inp_rd_0_data_bits_0_10; // @[Core.scala 68:20]
  wire [7:0] load_io_inp_rd_0_data_bits_0_11; // @[Core.scala 68:20]
  wire [7:0] load_io_inp_rd_0_data_bits_0_12; // @[Core.scala 68:20]
  wire [7:0] load_io_inp_rd_0_data_bits_0_13; // @[Core.scala 68:20]
  wire [7:0] load_io_inp_rd_0_data_bits_0_14; // @[Core.scala 68:20]
  wire [7:0] load_io_inp_rd_0_data_bits_0_15; // @[Core.scala 68:20]
  wire  load_io_wgt_rd_0_idx_valid; // @[Core.scala 68:20]
  wire [5:0] load_io_wgt_rd_0_idx_bits; // @[Core.scala 68:20]
  wire  load_io_wgt_rd_0_data_valid; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_0_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_0_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_0_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_0_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_0_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_0_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_0_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_0_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_0_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_0_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_0_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_0_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_0_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_0_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_0_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_0_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_1_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_1_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_1_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_1_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_1_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_1_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_1_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_1_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_1_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_1_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_1_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_1_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_1_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_1_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_1_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_1_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_2_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_2_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_2_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_2_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_2_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_2_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_2_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_2_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_2_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_2_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_2_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_2_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_2_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_2_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_2_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_2_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_3_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_3_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_3_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_3_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_3_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_3_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_3_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_3_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_3_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_3_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_3_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_3_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_3_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_3_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_3_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_3_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_4_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_4_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_4_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_4_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_4_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_4_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_4_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_4_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_4_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_4_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_4_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_4_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_4_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_4_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_4_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_4_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_5_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_5_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_5_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_5_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_5_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_5_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_5_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_5_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_5_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_5_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_5_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_5_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_5_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_5_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_5_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_5_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_6_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_6_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_6_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_6_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_6_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_6_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_6_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_6_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_6_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_6_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_6_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_6_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_6_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_6_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_6_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_6_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_7_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_7_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_7_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_7_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_7_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_7_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_7_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_7_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_7_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_7_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_7_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_7_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_7_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_7_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_7_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_7_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_8_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_8_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_8_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_8_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_8_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_8_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_8_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_8_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_8_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_8_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_8_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_8_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_8_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_8_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_8_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_8_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_9_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_9_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_9_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_9_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_9_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_9_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_9_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_9_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_9_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_9_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_9_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_9_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_9_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_9_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_9_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_9_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_10_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_10_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_10_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_10_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_10_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_10_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_10_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_10_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_10_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_10_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_10_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_10_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_10_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_10_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_10_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_10_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_11_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_11_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_11_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_11_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_11_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_11_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_11_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_11_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_11_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_11_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_11_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_11_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_11_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_11_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_11_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_11_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_12_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_12_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_12_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_12_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_12_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_12_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_12_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_12_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_12_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_12_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_12_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_12_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_12_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_12_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_12_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_12_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_13_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_13_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_13_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_13_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_13_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_13_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_13_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_13_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_13_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_13_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_13_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_13_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_13_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_13_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_13_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_13_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_14_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_14_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_14_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_14_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_14_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_14_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_14_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_14_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_14_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_14_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_14_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_14_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_14_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_14_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_14_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_14_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_15_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_15_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_15_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_15_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_15_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_15_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_15_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_15_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_15_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_15_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_15_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_15_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_15_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_15_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_15_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_15_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_16_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_16_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_16_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_16_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_16_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_16_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_16_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_16_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_16_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_16_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_16_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_16_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_16_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_16_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_16_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_16_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_17_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_17_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_17_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_17_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_17_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_17_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_17_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_17_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_17_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_17_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_17_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_17_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_17_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_17_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_17_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_17_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_18_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_18_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_18_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_18_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_18_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_18_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_18_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_18_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_18_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_18_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_18_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_18_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_18_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_18_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_18_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_18_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_19_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_19_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_19_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_19_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_19_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_19_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_19_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_19_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_19_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_19_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_19_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_19_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_19_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_19_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_19_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_19_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_20_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_20_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_20_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_20_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_20_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_20_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_20_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_20_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_20_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_20_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_20_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_20_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_20_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_20_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_20_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_20_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_21_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_21_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_21_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_21_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_21_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_21_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_21_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_21_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_21_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_21_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_21_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_21_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_21_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_21_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_21_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_21_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_22_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_22_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_22_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_22_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_22_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_22_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_22_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_22_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_22_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_22_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_22_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_22_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_22_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_22_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_22_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_22_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_23_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_23_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_23_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_23_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_23_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_23_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_23_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_23_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_23_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_23_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_23_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_23_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_23_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_23_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_23_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_23_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_24_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_24_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_24_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_24_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_24_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_24_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_24_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_24_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_24_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_24_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_24_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_24_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_24_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_24_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_24_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_24_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_25_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_25_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_25_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_25_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_25_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_25_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_25_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_25_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_25_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_25_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_25_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_25_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_25_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_25_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_25_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_25_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_26_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_26_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_26_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_26_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_26_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_26_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_26_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_26_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_26_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_26_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_26_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_26_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_26_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_26_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_26_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_26_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_27_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_27_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_27_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_27_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_27_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_27_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_27_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_27_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_27_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_27_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_27_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_27_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_27_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_27_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_27_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_27_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_28_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_28_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_28_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_28_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_28_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_28_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_28_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_28_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_28_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_28_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_28_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_28_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_28_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_28_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_28_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_28_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_29_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_29_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_29_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_29_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_29_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_29_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_29_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_29_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_29_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_29_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_29_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_29_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_29_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_29_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_29_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_29_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_30_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_30_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_30_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_30_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_30_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_30_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_30_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_30_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_30_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_30_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_30_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_30_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_30_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_30_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_30_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_30_15; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_31_0; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_31_1; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_31_2; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_31_3; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_31_4; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_31_5; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_31_6; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_31_7; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_31_8; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_31_9; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_31_10; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_31_11; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_31_12; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_31_13; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_31_14; // @[Core.scala 68:20]
  wire [7:0] load_io_wgt_rd_0_data_bits_31_15; // @[Core.scala 68:20]
  wire  compute_clock; // @[Core.scala 69:23]
  wire  compute_reset; // @[Core.scala 69:23]
  wire  compute_io_i_post_0; // @[Core.scala 69:23]
  wire  compute_io_i_post_1; // @[Core.scala 69:23]
  wire  compute_io_o_post_0; // @[Core.scala 69:23]
  wire  compute_io_o_post_1; // @[Core.scala 69:23]
  wire  compute_io_inst_ready; // @[Core.scala 69:23]
  wire  compute_io_inst_valid; // @[Core.scala 69:23]
  wire [127:0] compute_io_inst_bits; // @[Core.scala 69:23]
  wire [31:0] compute_io_uop_baddr; // @[Core.scala 69:23]
  wire [31:0] compute_io_acc_baddr; // @[Core.scala 69:23]
  wire  compute_io_vme_rd_0_cmd_ready; // @[Core.scala 69:23]
  wire  compute_io_vme_rd_0_cmd_valid; // @[Core.scala 69:23]
  wire [31:0] compute_io_vme_rd_0_cmd_bits_addr; // @[Core.scala 69:23]
  wire [3:0] compute_io_vme_rd_0_cmd_bits_len; // @[Core.scala 69:23]
  wire [20:0] compute_io_vme_rd_0_cmd_bits_tag; // @[Core.scala 69:23]
  wire  compute_io_vme_rd_0_data_valid; // @[Core.scala 69:23]
  wire [63:0] compute_io_vme_rd_0_data_bits_data; // @[Core.scala 69:23]
  wire [20:0] compute_io_vme_rd_0_data_bits_tag; // @[Core.scala 69:23]
  wire  compute_io_vme_rd_0_data_bits_last; // @[Core.scala 69:23]
  wire  compute_io_vme_rd_1_cmd_ready; // @[Core.scala 69:23]
  wire  compute_io_vme_rd_1_cmd_valid; // @[Core.scala 69:23]
  wire [31:0] compute_io_vme_rd_1_cmd_bits_addr; // @[Core.scala 69:23]
  wire [3:0] compute_io_vme_rd_1_cmd_bits_len; // @[Core.scala 69:23]
  wire [20:0] compute_io_vme_rd_1_cmd_bits_tag; // @[Core.scala 69:23]
  wire  compute_io_vme_rd_1_data_valid; // @[Core.scala 69:23]
  wire [63:0] compute_io_vme_rd_1_data_bits_data; // @[Core.scala 69:23]
  wire [20:0] compute_io_vme_rd_1_data_bits_tag; // @[Core.scala 69:23]
  wire  compute_io_inp_rd_0_idx_valid; // @[Core.scala 69:23]
  wire [6:0] compute_io_inp_rd_0_idx_bits; // @[Core.scala 69:23]
  wire  compute_io_inp_rd_0_data_valid; // @[Core.scala 69:23]
  wire [7:0] compute_io_inp_rd_0_data_bits_0_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_inp_rd_0_data_bits_0_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_inp_rd_0_data_bits_0_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_inp_rd_0_data_bits_0_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_inp_rd_0_data_bits_0_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_inp_rd_0_data_bits_0_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_inp_rd_0_data_bits_0_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_inp_rd_0_data_bits_0_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_inp_rd_0_data_bits_0_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_inp_rd_0_data_bits_0_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_inp_rd_0_data_bits_0_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_inp_rd_0_data_bits_0_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_inp_rd_0_data_bits_0_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_inp_rd_0_data_bits_0_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_inp_rd_0_data_bits_0_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_inp_rd_0_data_bits_0_15; // @[Core.scala 69:23]
  wire  compute_io_wgt_rd_0_idx_valid; // @[Core.scala 69:23]
  wire [5:0] compute_io_wgt_rd_0_idx_bits; // @[Core.scala 69:23]
  wire  compute_io_wgt_rd_0_data_valid; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_0_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_0_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_0_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_0_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_0_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_0_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_0_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_0_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_0_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_0_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_0_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_0_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_0_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_0_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_0_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_0_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_1_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_1_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_1_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_1_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_1_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_1_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_1_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_1_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_1_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_1_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_1_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_1_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_1_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_1_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_1_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_1_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_2_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_2_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_2_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_2_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_2_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_2_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_2_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_2_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_2_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_2_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_2_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_2_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_2_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_2_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_2_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_2_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_3_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_3_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_3_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_3_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_3_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_3_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_3_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_3_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_3_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_3_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_3_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_3_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_3_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_3_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_3_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_3_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_4_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_4_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_4_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_4_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_4_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_4_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_4_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_4_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_4_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_4_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_4_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_4_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_4_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_4_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_4_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_4_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_5_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_5_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_5_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_5_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_5_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_5_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_5_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_5_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_5_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_5_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_5_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_5_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_5_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_5_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_5_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_5_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_6_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_6_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_6_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_6_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_6_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_6_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_6_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_6_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_6_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_6_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_6_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_6_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_6_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_6_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_6_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_6_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_7_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_7_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_7_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_7_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_7_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_7_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_7_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_7_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_7_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_7_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_7_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_7_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_7_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_7_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_7_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_7_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_8_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_8_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_8_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_8_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_8_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_8_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_8_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_8_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_8_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_8_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_8_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_8_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_8_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_8_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_8_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_8_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_9_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_9_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_9_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_9_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_9_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_9_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_9_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_9_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_9_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_9_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_9_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_9_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_9_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_9_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_9_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_9_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_10_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_10_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_10_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_10_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_10_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_10_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_10_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_10_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_10_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_10_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_10_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_10_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_10_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_10_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_10_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_10_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_11_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_11_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_11_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_11_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_11_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_11_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_11_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_11_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_11_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_11_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_11_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_11_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_11_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_11_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_11_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_11_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_12_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_12_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_12_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_12_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_12_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_12_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_12_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_12_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_12_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_12_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_12_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_12_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_12_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_12_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_12_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_12_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_13_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_13_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_13_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_13_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_13_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_13_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_13_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_13_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_13_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_13_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_13_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_13_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_13_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_13_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_13_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_13_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_14_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_14_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_14_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_14_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_14_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_14_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_14_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_14_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_14_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_14_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_14_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_14_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_14_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_14_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_14_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_14_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_15_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_15_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_15_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_15_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_15_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_15_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_15_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_15_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_15_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_15_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_15_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_15_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_15_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_15_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_15_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_15_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_16_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_16_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_16_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_16_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_16_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_16_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_16_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_16_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_16_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_16_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_16_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_16_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_16_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_16_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_16_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_16_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_17_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_17_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_17_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_17_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_17_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_17_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_17_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_17_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_17_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_17_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_17_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_17_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_17_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_17_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_17_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_17_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_18_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_18_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_18_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_18_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_18_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_18_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_18_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_18_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_18_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_18_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_18_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_18_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_18_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_18_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_18_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_18_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_19_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_19_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_19_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_19_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_19_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_19_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_19_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_19_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_19_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_19_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_19_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_19_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_19_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_19_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_19_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_19_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_20_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_20_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_20_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_20_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_20_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_20_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_20_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_20_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_20_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_20_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_20_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_20_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_20_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_20_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_20_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_20_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_21_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_21_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_21_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_21_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_21_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_21_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_21_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_21_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_21_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_21_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_21_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_21_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_21_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_21_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_21_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_21_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_22_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_22_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_22_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_22_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_22_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_22_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_22_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_22_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_22_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_22_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_22_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_22_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_22_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_22_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_22_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_22_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_23_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_23_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_23_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_23_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_23_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_23_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_23_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_23_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_23_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_23_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_23_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_23_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_23_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_23_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_23_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_23_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_24_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_24_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_24_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_24_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_24_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_24_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_24_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_24_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_24_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_24_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_24_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_24_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_24_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_24_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_24_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_24_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_25_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_25_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_25_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_25_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_25_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_25_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_25_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_25_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_25_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_25_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_25_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_25_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_25_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_25_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_25_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_25_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_26_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_26_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_26_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_26_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_26_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_26_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_26_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_26_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_26_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_26_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_26_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_26_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_26_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_26_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_26_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_26_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_27_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_27_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_27_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_27_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_27_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_27_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_27_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_27_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_27_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_27_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_27_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_27_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_27_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_27_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_27_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_27_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_28_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_28_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_28_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_28_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_28_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_28_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_28_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_28_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_28_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_28_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_28_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_28_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_28_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_28_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_28_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_28_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_29_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_29_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_29_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_29_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_29_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_29_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_29_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_29_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_29_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_29_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_29_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_29_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_29_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_29_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_29_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_29_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_30_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_30_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_30_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_30_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_30_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_30_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_30_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_30_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_30_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_30_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_30_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_30_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_30_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_30_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_30_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_30_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_31_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_31_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_31_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_31_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_31_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_31_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_31_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_31_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_31_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_31_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_31_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_31_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_31_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_31_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_31_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_wgt_rd_0_data_bits_31_15; // @[Core.scala 69:23]
  wire  compute_io_out_wr_0_valid; // @[Core.scala 69:23]
  wire [6:0] compute_io_out_wr_0_bits_idx; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_0; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_1; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_2; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_3; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_4; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_5; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_6; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_7; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_8; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_9; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_10; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_11; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_12; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_13; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_14; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_15; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_16; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_17; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_18; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_19; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_20; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_21; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_22; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_23; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_24; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_25; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_26; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_27; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_28; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_29; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_30; // @[Core.scala 69:23]
  wire [7:0] compute_io_out_wr_0_bits_data_0_31; // @[Core.scala 69:23]
  wire  compute_io_finish; // @[Core.scala 69:23]
  wire  compute_io_acc_wr_event; // @[Core.scala 69:23]
  wire  store_clock; // @[Core.scala 70:21]
  wire  store_reset; // @[Core.scala 70:21]
  wire  store_io_i_post; // @[Core.scala 70:21]
  wire  store_io_o_post; // @[Core.scala 70:21]
  wire  store_io_inst_ready; // @[Core.scala 70:21]
  wire  store_io_inst_valid; // @[Core.scala 70:21]
  wire [127:0] store_io_inst_bits; // @[Core.scala 70:21]
  wire [31:0] store_io_out_baddr; // @[Core.scala 70:21]
  wire  store_io_vme_wr_cmd_ready; // @[Core.scala 70:21]
  wire  store_io_vme_wr_cmd_valid; // @[Core.scala 70:21]
  wire [31:0] store_io_vme_wr_cmd_bits_addr; // @[Core.scala 70:21]
  wire [3:0] store_io_vme_wr_cmd_bits_len; // @[Core.scala 70:21]
  wire  store_io_vme_wr_data_ready; // @[Core.scala 70:21]
  wire  store_io_vme_wr_data_valid; // @[Core.scala 70:21]
  wire [63:0] store_io_vme_wr_data_bits_data; // @[Core.scala 70:21]
  wire  store_io_vme_wr_ack; // @[Core.scala 70:21]
  wire  store_io_out_wr_0_valid; // @[Core.scala 70:21]
  wire [6:0] store_io_out_wr_0_bits_idx; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_0; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_1; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_2; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_3; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_4; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_5; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_6; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_7; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_8; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_9; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_10; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_11; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_12; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_13; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_14; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_15; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_16; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_17; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_18; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_19; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_20; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_21; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_22; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_23; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_24; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_25; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_26; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_27; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_28; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_29; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_30; // @[Core.scala 70:21]
  wire [7:0] store_io_out_wr_0_bits_data_0_31; // @[Core.scala 70:21]
  wire  ecounters_clock; // @[Core.scala 71:25]
  wire  ecounters_reset; // @[Core.scala 71:25]
  wire  ecounters_io_launch; // @[Core.scala 71:25]
  wire  ecounters_io_finish; // @[Core.scala 71:25]
  wire  ecounters_io_ecnt_0_valid; // @[Core.scala 71:25]
  wire [31:0] ecounters_io_ecnt_0_bits; // @[Core.scala 71:25]
  wire  ecounters_io_ucnt_0_valid; // @[Core.scala 71:25]
  wire [31:0] ecounters_io_ucnt_0_bits; // @[Core.scala 71:25]
  wire  ecounters_io_acc_wr_event; // @[Core.scala 71:25]
  reg  finish; // @[Core.scala 119:23]
  Fetch fetch ( // @[Core.scala 67:21]
    .clock(fetch_clock),
    .reset(fetch_reset),
    .io_launch(fetch_io_launch),
    .io_ins_baddr(fetch_io_ins_baddr),
    .io_ins_count(fetch_io_ins_count),
    .io_vme_rd_cmd_ready(fetch_io_vme_rd_cmd_ready),
    .io_vme_rd_cmd_valid(fetch_io_vme_rd_cmd_valid),
    .io_vme_rd_cmd_bits_addr(fetch_io_vme_rd_cmd_bits_addr),
    .io_vme_rd_cmd_bits_len(fetch_io_vme_rd_cmd_bits_len),
    .io_vme_rd_data_ready(fetch_io_vme_rd_data_ready),
    .io_vme_rd_data_valid(fetch_io_vme_rd_data_valid),
    .io_vme_rd_data_bits_data(fetch_io_vme_rd_data_bits_data),
    .io_inst_ld_ready(fetch_io_inst_ld_ready),
    .io_inst_ld_valid(fetch_io_inst_ld_valid),
    .io_inst_ld_bits(fetch_io_inst_ld_bits),
    .io_inst_co_ready(fetch_io_inst_co_ready),
    .io_inst_co_valid(fetch_io_inst_co_valid),
    .io_inst_co_bits(fetch_io_inst_co_bits),
    .io_inst_st_ready(fetch_io_inst_st_ready),
    .io_inst_st_valid(fetch_io_inst_st_valid),
    .io_inst_st_bits(fetch_io_inst_st_bits)
  );
  Load load ( // @[Core.scala 68:20]
    .clock(load_clock),
    .reset(load_reset),
    .io_i_post(load_io_i_post),
    .io_o_post(load_io_o_post),
    .io_inst_ready(load_io_inst_ready),
    .io_inst_valid(load_io_inst_valid),
    .io_inst_bits(load_io_inst_bits),
    .io_inp_baddr(load_io_inp_baddr),
    .io_wgt_baddr(load_io_wgt_baddr),
    .io_vme_rd_0_cmd_ready(load_io_vme_rd_0_cmd_ready),
    .io_vme_rd_0_cmd_valid(load_io_vme_rd_0_cmd_valid),
    .io_vme_rd_0_cmd_bits_addr(load_io_vme_rd_0_cmd_bits_addr),
    .io_vme_rd_0_cmd_bits_len(load_io_vme_rd_0_cmd_bits_len),
    .io_vme_rd_0_cmd_bits_tag(load_io_vme_rd_0_cmd_bits_tag),
    .io_vme_rd_0_data_valid(load_io_vme_rd_0_data_valid),
    .io_vme_rd_0_data_bits_data(load_io_vme_rd_0_data_bits_data),
    .io_vme_rd_0_data_bits_tag(load_io_vme_rd_0_data_bits_tag),
    .io_vme_rd_1_cmd_ready(load_io_vme_rd_1_cmd_ready),
    .io_vme_rd_1_cmd_valid(load_io_vme_rd_1_cmd_valid),
    .io_vme_rd_1_cmd_bits_addr(load_io_vme_rd_1_cmd_bits_addr),
    .io_vme_rd_1_cmd_bits_len(load_io_vme_rd_1_cmd_bits_len),
    .io_vme_rd_1_cmd_bits_tag(load_io_vme_rd_1_cmd_bits_tag),
    .io_vme_rd_1_data_valid(load_io_vme_rd_1_data_valid),
    .io_vme_rd_1_data_bits_data(load_io_vme_rd_1_data_bits_data),
    .io_vme_rd_1_data_bits_tag(load_io_vme_rd_1_data_bits_tag),
    .io_inp_rd_0_idx_valid(load_io_inp_rd_0_idx_valid),
    .io_inp_rd_0_idx_bits(load_io_inp_rd_0_idx_bits),
    .io_inp_rd_0_data_valid(load_io_inp_rd_0_data_valid),
    .io_inp_rd_0_data_bits_0_0(load_io_inp_rd_0_data_bits_0_0),
    .io_inp_rd_0_data_bits_0_1(load_io_inp_rd_0_data_bits_0_1),
    .io_inp_rd_0_data_bits_0_2(load_io_inp_rd_0_data_bits_0_2),
    .io_inp_rd_0_data_bits_0_3(load_io_inp_rd_0_data_bits_0_3),
    .io_inp_rd_0_data_bits_0_4(load_io_inp_rd_0_data_bits_0_4),
    .io_inp_rd_0_data_bits_0_5(load_io_inp_rd_0_data_bits_0_5),
    .io_inp_rd_0_data_bits_0_6(load_io_inp_rd_0_data_bits_0_6),
    .io_inp_rd_0_data_bits_0_7(load_io_inp_rd_0_data_bits_0_7),
    .io_inp_rd_0_data_bits_0_8(load_io_inp_rd_0_data_bits_0_8),
    .io_inp_rd_0_data_bits_0_9(load_io_inp_rd_0_data_bits_0_9),
    .io_inp_rd_0_data_bits_0_10(load_io_inp_rd_0_data_bits_0_10),
    .io_inp_rd_0_data_bits_0_11(load_io_inp_rd_0_data_bits_0_11),
    .io_inp_rd_0_data_bits_0_12(load_io_inp_rd_0_data_bits_0_12),
    .io_inp_rd_0_data_bits_0_13(load_io_inp_rd_0_data_bits_0_13),
    .io_inp_rd_0_data_bits_0_14(load_io_inp_rd_0_data_bits_0_14),
    .io_inp_rd_0_data_bits_0_15(load_io_inp_rd_0_data_bits_0_15),
    .io_wgt_rd_0_idx_valid(load_io_wgt_rd_0_idx_valid),
    .io_wgt_rd_0_idx_bits(load_io_wgt_rd_0_idx_bits),
    .io_wgt_rd_0_data_valid(load_io_wgt_rd_0_data_valid),
    .io_wgt_rd_0_data_bits_0_0(load_io_wgt_rd_0_data_bits_0_0),
    .io_wgt_rd_0_data_bits_0_1(load_io_wgt_rd_0_data_bits_0_1),
    .io_wgt_rd_0_data_bits_0_2(load_io_wgt_rd_0_data_bits_0_2),
    .io_wgt_rd_0_data_bits_0_3(load_io_wgt_rd_0_data_bits_0_3),
    .io_wgt_rd_0_data_bits_0_4(load_io_wgt_rd_0_data_bits_0_4),
    .io_wgt_rd_0_data_bits_0_5(load_io_wgt_rd_0_data_bits_0_5),
    .io_wgt_rd_0_data_bits_0_6(load_io_wgt_rd_0_data_bits_0_6),
    .io_wgt_rd_0_data_bits_0_7(load_io_wgt_rd_0_data_bits_0_7),
    .io_wgt_rd_0_data_bits_0_8(load_io_wgt_rd_0_data_bits_0_8),
    .io_wgt_rd_0_data_bits_0_9(load_io_wgt_rd_0_data_bits_0_9),
    .io_wgt_rd_0_data_bits_0_10(load_io_wgt_rd_0_data_bits_0_10),
    .io_wgt_rd_0_data_bits_0_11(load_io_wgt_rd_0_data_bits_0_11),
    .io_wgt_rd_0_data_bits_0_12(load_io_wgt_rd_0_data_bits_0_12),
    .io_wgt_rd_0_data_bits_0_13(load_io_wgt_rd_0_data_bits_0_13),
    .io_wgt_rd_0_data_bits_0_14(load_io_wgt_rd_0_data_bits_0_14),
    .io_wgt_rd_0_data_bits_0_15(load_io_wgt_rd_0_data_bits_0_15),
    .io_wgt_rd_0_data_bits_1_0(load_io_wgt_rd_0_data_bits_1_0),
    .io_wgt_rd_0_data_bits_1_1(load_io_wgt_rd_0_data_bits_1_1),
    .io_wgt_rd_0_data_bits_1_2(load_io_wgt_rd_0_data_bits_1_2),
    .io_wgt_rd_0_data_bits_1_3(load_io_wgt_rd_0_data_bits_1_3),
    .io_wgt_rd_0_data_bits_1_4(load_io_wgt_rd_0_data_bits_1_4),
    .io_wgt_rd_0_data_bits_1_5(load_io_wgt_rd_0_data_bits_1_5),
    .io_wgt_rd_0_data_bits_1_6(load_io_wgt_rd_0_data_bits_1_6),
    .io_wgt_rd_0_data_bits_1_7(load_io_wgt_rd_0_data_bits_1_7),
    .io_wgt_rd_0_data_bits_1_8(load_io_wgt_rd_0_data_bits_1_8),
    .io_wgt_rd_0_data_bits_1_9(load_io_wgt_rd_0_data_bits_1_9),
    .io_wgt_rd_0_data_bits_1_10(load_io_wgt_rd_0_data_bits_1_10),
    .io_wgt_rd_0_data_bits_1_11(load_io_wgt_rd_0_data_bits_1_11),
    .io_wgt_rd_0_data_bits_1_12(load_io_wgt_rd_0_data_bits_1_12),
    .io_wgt_rd_0_data_bits_1_13(load_io_wgt_rd_0_data_bits_1_13),
    .io_wgt_rd_0_data_bits_1_14(load_io_wgt_rd_0_data_bits_1_14),
    .io_wgt_rd_0_data_bits_1_15(load_io_wgt_rd_0_data_bits_1_15),
    .io_wgt_rd_0_data_bits_2_0(load_io_wgt_rd_0_data_bits_2_0),
    .io_wgt_rd_0_data_bits_2_1(load_io_wgt_rd_0_data_bits_2_1),
    .io_wgt_rd_0_data_bits_2_2(load_io_wgt_rd_0_data_bits_2_2),
    .io_wgt_rd_0_data_bits_2_3(load_io_wgt_rd_0_data_bits_2_3),
    .io_wgt_rd_0_data_bits_2_4(load_io_wgt_rd_0_data_bits_2_4),
    .io_wgt_rd_0_data_bits_2_5(load_io_wgt_rd_0_data_bits_2_5),
    .io_wgt_rd_0_data_bits_2_6(load_io_wgt_rd_0_data_bits_2_6),
    .io_wgt_rd_0_data_bits_2_7(load_io_wgt_rd_0_data_bits_2_7),
    .io_wgt_rd_0_data_bits_2_8(load_io_wgt_rd_0_data_bits_2_8),
    .io_wgt_rd_0_data_bits_2_9(load_io_wgt_rd_0_data_bits_2_9),
    .io_wgt_rd_0_data_bits_2_10(load_io_wgt_rd_0_data_bits_2_10),
    .io_wgt_rd_0_data_bits_2_11(load_io_wgt_rd_0_data_bits_2_11),
    .io_wgt_rd_0_data_bits_2_12(load_io_wgt_rd_0_data_bits_2_12),
    .io_wgt_rd_0_data_bits_2_13(load_io_wgt_rd_0_data_bits_2_13),
    .io_wgt_rd_0_data_bits_2_14(load_io_wgt_rd_0_data_bits_2_14),
    .io_wgt_rd_0_data_bits_2_15(load_io_wgt_rd_0_data_bits_2_15),
    .io_wgt_rd_0_data_bits_3_0(load_io_wgt_rd_0_data_bits_3_0),
    .io_wgt_rd_0_data_bits_3_1(load_io_wgt_rd_0_data_bits_3_1),
    .io_wgt_rd_0_data_bits_3_2(load_io_wgt_rd_0_data_bits_3_2),
    .io_wgt_rd_0_data_bits_3_3(load_io_wgt_rd_0_data_bits_3_3),
    .io_wgt_rd_0_data_bits_3_4(load_io_wgt_rd_0_data_bits_3_4),
    .io_wgt_rd_0_data_bits_3_5(load_io_wgt_rd_0_data_bits_3_5),
    .io_wgt_rd_0_data_bits_3_6(load_io_wgt_rd_0_data_bits_3_6),
    .io_wgt_rd_0_data_bits_3_7(load_io_wgt_rd_0_data_bits_3_7),
    .io_wgt_rd_0_data_bits_3_8(load_io_wgt_rd_0_data_bits_3_8),
    .io_wgt_rd_0_data_bits_3_9(load_io_wgt_rd_0_data_bits_3_9),
    .io_wgt_rd_0_data_bits_3_10(load_io_wgt_rd_0_data_bits_3_10),
    .io_wgt_rd_0_data_bits_3_11(load_io_wgt_rd_0_data_bits_3_11),
    .io_wgt_rd_0_data_bits_3_12(load_io_wgt_rd_0_data_bits_3_12),
    .io_wgt_rd_0_data_bits_3_13(load_io_wgt_rd_0_data_bits_3_13),
    .io_wgt_rd_0_data_bits_3_14(load_io_wgt_rd_0_data_bits_3_14),
    .io_wgt_rd_0_data_bits_3_15(load_io_wgt_rd_0_data_bits_3_15),
    .io_wgt_rd_0_data_bits_4_0(load_io_wgt_rd_0_data_bits_4_0),
    .io_wgt_rd_0_data_bits_4_1(load_io_wgt_rd_0_data_bits_4_1),
    .io_wgt_rd_0_data_bits_4_2(load_io_wgt_rd_0_data_bits_4_2),
    .io_wgt_rd_0_data_bits_4_3(load_io_wgt_rd_0_data_bits_4_3),
    .io_wgt_rd_0_data_bits_4_4(load_io_wgt_rd_0_data_bits_4_4),
    .io_wgt_rd_0_data_bits_4_5(load_io_wgt_rd_0_data_bits_4_5),
    .io_wgt_rd_0_data_bits_4_6(load_io_wgt_rd_0_data_bits_4_6),
    .io_wgt_rd_0_data_bits_4_7(load_io_wgt_rd_0_data_bits_4_7),
    .io_wgt_rd_0_data_bits_4_8(load_io_wgt_rd_0_data_bits_4_8),
    .io_wgt_rd_0_data_bits_4_9(load_io_wgt_rd_0_data_bits_4_9),
    .io_wgt_rd_0_data_bits_4_10(load_io_wgt_rd_0_data_bits_4_10),
    .io_wgt_rd_0_data_bits_4_11(load_io_wgt_rd_0_data_bits_4_11),
    .io_wgt_rd_0_data_bits_4_12(load_io_wgt_rd_0_data_bits_4_12),
    .io_wgt_rd_0_data_bits_4_13(load_io_wgt_rd_0_data_bits_4_13),
    .io_wgt_rd_0_data_bits_4_14(load_io_wgt_rd_0_data_bits_4_14),
    .io_wgt_rd_0_data_bits_4_15(load_io_wgt_rd_0_data_bits_4_15),
    .io_wgt_rd_0_data_bits_5_0(load_io_wgt_rd_0_data_bits_5_0),
    .io_wgt_rd_0_data_bits_5_1(load_io_wgt_rd_0_data_bits_5_1),
    .io_wgt_rd_0_data_bits_5_2(load_io_wgt_rd_0_data_bits_5_2),
    .io_wgt_rd_0_data_bits_5_3(load_io_wgt_rd_0_data_bits_5_3),
    .io_wgt_rd_0_data_bits_5_4(load_io_wgt_rd_0_data_bits_5_4),
    .io_wgt_rd_0_data_bits_5_5(load_io_wgt_rd_0_data_bits_5_5),
    .io_wgt_rd_0_data_bits_5_6(load_io_wgt_rd_0_data_bits_5_6),
    .io_wgt_rd_0_data_bits_5_7(load_io_wgt_rd_0_data_bits_5_7),
    .io_wgt_rd_0_data_bits_5_8(load_io_wgt_rd_0_data_bits_5_8),
    .io_wgt_rd_0_data_bits_5_9(load_io_wgt_rd_0_data_bits_5_9),
    .io_wgt_rd_0_data_bits_5_10(load_io_wgt_rd_0_data_bits_5_10),
    .io_wgt_rd_0_data_bits_5_11(load_io_wgt_rd_0_data_bits_5_11),
    .io_wgt_rd_0_data_bits_5_12(load_io_wgt_rd_0_data_bits_5_12),
    .io_wgt_rd_0_data_bits_5_13(load_io_wgt_rd_0_data_bits_5_13),
    .io_wgt_rd_0_data_bits_5_14(load_io_wgt_rd_0_data_bits_5_14),
    .io_wgt_rd_0_data_bits_5_15(load_io_wgt_rd_0_data_bits_5_15),
    .io_wgt_rd_0_data_bits_6_0(load_io_wgt_rd_0_data_bits_6_0),
    .io_wgt_rd_0_data_bits_6_1(load_io_wgt_rd_0_data_bits_6_1),
    .io_wgt_rd_0_data_bits_6_2(load_io_wgt_rd_0_data_bits_6_2),
    .io_wgt_rd_0_data_bits_6_3(load_io_wgt_rd_0_data_bits_6_3),
    .io_wgt_rd_0_data_bits_6_4(load_io_wgt_rd_0_data_bits_6_4),
    .io_wgt_rd_0_data_bits_6_5(load_io_wgt_rd_0_data_bits_6_5),
    .io_wgt_rd_0_data_bits_6_6(load_io_wgt_rd_0_data_bits_6_6),
    .io_wgt_rd_0_data_bits_6_7(load_io_wgt_rd_0_data_bits_6_7),
    .io_wgt_rd_0_data_bits_6_8(load_io_wgt_rd_0_data_bits_6_8),
    .io_wgt_rd_0_data_bits_6_9(load_io_wgt_rd_0_data_bits_6_9),
    .io_wgt_rd_0_data_bits_6_10(load_io_wgt_rd_0_data_bits_6_10),
    .io_wgt_rd_0_data_bits_6_11(load_io_wgt_rd_0_data_bits_6_11),
    .io_wgt_rd_0_data_bits_6_12(load_io_wgt_rd_0_data_bits_6_12),
    .io_wgt_rd_0_data_bits_6_13(load_io_wgt_rd_0_data_bits_6_13),
    .io_wgt_rd_0_data_bits_6_14(load_io_wgt_rd_0_data_bits_6_14),
    .io_wgt_rd_0_data_bits_6_15(load_io_wgt_rd_0_data_bits_6_15),
    .io_wgt_rd_0_data_bits_7_0(load_io_wgt_rd_0_data_bits_7_0),
    .io_wgt_rd_0_data_bits_7_1(load_io_wgt_rd_0_data_bits_7_1),
    .io_wgt_rd_0_data_bits_7_2(load_io_wgt_rd_0_data_bits_7_2),
    .io_wgt_rd_0_data_bits_7_3(load_io_wgt_rd_0_data_bits_7_3),
    .io_wgt_rd_0_data_bits_7_4(load_io_wgt_rd_0_data_bits_7_4),
    .io_wgt_rd_0_data_bits_7_5(load_io_wgt_rd_0_data_bits_7_5),
    .io_wgt_rd_0_data_bits_7_6(load_io_wgt_rd_0_data_bits_7_6),
    .io_wgt_rd_0_data_bits_7_7(load_io_wgt_rd_0_data_bits_7_7),
    .io_wgt_rd_0_data_bits_7_8(load_io_wgt_rd_0_data_bits_7_8),
    .io_wgt_rd_0_data_bits_7_9(load_io_wgt_rd_0_data_bits_7_9),
    .io_wgt_rd_0_data_bits_7_10(load_io_wgt_rd_0_data_bits_7_10),
    .io_wgt_rd_0_data_bits_7_11(load_io_wgt_rd_0_data_bits_7_11),
    .io_wgt_rd_0_data_bits_7_12(load_io_wgt_rd_0_data_bits_7_12),
    .io_wgt_rd_0_data_bits_7_13(load_io_wgt_rd_0_data_bits_7_13),
    .io_wgt_rd_0_data_bits_7_14(load_io_wgt_rd_0_data_bits_7_14),
    .io_wgt_rd_0_data_bits_7_15(load_io_wgt_rd_0_data_bits_7_15),
    .io_wgt_rd_0_data_bits_8_0(load_io_wgt_rd_0_data_bits_8_0),
    .io_wgt_rd_0_data_bits_8_1(load_io_wgt_rd_0_data_bits_8_1),
    .io_wgt_rd_0_data_bits_8_2(load_io_wgt_rd_0_data_bits_8_2),
    .io_wgt_rd_0_data_bits_8_3(load_io_wgt_rd_0_data_bits_8_3),
    .io_wgt_rd_0_data_bits_8_4(load_io_wgt_rd_0_data_bits_8_4),
    .io_wgt_rd_0_data_bits_8_5(load_io_wgt_rd_0_data_bits_8_5),
    .io_wgt_rd_0_data_bits_8_6(load_io_wgt_rd_0_data_bits_8_6),
    .io_wgt_rd_0_data_bits_8_7(load_io_wgt_rd_0_data_bits_8_7),
    .io_wgt_rd_0_data_bits_8_8(load_io_wgt_rd_0_data_bits_8_8),
    .io_wgt_rd_0_data_bits_8_9(load_io_wgt_rd_0_data_bits_8_9),
    .io_wgt_rd_0_data_bits_8_10(load_io_wgt_rd_0_data_bits_8_10),
    .io_wgt_rd_0_data_bits_8_11(load_io_wgt_rd_0_data_bits_8_11),
    .io_wgt_rd_0_data_bits_8_12(load_io_wgt_rd_0_data_bits_8_12),
    .io_wgt_rd_0_data_bits_8_13(load_io_wgt_rd_0_data_bits_8_13),
    .io_wgt_rd_0_data_bits_8_14(load_io_wgt_rd_0_data_bits_8_14),
    .io_wgt_rd_0_data_bits_8_15(load_io_wgt_rd_0_data_bits_8_15),
    .io_wgt_rd_0_data_bits_9_0(load_io_wgt_rd_0_data_bits_9_0),
    .io_wgt_rd_0_data_bits_9_1(load_io_wgt_rd_0_data_bits_9_1),
    .io_wgt_rd_0_data_bits_9_2(load_io_wgt_rd_0_data_bits_9_2),
    .io_wgt_rd_0_data_bits_9_3(load_io_wgt_rd_0_data_bits_9_3),
    .io_wgt_rd_0_data_bits_9_4(load_io_wgt_rd_0_data_bits_9_4),
    .io_wgt_rd_0_data_bits_9_5(load_io_wgt_rd_0_data_bits_9_5),
    .io_wgt_rd_0_data_bits_9_6(load_io_wgt_rd_0_data_bits_9_6),
    .io_wgt_rd_0_data_bits_9_7(load_io_wgt_rd_0_data_bits_9_7),
    .io_wgt_rd_0_data_bits_9_8(load_io_wgt_rd_0_data_bits_9_8),
    .io_wgt_rd_0_data_bits_9_9(load_io_wgt_rd_0_data_bits_9_9),
    .io_wgt_rd_0_data_bits_9_10(load_io_wgt_rd_0_data_bits_9_10),
    .io_wgt_rd_0_data_bits_9_11(load_io_wgt_rd_0_data_bits_9_11),
    .io_wgt_rd_0_data_bits_9_12(load_io_wgt_rd_0_data_bits_9_12),
    .io_wgt_rd_0_data_bits_9_13(load_io_wgt_rd_0_data_bits_9_13),
    .io_wgt_rd_0_data_bits_9_14(load_io_wgt_rd_0_data_bits_9_14),
    .io_wgt_rd_0_data_bits_9_15(load_io_wgt_rd_0_data_bits_9_15),
    .io_wgt_rd_0_data_bits_10_0(load_io_wgt_rd_0_data_bits_10_0),
    .io_wgt_rd_0_data_bits_10_1(load_io_wgt_rd_0_data_bits_10_1),
    .io_wgt_rd_0_data_bits_10_2(load_io_wgt_rd_0_data_bits_10_2),
    .io_wgt_rd_0_data_bits_10_3(load_io_wgt_rd_0_data_bits_10_3),
    .io_wgt_rd_0_data_bits_10_4(load_io_wgt_rd_0_data_bits_10_4),
    .io_wgt_rd_0_data_bits_10_5(load_io_wgt_rd_0_data_bits_10_5),
    .io_wgt_rd_0_data_bits_10_6(load_io_wgt_rd_0_data_bits_10_6),
    .io_wgt_rd_0_data_bits_10_7(load_io_wgt_rd_0_data_bits_10_7),
    .io_wgt_rd_0_data_bits_10_8(load_io_wgt_rd_0_data_bits_10_8),
    .io_wgt_rd_0_data_bits_10_9(load_io_wgt_rd_0_data_bits_10_9),
    .io_wgt_rd_0_data_bits_10_10(load_io_wgt_rd_0_data_bits_10_10),
    .io_wgt_rd_0_data_bits_10_11(load_io_wgt_rd_0_data_bits_10_11),
    .io_wgt_rd_0_data_bits_10_12(load_io_wgt_rd_0_data_bits_10_12),
    .io_wgt_rd_0_data_bits_10_13(load_io_wgt_rd_0_data_bits_10_13),
    .io_wgt_rd_0_data_bits_10_14(load_io_wgt_rd_0_data_bits_10_14),
    .io_wgt_rd_0_data_bits_10_15(load_io_wgt_rd_0_data_bits_10_15),
    .io_wgt_rd_0_data_bits_11_0(load_io_wgt_rd_0_data_bits_11_0),
    .io_wgt_rd_0_data_bits_11_1(load_io_wgt_rd_0_data_bits_11_1),
    .io_wgt_rd_0_data_bits_11_2(load_io_wgt_rd_0_data_bits_11_2),
    .io_wgt_rd_0_data_bits_11_3(load_io_wgt_rd_0_data_bits_11_3),
    .io_wgt_rd_0_data_bits_11_4(load_io_wgt_rd_0_data_bits_11_4),
    .io_wgt_rd_0_data_bits_11_5(load_io_wgt_rd_0_data_bits_11_5),
    .io_wgt_rd_0_data_bits_11_6(load_io_wgt_rd_0_data_bits_11_6),
    .io_wgt_rd_0_data_bits_11_7(load_io_wgt_rd_0_data_bits_11_7),
    .io_wgt_rd_0_data_bits_11_8(load_io_wgt_rd_0_data_bits_11_8),
    .io_wgt_rd_0_data_bits_11_9(load_io_wgt_rd_0_data_bits_11_9),
    .io_wgt_rd_0_data_bits_11_10(load_io_wgt_rd_0_data_bits_11_10),
    .io_wgt_rd_0_data_bits_11_11(load_io_wgt_rd_0_data_bits_11_11),
    .io_wgt_rd_0_data_bits_11_12(load_io_wgt_rd_0_data_bits_11_12),
    .io_wgt_rd_0_data_bits_11_13(load_io_wgt_rd_0_data_bits_11_13),
    .io_wgt_rd_0_data_bits_11_14(load_io_wgt_rd_0_data_bits_11_14),
    .io_wgt_rd_0_data_bits_11_15(load_io_wgt_rd_0_data_bits_11_15),
    .io_wgt_rd_0_data_bits_12_0(load_io_wgt_rd_0_data_bits_12_0),
    .io_wgt_rd_0_data_bits_12_1(load_io_wgt_rd_0_data_bits_12_1),
    .io_wgt_rd_0_data_bits_12_2(load_io_wgt_rd_0_data_bits_12_2),
    .io_wgt_rd_0_data_bits_12_3(load_io_wgt_rd_0_data_bits_12_3),
    .io_wgt_rd_0_data_bits_12_4(load_io_wgt_rd_0_data_bits_12_4),
    .io_wgt_rd_0_data_bits_12_5(load_io_wgt_rd_0_data_bits_12_5),
    .io_wgt_rd_0_data_bits_12_6(load_io_wgt_rd_0_data_bits_12_6),
    .io_wgt_rd_0_data_bits_12_7(load_io_wgt_rd_0_data_bits_12_7),
    .io_wgt_rd_0_data_bits_12_8(load_io_wgt_rd_0_data_bits_12_8),
    .io_wgt_rd_0_data_bits_12_9(load_io_wgt_rd_0_data_bits_12_9),
    .io_wgt_rd_0_data_bits_12_10(load_io_wgt_rd_0_data_bits_12_10),
    .io_wgt_rd_0_data_bits_12_11(load_io_wgt_rd_0_data_bits_12_11),
    .io_wgt_rd_0_data_bits_12_12(load_io_wgt_rd_0_data_bits_12_12),
    .io_wgt_rd_0_data_bits_12_13(load_io_wgt_rd_0_data_bits_12_13),
    .io_wgt_rd_0_data_bits_12_14(load_io_wgt_rd_0_data_bits_12_14),
    .io_wgt_rd_0_data_bits_12_15(load_io_wgt_rd_0_data_bits_12_15),
    .io_wgt_rd_0_data_bits_13_0(load_io_wgt_rd_0_data_bits_13_0),
    .io_wgt_rd_0_data_bits_13_1(load_io_wgt_rd_0_data_bits_13_1),
    .io_wgt_rd_0_data_bits_13_2(load_io_wgt_rd_0_data_bits_13_2),
    .io_wgt_rd_0_data_bits_13_3(load_io_wgt_rd_0_data_bits_13_3),
    .io_wgt_rd_0_data_bits_13_4(load_io_wgt_rd_0_data_bits_13_4),
    .io_wgt_rd_0_data_bits_13_5(load_io_wgt_rd_0_data_bits_13_5),
    .io_wgt_rd_0_data_bits_13_6(load_io_wgt_rd_0_data_bits_13_6),
    .io_wgt_rd_0_data_bits_13_7(load_io_wgt_rd_0_data_bits_13_7),
    .io_wgt_rd_0_data_bits_13_8(load_io_wgt_rd_0_data_bits_13_8),
    .io_wgt_rd_0_data_bits_13_9(load_io_wgt_rd_0_data_bits_13_9),
    .io_wgt_rd_0_data_bits_13_10(load_io_wgt_rd_0_data_bits_13_10),
    .io_wgt_rd_0_data_bits_13_11(load_io_wgt_rd_0_data_bits_13_11),
    .io_wgt_rd_0_data_bits_13_12(load_io_wgt_rd_0_data_bits_13_12),
    .io_wgt_rd_0_data_bits_13_13(load_io_wgt_rd_0_data_bits_13_13),
    .io_wgt_rd_0_data_bits_13_14(load_io_wgt_rd_0_data_bits_13_14),
    .io_wgt_rd_0_data_bits_13_15(load_io_wgt_rd_0_data_bits_13_15),
    .io_wgt_rd_0_data_bits_14_0(load_io_wgt_rd_0_data_bits_14_0),
    .io_wgt_rd_0_data_bits_14_1(load_io_wgt_rd_0_data_bits_14_1),
    .io_wgt_rd_0_data_bits_14_2(load_io_wgt_rd_0_data_bits_14_2),
    .io_wgt_rd_0_data_bits_14_3(load_io_wgt_rd_0_data_bits_14_3),
    .io_wgt_rd_0_data_bits_14_4(load_io_wgt_rd_0_data_bits_14_4),
    .io_wgt_rd_0_data_bits_14_5(load_io_wgt_rd_0_data_bits_14_5),
    .io_wgt_rd_0_data_bits_14_6(load_io_wgt_rd_0_data_bits_14_6),
    .io_wgt_rd_0_data_bits_14_7(load_io_wgt_rd_0_data_bits_14_7),
    .io_wgt_rd_0_data_bits_14_8(load_io_wgt_rd_0_data_bits_14_8),
    .io_wgt_rd_0_data_bits_14_9(load_io_wgt_rd_0_data_bits_14_9),
    .io_wgt_rd_0_data_bits_14_10(load_io_wgt_rd_0_data_bits_14_10),
    .io_wgt_rd_0_data_bits_14_11(load_io_wgt_rd_0_data_bits_14_11),
    .io_wgt_rd_0_data_bits_14_12(load_io_wgt_rd_0_data_bits_14_12),
    .io_wgt_rd_0_data_bits_14_13(load_io_wgt_rd_0_data_bits_14_13),
    .io_wgt_rd_0_data_bits_14_14(load_io_wgt_rd_0_data_bits_14_14),
    .io_wgt_rd_0_data_bits_14_15(load_io_wgt_rd_0_data_bits_14_15),
    .io_wgt_rd_0_data_bits_15_0(load_io_wgt_rd_0_data_bits_15_0),
    .io_wgt_rd_0_data_bits_15_1(load_io_wgt_rd_0_data_bits_15_1),
    .io_wgt_rd_0_data_bits_15_2(load_io_wgt_rd_0_data_bits_15_2),
    .io_wgt_rd_0_data_bits_15_3(load_io_wgt_rd_0_data_bits_15_3),
    .io_wgt_rd_0_data_bits_15_4(load_io_wgt_rd_0_data_bits_15_4),
    .io_wgt_rd_0_data_bits_15_5(load_io_wgt_rd_0_data_bits_15_5),
    .io_wgt_rd_0_data_bits_15_6(load_io_wgt_rd_0_data_bits_15_6),
    .io_wgt_rd_0_data_bits_15_7(load_io_wgt_rd_0_data_bits_15_7),
    .io_wgt_rd_0_data_bits_15_8(load_io_wgt_rd_0_data_bits_15_8),
    .io_wgt_rd_0_data_bits_15_9(load_io_wgt_rd_0_data_bits_15_9),
    .io_wgt_rd_0_data_bits_15_10(load_io_wgt_rd_0_data_bits_15_10),
    .io_wgt_rd_0_data_bits_15_11(load_io_wgt_rd_0_data_bits_15_11),
    .io_wgt_rd_0_data_bits_15_12(load_io_wgt_rd_0_data_bits_15_12),
    .io_wgt_rd_0_data_bits_15_13(load_io_wgt_rd_0_data_bits_15_13),
    .io_wgt_rd_0_data_bits_15_14(load_io_wgt_rd_0_data_bits_15_14),
    .io_wgt_rd_0_data_bits_15_15(load_io_wgt_rd_0_data_bits_15_15),
    .io_wgt_rd_0_data_bits_16_0(load_io_wgt_rd_0_data_bits_16_0),
    .io_wgt_rd_0_data_bits_16_1(load_io_wgt_rd_0_data_bits_16_1),
    .io_wgt_rd_0_data_bits_16_2(load_io_wgt_rd_0_data_bits_16_2),
    .io_wgt_rd_0_data_bits_16_3(load_io_wgt_rd_0_data_bits_16_3),
    .io_wgt_rd_0_data_bits_16_4(load_io_wgt_rd_0_data_bits_16_4),
    .io_wgt_rd_0_data_bits_16_5(load_io_wgt_rd_0_data_bits_16_5),
    .io_wgt_rd_0_data_bits_16_6(load_io_wgt_rd_0_data_bits_16_6),
    .io_wgt_rd_0_data_bits_16_7(load_io_wgt_rd_0_data_bits_16_7),
    .io_wgt_rd_0_data_bits_16_8(load_io_wgt_rd_0_data_bits_16_8),
    .io_wgt_rd_0_data_bits_16_9(load_io_wgt_rd_0_data_bits_16_9),
    .io_wgt_rd_0_data_bits_16_10(load_io_wgt_rd_0_data_bits_16_10),
    .io_wgt_rd_0_data_bits_16_11(load_io_wgt_rd_0_data_bits_16_11),
    .io_wgt_rd_0_data_bits_16_12(load_io_wgt_rd_0_data_bits_16_12),
    .io_wgt_rd_0_data_bits_16_13(load_io_wgt_rd_0_data_bits_16_13),
    .io_wgt_rd_0_data_bits_16_14(load_io_wgt_rd_0_data_bits_16_14),
    .io_wgt_rd_0_data_bits_16_15(load_io_wgt_rd_0_data_bits_16_15),
    .io_wgt_rd_0_data_bits_17_0(load_io_wgt_rd_0_data_bits_17_0),
    .io_wgt_rd_0_data_bits_17_1(load_io_wgt_rd_0_data_bits_17_1),
    .io_wgt_rd_0_data_bits_17_2(load_io_wgt_rd_0_data_bits_17_2),
    .io_wgt_rd_0_data_bits_17_3(load_io_wgt_rd_0_data_bits_17_3),
    .io_wgt_rd_0_data_bits_17_4(load_io_wgt_rd_0_data_bits_17_4),
    .io_wgt_rd_0_data_bits_17_5(load_io_wgt_rd_0_data_bits_17_5),
    .io_wgt_rd_0_data_bits_17_6(load_io_wgt_rd_0_data_bits_17_6),
    .io_wgt_rd_0_data_bits_17_7(load_io_wgt_rd_0_data_bits_17_7),
    .io_wgt_rd_0_data_bits_17_8(load_io_wgt_rd_0_data_bits_17_8),
    .io_wgt_rd_0_data_bits_17_9(load_io_wgt_rd_0_data_bits_17_9),
    .io_wgt_rd_0_data_bits_17_10(load_io_wgt_rd_0_data_bits_17_10),
    .io_wgt_rd_0_data_bits_17_11(load_io_wgt_rd_0_data_bits_17_11),
    .io_wgt_rd_0_data_bits_17_12(load_io_wgt_rd_0_data_bits_17_12),
    .io_wgt_rd_0_data_bits_17_13(load_io_wgt_rd_0_data_bits_17_13),
    .io_wgt_rd_0_data_bits_17_14(load_io_wgt_rd_0_data_bits_17_14),
    .io_wgt_rd_0_data_bits_17_15(load_io_wgt_rd_0_data_bits_17_15),
    .io_wgt_rd_0_data_bits_18_0(load_io_wgt_rd_0_data_bits_18_0),
    .io_wgt_rd_0_data_bits_18_1(load_io_wgt_rd_0_data_bits_18_1),
    .io_wgt_rd_0_data_bits_18_2(load_io_wgt_rd_0_data_bits_18_2),
    .io_wgt_rd_0_data_bits_18_3(load_io_wgt_rd_0_data_bits_18_3),
    .io_wgt_rd_0_data_bits_18_4(load_io_wgt_rd_0_data_bits_18_4),
    .io_wgt_rd_0_data_bits_18_5(load_io_wgt_rd_0_data_bits_18_5),
    .io_wgt_rd_0_data_bits_18_6(load_io_wgt_rd_0_data_bits_18_6),
    .io_wgt_rd_0_data_bits_18_7(load_io_wgt_rd_0_data_bits_18_7),
    .io_wgt_rd_0_data_bits_18_8(load_io_wgt_rd_0_data_bits_18_8),
    .io_wgt_rd_0_data_bits_18_9(load_io_wgt_rd_0_data_bits_18_9),
    .io_wgt_rd_0_data_bits_18_10(load_io_wgt_rd_0_data_bits_18_10),
    .io_wgt_rd_0_data_bits_18_11(load_io_wgt_rd_0_data_bits_18_11),
    .io_wgt_rd_0_data_bits_18_12(load_io_wgt_rd_0_data_bits_18_12),
    .io_wgt_rd_0_data_bits_18_13(load_io_wgt_rd_0_data_bits_18_13),
    .io_wgt_rd_0_data_bits_18_14(load_io_wgt_rd_0_data_bits_18_14),
    .io_wgt_rd_0_data_bits_18_15(load_io_wgt_rd_0_data_bits_18_15),
    .io_wgt_rd_0_data_bits_19_0(load_io_wgt_rd_0_data_bits_19_0),
    .io_wgt_rd_0_data_bits_19_1(load_io_wgt_rd_0_data_bits_19_1),
    .io_wgt_rd_0_data_bits_19_2(load_io_wgt_rd_0_data_bits_19_2),
    .io_wgt_rd_0_data_bits_19_3(load_io_wgt_rd_0_data_bits_19_3),
    .io_wgt_rd_0_data_bits_19_4(load_io_wgt_rd_0_data_bits_19_4),
    .io_wgt_rd_0_data_bits_19_5(load_io_wgt_rd_0_data_bits_19_5),
    .io_wgt_rd_0_data_bits_19_6(load_io_wgt_rd_0_data_bits_19_6),
    .io_wgt_rd_0_data_bits_19_7(load_io_wgt_rd_0_data_bits_19_7),
    .io_wgt_rd_0_data_bits_19_8(load_io_wgt_rd_0_data_bits_19_8),
    .io_wgt_rd_0_data_bits_19_9(load_io_wgt_rd_0_data_bits_19_9),
    .io_wgt_rd_0_data_bits_19_10(load_io_wgt_rd_0_data_bits_19_10),
    .io_wgt_rd_0_data_bits_19_11(load_io_wgt_rd_0_data_bits_19_11),
    .io_wgt_rd_0_data_bits_19_12(load_io_wgt_rd_0_data_bits_19_12),
    .io_wgt_rd_0_data_bits_19_13(load_io_wgt_rd_0_data_bits_19_13),
    .io_wgt_rd_0_data_bits_19_14(load_io_wgt_rd_0_data_bits_19_14),
    .io_wgt_rd_0_data_bits_19_15(load_io_wgt_rd_0_data_bits_19_15),
    .io_wgt_rd_0_data_bits_20_0(load_io_wgt_rd_0_data_bits_20_0),
    .io_wgt_rd_0_data_bits_20_1(load_io_wgt_rd_0_data_bits_20_1),
    .io_wgt_rd_0_data_bits_20_2(load_io_wgt_rd_0_data_bits_20_2),
    .io_wgt_rd_0_data_bits_20_3(load_io_wgt_rd_0_data_bits_20_3),
    .io_wgt_rd_0_data_bits_20_4(load_io_wgt_rd_0_data_bits_20_4),
    .io_wgt_rd_0_data_bits_20_5(load_io_wgt_rd_0_data_bits_20_5),
    .io_wgt_rd_0_data_bits_20_6(load_io_wgt_rd_0_data_bits_20_6),
    .io_wgt_rd_0_data_bits_20_7(load_io_wgt_rd_0_data_bits_20_7),
    .io_wgt_rd_0_data_bits_20_8(load_io_wgt_rd_0_data_bits_20_8),
    .io_wgt_rd_0_data_bits_20_9(load_io_wgt_rd_0_data_bits_20_9),
    .io_wgt_rd_0_data_bits_20_10(load_io_wgt_rd_0_data_bits_20_10),
    .io_wgt_rd_0_data_bits_20_11(load_io_wgt_rd_0_data_bits_20_11),
    .io_wgt_rd_0_data_bits_20_12(load_io_wgt_rd_0_data_bits_20_12),
    .io_wgt_rd_0_data_bits_20_13(load_io_wgt_rd_0_data_bits_20_13),
    .io_wgt_rd_0_data_bits_20_14(load_io_wgt_rd_0_data_bits_20_14),
    .io_wgt_rd_0_data_bits_20_15(load_io_wgt_rd_0_data_bits_20_15),
    .io_wgt_rd_0_data_bits_21_0(load_io_wgt_rd_0_data_bits_21_0),
    .io_wgt_rd_0_data_bits_21_1(load_io_wgt_rd_0_data_bits_21_1),
    .io_wgt_rd_0_data_bits_21_2(load_io_wgt_rd_0_data_bits_21_2),
    .io_wgt_rd_0_data_bits_21_3(load_io_wgt_rd_0_data_bits_21_3),
    .io_wgt_rd_0_data_bits_21_4(load_io_wgt_rd_0_data_bits_21_4),
    .io_wgt_rd_0_data_bits_21_5(load_io_wgt_rd_0_data_bits_21_5),
    .io_wgt_rd_0_data_bits_21_6(load_io_wgt_rd_0_data_bits_21_6),
    .io_wgt_rd_0_data_bits_21_7(load_io_wgt_rd_0_data_bits_21_7),
    .io_wgt_rd_0_data_bits_21_8(load_io_wgt_rd_0_data_bits_21_8),
    .io_wgt_rd_0_data_bits_21_9(load_io_wgt_rd_0_data_bits_21_9),
    .io_wgt_rd_0_data_bits_21_10(load_io_wgt_rd_0_data_bits_21_10),
    .io_wgt_rd_0_data_bits_21_11(load_io_wgt_rd_0_data_bits_21_11),
    .io_wgt_rd_0_data_bits_21_12(load_io_wgt_rd_0_data_bits_21_12),
    .io_wgt_rd_0_data_bits_21_13(load_io_wgt_rd_0_data_bits_21_13),
    .io_wgt_rd_0_data_bits_21_14(load_io_wgt_rd_0_data_bits_21_14),
    .io_wgt_rd_0_data_bits_21_15(load_io_wgt_rd_0_data_bits_21_15),
    .io_wgt_rd_0_data_bits_22_0(load_io_wgt_rd_0_data_bits_22_0),
    .io_wgt_rd_0_data_bits_22_1(load_io_wgt_rd_0_data_bits_22_1),
    .io_wgt_rd_0_data_bits_22_2(load_io_wgt_rd_0_data_bits_22_2),
    .io_wgt_rd_0_data_bits_22_3(load_io_wgt_rd_0_data_bits_22_3),
    .io_wgt_rd_0_data_bits_22_4(load_io_wgt_rd_0_data_bits_22_4),
    .io_wgt_rd_0_data_bits_22_5(load_io_wgt_rd_0_data_bits_22_5),
    .io_wgt_rd_0_data_bits_22_6(load_io_wgt_rd_0_data_bits_22_6),
    .io_wgt_rd_0_data_bits_22_7(load_io_wgt_rd_0_data_bits_22_7),
    .io_wgt_rd_0_data_bits_22_8(load_io_wgt_rd_0_data_bits_22_8),
    .io_wgt_rd_0_data_bits_22_9(load_io_wgt_rd_0_data_bits_22_9),
    .io_wgt_rd_0_data_bits_22_10(load_io_wgt_rd_0_data_bits_22_10),
    .io_wgt_rd_0_data_bits_22_11(load_io_wgt_rd_0_data_bits_22_11),
    .io_wgt_rd_0_data_bits_22_12(load_io_wgt_rd_0_data_bits_22_12),
    .io_wgt_rd_0_data_bits_22_13(load_io_wgt_rd_0_data_bits_22_13),
    .io_wgt_rd_0_data_bits_22_14(load_io_wgt_rd_0_data_bits_22_14),
    .io_wgt_rd_0_data_bits_22_15(load_io_wgt_rd_0_data_bits_22_15),
    .io_wgt_rd_0_data_bits_23_0(load_io_wgt_rd_0_data_bits_23_0),
    .io_wgt_rd_0_data_bits_23_1(load_io_wgt_rd_0_data_bits_23_1),
    .io_wgt_rd_0_data_bits_23_2(load_io_wgt_rd_0_data_bits_23_2),
    .io_wgt_rd_0_data_bits_23_3(load_io_wgt_rd_0_data_bits_23_3),
    .io_wgt_rd_0_data_bits_23_4(load_io_wgt_rd_0_data_bits_23_4),
    .io_wgt_rd_0_data_bits_23_5(load_io_wgt_rd_0_data_bits_23_5),
    .io_wgt_rd_0_data_bits_23_6(load_io_wgt_rd_0_data_bits_23_6),
    .io_wgt_rd_0_data_bits_23_7(load_io_wgt_rd_0_data_bits_23_7),
    .io_wgt_rd_0_data_bits_23_8(load_io_wgt_rd_0_data_bits_23_8),
    .io_wgt_rd_0_data_bits_23_9(load_io_wgt_rd_0_data_bits_23_9),
    .io_wgt_rd_0_data_bits_23_10(load_io_wgt_rd_0_data_bits_23_10),
    .io_wgt_rd_0_data_bits_23_11(load_io_wgt_rd_0_data_bits_23_11),
    .io_wgt_rd_0_data_bits_23_12(load_io_wgt_rd_0_data_bits_23_12),
    .io_wgt_rd_0_data_bits_23_13(load_io_wgt_rd_0_data_bits_23_13),
    .io_wgt_rd_0_data_bits_23_14(load_io_wgt_rd_0_data_bits_23_14),
    .io_wgt_rd_0_data_bits_23_15(load_io_wgt_rd_0_data_bits_23_15),
    .io_wgt_rd_0_data_bits_24_0(load_io_wgt_rd_0_data_bits_24_0),
    .io_wgt_rd_0_data_bits_24_1(load_io_wgt_rd_0_data_bits_24_1),
    .io_wgt_rd_0_data_bits_24_2(load_io_wgt_rd_0_data_bits_24_2),
    .io_wgt_rd_0_data_bits_24_3(load_io_wgt_rd_0_data_bits_24_3),
    .io_wgt_rd_0_data_bits_24_4(load_io_wgt_rd_0_data_bits_24_4),
    .io_wgt_rd_0_data_bits_24_5(load_io_wgt_rd_0_data_bits_24_5),
    .io_wgt_rd_0_data_bits_24_6(load_io_wgt_rd_0_data_bits_24_6),
    .io_wgt_rd_0_data_bits_24_7(load_io_wgt_rd_0_data_bits_24_7),
    .io_wgt_rd_0_data_bits_24_8(load_io_wgt_rd_0_data_bits_24_8),
    .io_wgt_rd_0_data_bits_24_9(load_io_wgt_rd_0_data_bits_24_9),
    .io_wgt_rd_0_data_bits_24_10(load_io_wgt_rd_0_data_bits_24_10),
    .io_wgt_rd_0_data_bits_24_11(load_io_wgt_rd_0_data_bits_24_11),
    .io_wgt_rd_0_data_bits_24_12(load_io_wgt_rd_0_data_bits_24_12),
    .io_wgt_rd_0_data_bits_24_13(load_io_wgt_rd_0_data_bits_24_13),
    .io_wgt_rd_0_data_bits_24_14(load_io_wgt_rd_0_data_bits_24_14),
    .io_wgt_rd_0_data_bits_24_15(load_io_wgt_rd_0_data_bits_24_15),
    .io_wgt_rd_0_data_bits_25_0(load_io_wgt_rd_0_data_bits_25_0),
    .io_wgt_rd_0_data_bits_25_1(load_io_wgt_rd_0_data_bits_25_1),
    .io_wgt_rd_0_data_bits_25_2(load_io_wgt_rd_0_data_bits_25_2),
    .io_wgt_rd_0_data_bits_25_3(load_io_wgt_rd_0_data_bits_25_3),
    .io_wgt_rd_0_data_bits_25_4(load_io_wgt_rd_0_data_bits_25_4),
    .io_wgt_rd_0_data_bits_25_5(load_io_wgt_rd_0_data_bits_25_5),
    .io_wgt_rd_0_data_bits_25_6(load_io_wgt_rd_0_data_bits_25_6),
    .io_wgt_rd_0_data_bits_25_7(load_io_wgt_rd_0_data_bits_25_7),
    .io_wgt_rd_0_data_bits_25_8(load_io_wgt_rd_0_data_bits_25_8),
    .io_wgt_rd_0_data_bits_25_9(load_io_wgt_rd_0_data_bits_25_9),
    .io_wgt_rd_0_data_bits_25_10(load_io_wgt_rd_0_data_bits_25_10),
    .io_wgt_rd_0_data_bits_25_11(load_io_wgt_rd_0_data_bits_25_11),
    .io_wgt_rd_0_data_bits_25_12(load_io_wgt_rd_0_data_bits_25_12),
    .io_wgt_rd_0_data_bits_25_13(load_io_wgt_rd_0_data_bits_25_13),
    .io_wgt_rd_0_data_bits_25_14(load_io_wgt_rd_0_data_bits_25_14),
    .io_wgt_rd_0_data_bits_25_15(load_io_wgt_rd_0_data_bits_25_15),
    .io_wgt_rd_0_data_bits_26_0(load_io_wgt_rd_0_data_bits_26_0),
    .io_wgt_rd_0_data_bits_26_1(load_io_wgt_rd_0_data_bits_26_1),
    .io_wgt_rd_0_data_bits_26_2(load_io_wgt_rd_0_data_bits_26_2),
    .io_wgt_rd_0_data_bits_26_3(load_io_wgt_rd_0_data_bits_26_3),
    .io_wgt_rd_0_data_bits_26_4(load_io_wgt_rd_0_data_bits_26_4),
    .io_wgt_rd_0_data_bits_26_5(load_io_wgt_rd_0_data_bits_26_5),
    .io_wgt_rd_0_data_bits_26_6(load_io_wgt_rd_0_data_bits_26_6),
    .io_wgt_rd_0_data_bits_26_7(load_io_wgt_rd_0_data_bits_26_7),
    .io_wgt_rd_0_data_bits_26_8(load_io_wgt_rd_0_data_bits_26_8),
    .io_wgt_rd_0_data_bits_26_9(load_io_wgt_rd_0_data_bits_26_9),
    .io_wgt_rd_0_data_bits_26_10(load_io_wgt_rd_0_data_bits_26_10),
    .io_wgt_rd_0_data_bits_26_11(load_io_wgt_rd_0_data_bits_26_11),
    .io_wgt_rd_0_data_bits_26_12(load_io_wgt_rd_0_data_bits_26_12),
    .io_wgt_rd_0_data_bits_26_13(load_io_wgt_rd_0_data_bits_26_13),
    .io_wgt_rd_0_data_bits_26_14(load_io_wgt_rd_0_data_bits_26_14),
    .io_wgt_rd_0_data_bits_26_15(load_io_wgt_rd_0_data_bits_26_15),
    .io_wgt_rd_0_data_bits_27_0(load_io_wgt_rd_0_data_bits_27_0),
    .io_wgt_rd_0_data_bits_27_1(load_io_wgt_rd_0_data_bits_27_1),
    .io_wgt_rd_0_data_bits_27_2(load_io_wgt_rd_0_data_bits_27_2),
    .io_wgt_rd_0_data_bits_27_3(load_io_wgt_rd_0_data_bits_27_3),
    .io_wgt_rd_0_data_bits_27_4(load_io_wgt_rd_0_data_bits_27_4),
    .io_wgt_rd_0_data_bits_27_5(load_io_wgt_rd_0_data_bits_27_5),
    .io_wgt_rd_0_data_bits_27_6(load_io_wgt_rd_0_data_bits_27_6),
    .io_wgt_rd_0_data_bits_27_7(load_io_wgt_rd_0_data_bits_27_7),
    .io_wgt_rd_0_data_bits_27_8(load_io_wgt_rd_0_data_bits_27_8),
    .io_wgt_rd_0_data_bits_27_9(load_io_wgt_rd_0_data_bits_27_9),
    .io_wgt_rd_0_data_bits_27_10(load_io_wgt_rd_0_data_bits_27_10),
    .io_wgt_rd_0_data_bits_27_11(load_io_wgt_rd_0_data_bits_27_11),
    .io_wgt_rd_0_data_bits_27_12(load_io_wgt_rd_0_data_bits_27_12),
    .io_wgt_rd_0_data_bits_27_13(load_io_wgt_rd_0_data_bits_27_13),
    .io_wgt_rd_0_data_bits_27_14(load_io_wgt_rd_0_data_bits_27_14),
    .io_wgt_rd_0_data_bits_27_15(load_io_wgt_rd_0_data_bits_27_15),
    .io_wgt_rd_0_data_bits_28_0(load_io_wgt_rd_0_data_bits_28_0),
    .io_wgt_rd_0_data_bits_28_1(load_io_wgt_rd_0_data_bits_28_1),
    .io_wgt_rd_0_data_bits_28_2(load_io_wgt_rd_0_data_bits_28_2),
    .io_wgt_rd_0_data_bits_28_3(load_io_wgt_rd_0_data_bits_28_3),
    .io_wgt_rd_0_data_bits_28_4(load_io_wgt_rd_0_data_bits_28_4),
    .io_wgt_rd_0_data_bits_28_5(load_io_wgt_rd_0_data_bits_28_5),
    .io_wgt_rd_0_data_bits_28_6(load_io_wgt_rd_0_data_bits_28_6),
    .io_wgt_rd_0_data_bits_28_7(load_io_wgt_rd_0_data_bits_28_7),
    .io_wgt_rd_0_data_bits_28_8(load_io_wgt_rd_0_data_bits_28_8),
    .io_wgt_rd_0_data_bits_28_9(load_io_wgt_rd_0_data_bits_28_9),
    .io_wgt_rd_0_data_bits_28_10(load_io_wgt_rd_0_data_bits_28_10),
    .io_wgt_rd_0_data_bits_28_11(load_io_wgt_rd_0_data_bits_28_11),
    .io_wgt_rd_0_data_bits_28_12(load_io_wgt_rd_0_data_bits_28_12),
    .io_wgt_rd_0_data_bits_28_13(load_io_wgt_rd_0_data_bits_28_13),
    .io_wgt_rd_0_data_bits_28_14(load_io_wgt_rd_0_data_bits_28_14),
    .io_wgt_rd_0_data_bits_28_15(load_io_wgt_rd_0_data_bits_28_15),
    .io_wgt_rd_0_data_bits_29_0(load_io_wgt_rd_0_data_bits_29_0),
    .io_wgt_rd_0_data_bits_29_1(load_io_wgt_rd_0_data_bits_29_1),
    .io_wgt_rd_0_data_bits_29_2(load_io_wgt_rd_0_data_bits_29_2),
    .io_wgt_rd_0_data_bits_29_3(load_io_wgt_rd_0_data_bits_29_3),
    .io_wgt_rd_0_data_bits_29_4(load_io_wgt_rd_0_data_bits_29_4),
    .io_wgt_rd_0_data_bits_29_5(load_io_wgt_rd_0_data_bits_29_5),
    .io_wgt_rd_0_data_bits_29_6(load_io_wgt_rd_0_data_bits_29_6),
    .io_wgt_rd_0_data_bits_29_7(load_io_wgt_rd_0_data_bits_29_7),
    .io_wgt_rd_0_data_bits_29_8(load_io_wgt_rd_0_data_bits_29_8),
    .io_wgt_rd_0_data_bits_29_9(load_io_wgt_rd_0_data_bits_29_9),
    .io_wgt_rd_0_data_bits_29_10(load_io_wgt_rd_0_data_bits_29_10),
    .io_wgt_rd_0_data_bits_29_11(load_io_wgt_rd_0_data_bits_29_11),
    .io_wgt_rd_0_data_bits_29_12(load_io_wgt_rd_0_data_bits_29_12),
    .io_wgt_rd_0_data_bits_29_13(load_io_wgt_rd_0_data_bits_29_13),
    .io_wgt_rd_0_data_bits_29_14(load_io_wgt_rd_0_data_bits_29_14),
    .io_wgt_rd_0_data_bits_29_15(load_io_wgt_rd_0_data_bits_29_15),
    .io_wgt_rd_0_data_bits_30_0(load_io_wgt_rd_0_data_bits_30_0),
    .io_wgt_rd_0_data_bits_30_1(load_io_wgt_rd_0_data_bits_30_1),
    .io_wgt_rd_0_data_bits_30_2(load_io_wgt_rd_0_data_bits_30_2),
    .io_wgt_rd_0_data_bits_30_3(load_io_wgt_rd_0_data_bits_30_3),
    .io_wgt_rd_0_data_bits_30_4(load_io_wgt_rd_0_data_bits_30_4),
    .io_wgt_rd_0_data_bits_30_5(load_io_wgt_rd_0_data_bits_30_5),
    .io_wgt_rd_0_data_bits_30_6(load_io_wgt_rd_0_data_bits_30_6),
    .io_wgt_rd_0_data_bits_30_7(load_io_wgt_rd_0_data_bits_30_7),
    .io_wgt_rd_0_data_bits_30_8(load_io_wgt_rd_0_data_bits_30_8),
    .io_wgt_rd_0_data_bits_30_9(load_io_wgt_rd_0_data_bits_30_9),
    .io_wgt_rd_0_data_bits_30_10(load_io_wgt_rd_0_data_bits_30_10),
    .io_wgt_rd_0_data_bits_30_11(load_io_wgt_rd_0_data_bits_30_11),
    .io_wgt_rd_0_data_bits_30_12(load_io_wgt_rd_0_data_bits_30_12),
    .io_wgt_rd_0_data_bits_30_13(load_io_wgt_rd_0_data_bits_30_13),
    .io_wgt_rd_0_data_bits_30_14(load_io_wgt_rd_0_data_bits_30_14),
    .io_wgt_rd_0_data_bits_30_15(load_io_wgt_rd_0_data_bits_30_15),
    .io_wgt_rd_0_data_bits_31_0(load_io_wgt_rd_0_data_bits_31_0),
    .io_wgt_rd_0_data_bits_31_1(load_io_wgt_rd_0_data_bits_31_1),
    .io_wgt_rd_0_data_bits_31_2(load_io_wgt_rd_0_data_bits_31_2),
    .io_wgt_rd_0_data_bits_31_3(load_io_wgt_rd_0_data_bits_31_3),
    .io_wgt_rd_0_data_bits_31_4(load_io_wgt_rd_0_data_bits_31_4),
    .io_wgt_rd_0_data_bits_31_5(load_io_wgt_rd_0_data_bits_31_5),
    .io_wgt_rd_0_data_bits_31_6(load_io_wgt_rd_0_data_bits_31_6),
    .io_wgt_rd_0_data_bits_31_7(load_io_wgt_rd_0_data_bits_31_7),
    .io_wgt_rd_0_data_bits_31_8(load_io_wgt_rd_0_data_bits_31_8),
    .io_wgt_rd_0_data_bits_31_9(load_io_wgt_rd_0_data_bits_31_9),
    .io_wgt_rd_0_data_bits_31_10(load_io_wgt_rd_0_data_bits_31_10),
    .io_wgt_rd_0_data_bits_31_11(load_io_wgt_rd_0_data_bits_31_11),
    .io_wgt_rd_0_data_bits_31_12(load_io_wgt_rd_0_data_bits_31_12),
    .io_wgt_rd_0_data_bits_31_13(load_io_wgt_rd_0_data_bits_31_13),
    .io_wgt_rd_0_data_bits_31_14(load_io_wgt_rd_0_data_bits_31_14),
    .io_wgt_rd_0_data_bits_31_15(load_io_wgt_rd_0_data_bits_31_15)
  );
  Compute compute ( // @[Core.scala 69:23]
    .clock(compute_clock),
    .reset(compute_reset),
    .io_i_post_0(compute_io_i_post_0),
    .io_i_post_1(compute_io_i_post_1),
    .io_o_post_0(compute_io_o_post_0),
    .io_o_post_1(compute_io_o_post_1),
    .io_inst_ready(compute_io_inst_ready),
    .io_inst_valid(compute_io_inst_valid),
    .io_inst_bits(compute_io_inst_bits),
    .io_uop_baddr(compute_io_uop_baddr),
    .io_acc_baddr(compute_io_acc_baddr),
    .io_vme_rd_0_cmd_ready(compute_io_vme_rd_0_cmd_ready),
    .io_vme_rd_0_cmd_valid(compute_io_vme_rd_0_cmd_valid),
    .io_vme_rd_0_cmd_bits_addr(compute_io_vme_rd_0_cmd_bits_addr),
    .io_vme_rd_0_cmd_bits_len(compute_io_vme_rd_0_cmd_bits_len),
    .io_vme_rd_0_cmd_bits_tag(compute_io_vme_rd_0_cmd_bits_tag),
    .io_vme_rd_0_data_valid(compute_io_vme_rd_0_data_valid),
    .io_vme_rd_0_data_bits_data(compute_io_vme_rd_0_data_bits_data),
    .io_vme_rd_0_data_bits_tag(compute_io_vme_rd_0_data_bits_tag),
    .io_vme_rd_0_data_bits_last(compute_io_vme_rd_0_data_bits_last),
    .io_vme_rd_1_cmd_ready(compute_io_vme_rd_1_cmd_ready),
    .io_vme_rd_1_cmd_valid(compute_io_vme_rd_1_cmd_valid),
    .io_vme_rd_1_cmd_bits_addr(compute_io_vme_rd_1_cmd_bits_addr),
    .io_vme_rd_1_cmd_bits_len(compute_io_vme_rd_1_cmd_bits_len),
    .io_vme_rd_1_cmd_bits_tag(compute_io_vme_rd_1_cmd_bits_tag),
    .io_vme_rd_1_data_valid(compute_io_vme_rd_1_data_valid),
    .io_vme_rd_1_data_bits_data(compute_io_vme_rd_1_data_bits_data),
    .io_vme_rd_1_data_bits_tag(compute_io_vme_rd_1_data_bits_tag),
    .io_inp_rd_0_idx_valid(compute_io_inp_rd_0_idx_valid),
    .io_inp_rd_0_idx_bits(compute_io_inp_rd_0_idx_bits),
    .io_inp_rd_0_data_valid(compute_io_inp_rd_0_data_valid),
    .io_inp_rd_0_data_bits_0_0(compute_io_inp_rd_0_data_bits_0_0),
    .io_inp_rd_0_data_bits_0_1(compute_io_inp_rd_0_data_bits_0_1),
    .io_inp_rd_0_data_bits_0_2(compute_io_inp_rd_0_data_bits_0_2),
    .io_inp_rd_0_data_bits_0_3(compute_io_inp_rd_0_data_bits_0_3),
    .io_inp_rd_0_data_bits_0_4(compute_io_inp_rd_0_data_bits_0_4),
    .io_inp_rd_0_data_bits_0_5(compute_io_inp_rd_0_data_bits_0_5),
    .io_inp_rd_0_data_bits_0_6(compute_io_inp_rd_0_data_bits_0_6),
    .io_inp_rd_0_data_bits_0_7(compute_io_inp_rd_0_data_bits_0_7),
    .io_inp_rd_0_data_bits_0_8(compute_io_inp_rd_0_data_bits_0_8),
    .io_inp_rd_0_data_bits_0_9(compute_io_inp_rd_0_data_bits_0_9),
    .io_inp_rd_0_data_bits_0_10(compute_io_inp_rd_0_data_bits_0_10),
    .io_inp_rd_0_data_bits_0_11(compute_io_inp_rd_0_data_bits_0_11),
    .io_inp_rd_0_data_bits_0_12(compute_io_inp_rd_0_data_bits_0_12),
    .io_inp_rd_0_data_bits_0_13(compute_io_inp_rd_0_data_bits_0_13),
    .io_inp_rd_0_data_bits_0_14(compute_io_inp_rd_0_data_bits_0_14),
    .io_inp_rd_0_data_bits_0_15(compute_io_inp_rd_0_data_bits_0_15),
    .io_wgt_rd_0_idx_valid(compute_io_wgt_rd_0_idx_valid),
    .io_wgt_rd_0_idx_bits(compute_io_wgt_rd_0_idx_bits),
    .io_wgt_rd_0_data_valid(compute_io_wgt_rd_0_data_valid),
    .io_wgt_rd_0_data_bits_0_0(compute_io_wgt_rd_0_data_bits_0_0),
    .io_wgt_rd_0_data_bits_0_1(compute_io_wgt_rd_0_data_bits_0_1),
    .io_wgt_rd_0_data_bits_0_2(compute_io_wgt_rd_0_data_bits_0_2),
    .io_wgt_rd_0_data_bits_0_3(compute_io_wgt_rd_0_data_bits_0_3),
    .io_wgt_rd_0_data_bits_0_4(compute_io_wgt_rd_0_data_bits_0_4),
    .io_wgt_rd_0_data_bits_0_5(compute_io_wgt_rd_0_data_bits_0_5),
    .io_wgt_rd_0_data_bits_0_6(compute_io_wgt_rd_0_data_bits_0_6),
    .io_wgt_rd_0_data_bits_0_7(compute_io_wgt_rd_0_data_bits_0_7),
    .io_wgt_rd_0_data_bits_0_8(compute_io_wgt_rd_0_data_bits_0_8),
    .io_wgt_rd_0_data_bits_0_9(compute_io_wgt_rd_0_data_bits_0_9),
    .io_wgt_rd_0_data_bits_0_10(compute_io_wgt_rd_0_data_bits_0_10),
    .io_wgt_rd_0_data_bits_0_11(compute_io_wgt_rd_0_data_bits_0_11),
    .io_wgt_rd_0_data_bits_0_12(compute_io_wgt_rd_0_data_bits_0_12),
    .io_wgt_rd_0_data_bits_0_13(compute_io_wgt_rd_0_data_bits_0_13),
    .io_wgt_rd_0_data_bits_0_14(compute_io_wgt_rd_0_data_bits_0_14),
    .io_wgt_rd_0_data_bits_0_15(compute_io_wgt_rd_0_data_bits_0_15),
    .io_wgt_rd_0_data_bits_1_0(compute_io_wgt_rd_0_data_bits_1_0),
    .io_wgt_rd_0_data_bits_1_1(compute_io_wgt_rd_0_data_bits_1_1),
    .io_wgt_rd_0_data_bits_1_2(compute_io_wgt_rd_0_data_bits_1_2),
    .io_wgt_rd_0_data_bits_1_3(compute_io_wgt_rd_0_data_bits_1_3),
    .io_wgt_rd_0_data_bits_1_4(compute_io_wgt_rd_0_data_bits_1_4),
    .io_wgt_rd_0_data_bits_1_5(compute_io_wgt_rd_0_data_bits_1_5),
    .io_wgt_rd_0_data_bits_1_6(compute_io_wgt_rd_0_data_bits_1_6),
    .io_wgt_rd_0_data_bits_1_7(compute_io_wgt_rd_0_data_bits_1_7),
    .io_wgt_rd_0_data_bits_1_8(compute_io_wgt_rd_0_data_bits_1_8),
    .io_wgt_rd_0_data_bits_1_9(compute_io_wgt_rd_0_data_bits_1_9),
    .io_wgt_rd_0_data_bits_1_10(compute_io_wgt_rd_0_data_bits_1_10),
    .io_wgt_rd_0_data_bits_1_11(compute_io_wgt_rd_0_data_bits_1_11),
    .io_wgt_rd_0_data_bits_1_12(compute_io_wgt_rd_0_data_bits_1_12),
    .io_wgt_rd_0_data_bits_1_13(compute_io_wgt_rd_0_data_bits_1_13),
    .io_wgt_rd_0_data_bits_1_14(compute_io_wgt_rd_0_data_bits_1_14),
    .io_wgt_rd_0_data_bits_1_15(compute_io_wgt_rd_0_data_bits_1_15),
    .io_wgt_rd_0_data_bits_2_0(compute_io_wgt_rd_0_data_bits_2_0),
    .io_wgt_rd_0_data_bits_2_1(compute_io_wgt_rd_0_data_bits_2_1),
    .io_wgt_rd_0_data_bits_2_2(compute_io_wgt_rd_0_data_bits_2_2),
    .io_wgt_rd_0_data_bits_2_3(compute_io_wgt_rd_0_data_bits_2_3),
    .io_wgt_rd_0_data_bits_2_4(compute_io_wgt_rd_0_data_bits_2_4),
    .io_wgt_rd_0_data_bits_2_5(compute_io_wgt_rd_0_data_bits_2_5),
    .io_wgt_rd_0_data_bits_2_6(compute_io_wgt_rd_0_data_bits_2_6),
    .io_wgt_rd_0_data_bits_2_7(compute_io_wgt_rd_0_data_bits_2_7),
    .io_wgt_rd_0_data_bits_2_8(compute_io_wgt_rd_0_data_bits_2_8),
    .io_wgt_rd_0_data_bits_2_9(compute_io_wgt_rd_0_data_bits_2_9),
    .io_wgt_rd_0_data_bits_2_10(compute_io_wgt_rd_0_data_bits_2_10),
    .io_wgt_rd_0_data_bits_2_11(compute_io_wgt_rd_0_data_bits_2_11),
    .io_wgt_rd_0_data_bits_2_12(compute_io_wgt_rd_0_data_bits_2_12),
    .io_wgt_rd_0_data_bits_2_13(compute_io_wgt_rd_0_data_bits_2_13),
    .io_wgt_rd_0_data_bits_2_14(compute_io_wgt_rd_0_data_bits_2_14),
    .io_wgt_rd_0_data_bits_2_15(compute_io_wgt_rd_0_data_bits_2_15),
    .io_wgt_rd_0_data_bits_3_0(compute_io_wgt_rd_0_data_bits_3_0),
    .io_wgt_rd_0_data_bits_3_1(compute_io_wgt_rd_0_data_bits_3_1),
    .io_wgt_rd_0_data_bits_3_2(compute_io_wgt_rd_0_data_bits_3_2),
    .io_wgt_rd_0_data_bits_3_3(compute_io_wgt_rd_0_data_bits_3_3),
    .io_wgt_rd_0_data_bits_3_4(compute_io_wgt_rd_0_data_bits_3_4),
    .io_wgt_rd_0_data_bits_3_5(compute_io_wgt_rd_0_data_bits_3_5),
    .io_wgt_rd_0_data_bits_3_6(compute_io_wgt_rd_0_data_bits_3_6),
    .io_wgt_rd_0_data_bits_3_7(compute_io_wgt_rd_0_data_bits_3_7),
    .io_wgt_rd_0_data_bits_3_8(compute_io_wgt_rd_0_data_bits_3_8),
    .io_wgt_rd_0_data_bits_3_9(compute_io_wgt_rd_0_data_bits_3_9),
    .io_wgt_rd_0_data_bits_3_10(compute_io_wgt_rd_0_data_bits_3_10),
    .io_wgt_rd_0_data_bits_3_11(compute_io_wgt_rd_0_data_bits_3_11),
    .io_wgt_rd_0_data_bits_3_12(compute_io_wgt_rd_0_data_bits_3_12),
    .io_wgt_rd_0_data_bits_3_13(compute_io_wgt_rd_0_data_bits_3_13),
    .io_wgt_rd_0_data_bits_3_14(compute_io_wgt_rd_0_data_bits_3_14),
    .io_wgt_rd_0_data_bits_3_15(compute_io_wgt_rd_0_data_bits_3_15),
    .io_wgt_rd_0_data_bits_4_0(compute_io_wgt_rd_0_data_bits_4_0),
    .io_wgt_rd_0_data_bits_4_1(compute_io_wgt_rd_0_data_bits_4_1),
    .io_wgt_rd_0_data_bits_4_2(compute_io_wgt_rd_0_data_bits_4_2),
    .io_wgt_rd_0_data_bits_4_3(compute_io_wgt_rd_0_data_bits_4_3),
    .io_wgt_rd_0_data_bits_4_4(compute_io_wgt_rd_0_data_bits_4_4),
    .io_wgt_rd_0_data_bits_4_5(compute_io_wgt_rd_0_data_bits_4_5),
    .io_wgt_rd_0_data_bits_4_6(compute_io_wgt_rd_0_data_bits_4_6),
    .io_wgt_rd_0_data_bits_4_7(compute_io_wgt_rd_0_data_bits_4_7),
    .io_wgt_rd_0_data_bits_4_8(compute_io_wgt_rd_0_data_bits_4_8),
    .io_wgt_rd_0_data_bits_4_9(compute_io_wgt_rd_0_data_bits_4_9),
    .io_wgt_rd_0_data_bits_4_10(compute_io_wgt_rd_0_data_bits_4_10),
    .io_wgt_rd_0_data_bits_4_11(compute_io_wgt_rd_0_data_bits_4_11),
    .io_wgt_rd_0_data_bits_4_12(compute_io_wgt_rd_0_data_bits_4_12),
    .io_wgt_rd_0_data_bits_4_13(compute_io_wgt_rd_0_data_bits_4_13),
    .io_wgt_rd_0_data_bits_4_14(compute_io_wgt_rd_0_data_bits_4_14),
    .io_wgt_rd_0_data_bits_4_15(compute_io_wgt_rd_0_data_bits_4_15),
    .io_wgt_rd_0_data_bits_5_0(compute_io_wgt_rd_0_data_bits_5_0),
    .io_wgt_rd_0_data_bits_5_1(compute_io_wgt_rd_0_data_bits_5_1),
    .io_wgt_rd_0_data_bits_5_2(compute_io_wgt_rd_0_data_bits_5_2),
    .io_wgt_rd_0_data_bits_5_3(compute_io_wgt_rd_0_data_bits_5_3),
    .io_wgt_rd_0_data_bits_5_4(compute_io_wgt_rd_0_data_bits_5_4),
    .io_wgt_rd_0_data_bits_5_5(compute_io_wgt_rd_0_data_bits_5_5),
    .io_wgt_rd_0_data_bits_5_6(compute_io_wgt_rd_0_data_bits_5_6),
    .io_wgt_rd_0_data_bits_5_7(compute_io_wgt_rd_0_data_bits_5_7),
    .io_wgt_rd_0_data_bits_5_8(compute_io_wgt_rd_0_data_bits_5_8),
    .io_wgt_rd_0_data_bits_5_9(compute_io_wgt_rd_0_data_bits_5_9),
    .io_wgt_rd_0_data_bits_5_10(compute_io_wgt_rd_0_data_bits_5_10),
    .io_wgt_rd_0_data_bits_5_11(compute_io_wgt_rd_0_data_bits_5_11),
    .io_wgt_rd_0_data_bits_5_12(compute_io_wgt_rd_0_data_bits_5_12),
    .io_wgt_rd_0_data_bits_5_13(compute_io_wgt_rd_0_data_bits_5_13),
    .io_wgt_rd_0_data_bits_5_14(compute_io_wgt_rd_0_data_bits_5_14),
    .io_wgt_rd_0_data_bits_5_15(compute_io_wgt_rd_0_data_bits_5_15),
    .io_wgt_rd_0_data_bits_6_0(compute_io_wgt_rd_0_data_bits_6_0),
    .io_wgt_rd_0_data_bits_6_1(compute_io_wgt_rd_0_data_bits_6_1),
    .io_wgt_rd_0_data_bits_6_2(compute_io_wgt_rd_0_data_bits_6_2),
    .io_wgt_rd_0_data_bits_6_3(compute_io_wgt_rd_0_data_bits_6_3),
    .io_wgt_rd_0_data_bits_6_4(compute_io_wgt_rd_0_data_bits_6_4),
    .io_wgt_rd_0_data_bits_6_5(compute_io_wgt_rd_0_data_bits_6_5),
    .io_wgt_rd_0_data_bits_6_6(compute_io_wgt_rd_0_data_bits_6_6),
    .io_wgt_rd_0_data_bits_6_7(compute_io_wgt_rd_0_data_bits_6_7),
    .io_wgt_rd_0_data_bits_6_8(compute_io_wgt_rd_0_data_bits_6_8),
    .io_wgt_rd_0_data_bits_6_9(compute_io_wgt_rd_0_data_bits_6_9),
    .io_wgt_rd_0_data_bits_6_10(compute_io_wgt_rd_0_data_bits_6_10),
    .io_wgt_rd_0_data_bits_6_11(compute_io_wgt_rd_0_data_bits_6_11),
    .io_wgt_rd_0_data_bits_6_12(compute_io_wgt_rd_0_data_bits_6_12),
    .io_wgt_rd_0_data_bits_6_13(compute_io_wgt_rd_0_data_bits_6_13),
    .io_wgt_rd_0_data_bits_6_14(compute_io_wgt_rd_0_data_bits_6_14),
    .io_wgt_rd_0_data_bits_6_15(compute_io_wgt_rd_0_data_bits_6_15),
    .io_wgt_rd_0_data_bits_7_0(compute_io_wgt_rd_0_data_bits_7_0),
    .io_wgt_rd_0_data_bits_7_1(compute_io_wgt_rd_0_data_bits_7_1),
    .io_wgt_rd_0_data_bits_7_2(compute_io_wgt_rd_0_data_bits_7_2),
    .io_wgt_rd_0_data_bits_7_3(compute_io_wgt_rd_0_data_bits_7_3),
    .io_wgt_rd_0_data_bits_7_4(compute_io_wgt_rd_0_data_bits_7_4),
    .io_wgt_rd_0_data_bits_7_5(compute_io_wgt_rd_0_data_bits_7_5),
    .io_wgt_rd_0_data_bits_7_6(compute_io_wgt_rd_0_data_bits_7_6),
    .io_wgt_rd_0_data_bits_7_7(compute_io_wgt_rd_0_data_bits_7_7),
    .io_wgt_rd_0_data_bits_7_8(compute_io_wgt_rd_0_data_bits_7_8),
    .io_wgt_rd_0_data_bits_7_9(compute_io_wgt_rd_0_data_bits_7_9),
    .io_wgt_rd_0_data_bits_7_10(compute_io_wgt_rd_0_data_bits_7_10),
    .io_wgt_rd_0_data_bits_7_11(compute_io_wgt_rd_0_data_bits_7_11),
    .io_wgt_rd_0_data_bits_7_12(compute_io_wgt_rd_0_data_bits_7_12),
    .io_wgt_rd_0_data_bits_7_13(compute_io_wgt_rd_0_data_bits_7_13),
    .io_wgt_rd_0_data_bits_7_14(compute_io_wgt_rd_0_data_bits_7_14),
    .io_wgt_rd_0_data_bits_7_15(compute_io_wgt_rd_0_data_bits_7_15),
    .io_wgt_rd_0_data_bits_8_0(compute_io_wgt_rd_0_data_bits_8_0),
    .io_wgt_rd_0_data_bits_8_1(compute_io_wgt_rd_0_data_bits_8_1),
    .io_wgt_rd_0_data_bits_8_2(compute_io_wgt_rd_0_data_bits_8_2),
    .io_wgt_rd_0_data_bits_8_3(compute_io_wgt_rd_0_data_bits_8_3),
    .io_wgt_rd_0_data_bits_8_4(compute_io_wgt_rd_0_data_bits_8_4),
    .io_wgt_rd_0_data_bits_8_5(compute_io_wgt_rd_0_data_bits_8_5),
    .io_wgt_rd_0_data_bits_8_6(compute_io_wgt_rd_0_data_bits_8_6),
    .io_wgt_rd_0_data_bits_8_7(compute_io_wgt_rd_0_data_bits_8_7),
    .io_wgt_rd_0_data_bits_8_8(compute_io_wgt_rd_0_data_bits_8_8),
    .io_wgt_rd_0_data_bits_8_9(compute_io_wgt_rd_0_data_bits_8_9),
    .io_wgt_rd_0_data_bits_8_10(compute_io_wgt_rd_0_data_bits_8_10),
    .io_wgt_rd_0_data_bits_8_11(compute_io_wgt_rd_0_data_bits_8_11),
    .io_wgt_rd_0_data_bits_8_12(compute_io_wgt_rd_0_data_bits_8_12),
    .io_wgt_rd_0_data_bits_8_13(compute_io_wgt_rd_0_data_bits_8_13),
    .io_wgt_rd_0_data_bits_8_14(compute_io_wgt_rd_0_data_bits_8_14),
    .io_wgt_rd_0_data_bits_8_15(compute_io_wgt_rd_0_data_bits_8_15),
    .io_wgt_rd_0_data_bits_9_0(compute_io_wgt_rd_0_data_bits_9_0),
    .io_wgt_rd_0_data_bits_9_1(compute_io_wgt_rd_0_data_bits_9_1),
    .io_wgt_rd_0_data_bits_9_2(compute_io_wgt_rd_0_data_bits_9_2),
    .io_wgt_rd_0_data_bits_9_3(compute_io_wgt_rd_0_data_bits_9_3),
    .io_wgt_rd_0_data_bits_9_4(compute_io_wgt_rd_0_data_bits_9_4),
    .io_wgt_rd_0_data_bits_9_5(compute_io_wgt_rd_0_data_bits_9_5),
    .io_wgt_rd_0_data_bits_9_6(compute_io_wgt_rd_0_data_bits_9_6),
    .io_wgt_rd_0_data_bits_9_7(compute_io_wgt_rd_0_data_bits_9_7),
    .io_wgt_rd_0_data_bits_9_8(compute_io_wgt_rd_0_data_bits_9_8),
    .io_wgt_rd_0_data_bits_9_9(compute_io_wgt_rd_0_data_bits_9_9),
    .io_wgt_rd_0_data_bits_9_10(compute_io_wgt_rd_0_data_bits_9_10),
    .io_wgt_rd_0_data_bits_9_11(compute_io_wgt_rd_0_data_bits_9_11),
    .io_wgt_rd_0_data_bits_9_12(compute_io_wgt_rd_0_data_bits_9_12),
    .io_wgt_rd_0_data_bits_9_13(compute_io_wgt_rd_0_data_bits_9_13),
    .io_wgt_rd_0_data_bits_9_14(compute_io_wgt_rd_0_data_bits_9_14),
    .io_wgt_rd_0_data_bits_9_15(compute_io_wgt_rd_0_data_bits_9_15),
    .io_wgt_rd_0_data_bits_10_0(compute_io_wgt_rd_0_data_bits_10_0),
    .io_wgt_rd_0_data_bits_10_1(compute_io_wgt_rd_0_data_bits_10_1),
    .io_wgt_rd_0_data_bits_10_2(compute_io_wgt_rd_0_data_bits_10_2),
    .io_wgt_rd_0_data_bits_10_3(compute_io_wgt_rd_0_data_bits_10_3),
    .io_wgt_rd_0_data_bits_10_4(compute_io_wgt_rd_0_data_bits_10_4),
    .io_wgt_rd_0_data_bits_10_5(compute_io_wgt_rd_0_data_bits_10_5),
    .io_wgt_rd_0_data_bits_10_6(compute_io_wgt_rd_0_data_bits_10_6),
    .io_wgt_rd_0_data_bits_10_7(compute_io_wgt_rd_0_data_bits_10_7),
    .io_wgt_rd_0_data_bits_10_8(compute_io_wgt_rd_0_data_bits_10_8),
    .io_wgt_rd_0_data_bits_10_9(compute_io_wgt_rd_0_data_bits_10_9),
    .io_wgt_rd_0_data_bits_10_10(compute_io_wgt_rd_0_data_bits_10_10),
    .io_wgt_rd_0_data_bits_10_11(compute_io_wgt_rd_0_data_bits_10_11),
    .io_wgt_rd_0_data_bits_10_12(compute_io_wgt_rd_0_data_bits_10_12),
    .io_wgt_rd_0_data_bits_10_13(compute_io_wgt_rd_0_data_bits_10_13),
    .io_wgt_rd_0_data_bits_10_14(compute_io_wgt_rd_0_data_bits_10_14),
    .io_wgt_rd_0_data_bits_10_15(compute_io_wgt_rd_0_data_bits_10_15),
    .io_wgt_rd_0_data_bits_11_0(compute_io_wgt_rd_0_data_bits_11_0),
    .io_wgt_rd_0_data_bits_11_1(compute_io_wgt_rd_0_data_bits_11_1),
    .io_wgt_rd_0_data_bits_11_2(compute_io_wgt_rd_0_data_bits_11_2),
    .io_wgt_rd_0_data_bits_11_3(compute_io_wgt_rd_0_data_bits_11_3),
    .io_wgt_rd_0_data_bits_11_4(compute_io_wgt_rd_0_data_bits_11_4),
    .io_wgt_rd_0_data_bits_11_5(compute_io_wgt_rd_0_data_bits_11_5),
    .io_wgt_rd_0_data_bits_11_6(compute_io_wgt_rd_0_data_bits_11_6),
    .io_wgt_rd_0_data_bits_11_7(compute_io_wgt_rd_0_data_bits_11_7),
    .io_wgt_rd_0_data_bits_11_8(compute_io_wgt_rd_0_data_bits_11_8),
    .io_wgt_rd_0_data_bits_11_9(compute_io_wgt_rd_0_data_bits_11_9),
    .io_wgt_rd_0_data_bits_11_10(compute_io_wgt_rd_0_data_bits_11_10),
    .io_wgt_rd_0_data_bits_11_11(compute_io_wgt_rd_0_data_bits_11_11),
    .io_wgt_rd_0_data_bits_11_12(compute_io_wgt_rd_0_data_bits_11_12),
    .io_wgt_rd_0_data_bits_11_13(compute_io_wgt_rd_0_data_bits_11_13),
    .io_wgt_rd_0_data_bits_11_14(compute_io_wgt_rd_0_data_bits_11_14),
    .io_wgt_rd_0_data_bits_11_15(compute_io_wgt_rd_0_data_bits_11_15),
    .io_wgt_rd_0_data_bits_12_0(compute_io_wgt_rd_0_data_bits_12_0),
    .io_wgt_rd_0_data_bits_12_1(compute_io_wgt_rd_0_data_bits_12_1),
    .io_wgt_rd_0_data_bits_12_2(compute_io_wgt_rd_0_data_bits_12_2),
    .io_wgt_rd_0_data_bits_12_3(compute_io_wgt_rd_0_data_bits_12_3),
    .io_wgt_rd_0_data_bits_12_4(compute_io_wgt_rd_0_data_bits_12_4),
    .io_wgt_rd_0_data_bits_12_5(compute_io_wgt_rd_0_data_bits_12_5),
    .io_wgt_rd_0_data_bits_12_6(compute_io_wgt_rd_0_data_bits_12_6),
    .io_wgt_rd_0_data_bits_12_7(compute_io_wgt_rd_0_data_bits_12_7),
    .io_wgt_rd_0_data_bits_12_8(compute_io_wgt_rd_0_data_bits_12_8),
    .io_wgt_rd_0_data_bits_12_9(compute_io_wgt_rd_0_data_bits_12_9),
    .io_wgt_rd_0_data_bits_12_10(compute_io_wgt_rd_0_data_bits_12_10),
    .io_wgt_rd_0_data_bits_12_11(compute_io_wgt_rd_0_data_bits_12_11),
    .io_wgt_rd_0_data_bits_12_12(compute_io_wgt_rd_0_data_bits_12_12),
    .io_wgt_rd_0_data_bits_12_13(compute_io_wgt_rd_0_data_bits_12_13),
    .io_wgt_rd_0_data_bits_12_14(compute_io_wgt_rd_0_data_bits_12_14),
    .io_wgt_rd_0_data_bits_12_15(compute_io_wgt_rd_0_data_bits_12_15),
    .io_wgt_rd_0_data_bits_13_0(compute_io_wgt_rd_0_data_bits_13_0),
    .io_wgt_rd_0_data_bits_13_1(compute_io_wgt_rd_0_data_bits_13_1),
    .io_wgt_rd_0_data_bits_13_2(compute_io_wgt_rd_0_data_bits_13_2),
    .io_wgt_rd_0_data_bits_13_3(compute_io_wgt_rd_0_data_bits_13_3),
    .io_wgt_rd_0_data_bits_13_4(compute_io_wgt_rd_0_data_bits_13_4),
    .io_wgt_rd_0_data_bits_13_5(compute_io_wgt_rd_0_data_bits_13_5),
    .io_wgt_rd_0_data_bits_13_6(compute_io_wgt_rd_0_data_bits_13_6),
    .io_wgt_rd_0_data_bits_13_7(compute_io_wgt_rd_0_data_bits_13_7),
    .io_wgt_rd_0_data_bits_13_8(compute_io_wgt_rd_0_data_bits_13_8),
    .io_wgt_rd_0_data_bits_13_9(compute_io_wgt_rd_0_data_bits_13_9),
    .io_wgt_rd_0_data_bits_13_10(compute_io_wgt_rd_0_data_bits_13_10),
    .io_wgt_rd_0_data_bits_13_11(compute_io_wgt_rd_0_data_bits_13_11),
    .io_wgt_rd_0_data_bits_13_12(compute_io_wgt_rd_0_data_bits_13_12),
    .io_wgt_rd_0_data_bits_13_13(compute_io_wgt_rd_0_data_bits_13_13),
    .io_wgt_rd_0_data_bits_13_14(compute_io_wgt_rd_0_data_bits_13_14),
    .io_wgt_rd_0_data_bits_13_15(compute_io_wgt_rd_0_data_bits_13_15),
    .io_wgt_rd_0_data_bits_14_0(compute_io_wgt_rd_0_data_bits_14_0),
    .io_wgt_rd_0_data_bits_14_1(compute_io_wgt_rd_0_data_bits_14_1),
    .io_wgt_rd_0_data_bits_14_2(compute_io_wgt_rd_0_data_bits_14_2),
    .io_wgt_rd_0_data_bits_14_3(compute_io_wgt_rd_0_data_bits_14_3),
    .io_wgt_rd_0_data_bits_14_4(compute_io_wgt_rd_0_data_bits_14_4),
    .io_wgt_rd_0_data_bits_14_5(compute_io_wgt_rd_0_data_bits_14_5),
    .io_wgt_rd_0_data_bits_14_6(compute_io_wgt_rd_0_data_bits_14_6),
    .io_wgt_rd_0_data_bits_14_7(compute_io_wgt_rd_0_data_bits_14_7),
    .io_wgt_rd_0_data_bits_14_8(compute_io_wgt_rd_0_data_bits_14_8),
    .io_wgt_rd_0_data_bits_14_9(compute_io_wgt_rd_0_data_bits_14_9),
    .io_wgt_rd_0_data_bits_14_10(compute_io_wgt_rd_0_data_bits_14_10),
    .io_wgt_rd_0_data_bits_14_11(compute_io_wgt_rd_0_data_bits_14_11),
    .io_wgt_rd_0_data_bits_14_12(compute_io_wgt_rd_0_data_bits_14_12),
    .io_wgt_rd_0_data_bits_14_13(compute_io_wgt_rd_0_data_bits_14_13),
    .io_wgt_rd_0_data_bits_14_14(compute_io_wgt_rd_0_data_bits_14_14),
    .io_wgt_rd_0_data_bits_14_15(compute_io_wgt_rd_0_data_bits_14_15),
    .io_wgt_rd_0_data_bits_15_0(compute_io_wgt_rd_0_data_bits_15_0),
    .io_wgt_rd_0_data_bits_15_1(compute_io_wgt_rd_0_data_bits_15_1),
    .io_wgt_rd_0_data_bits_15_2(compute_io_wgt_rd_0_data_bits_15_2),
    .io_wgt_rd_0_data_bits_15_3(compute_io_wgt_rd_0_data_bits_15_3),
    .io_wgt_rd_0_data_bits_15_4(compute_io_wgt_rd_0_data_bits_15_4),
    .io_wgt_rd_0_data_bits_15_5(compute_io_wgt_rd_0_data_bits_15_5),
    .io_wgt_rd_0_data_bits_15_6(compute_io_wgt_rd_0_data_bits_15_6),
    .io_wgt_rd_0_data_bits_15_7(compute_io_wgt_rd_0_data_bits_15_7),
    .io_wgt_rd_0_data_bits_15_8(compute_io_wgt_rd_0_data_bits_15_8),
    .io_wgt_rd_0_data_bits_15_9(compute_io_wgt_rd_0_data_bits_15_9),
    .io_wgt_rd_0_data_bits_15_10(compute_io_wgt_rd_0_data_bits_15_10),
    .io_wgt_rd_0_data_bits_15_11(compute_io_wgt_rd_0_data_bits_15_11),
    .io_wgt_rd_0_data_bits_15_12(compute_io_wgt_rd_0_data_bits_15_12),
    .io_wgt_rd_0_data_bits_15_13(compute_io_wgt_rd_0_data_bits_15_13),
    .io_wgt_rd_0_data_bits_15_14(compute_io_wgt_rd_0_data_bits_15_14),
    .io_wgt_rd_0_data_bits_15_15(compute_io_wgt_rd_0_data_bits_15_15),
    .io_wgt_rd_0_data_bits_16_0(compute_io_wgt_rd_0_data_bits_16_0),
    .io_wgt_rd_0_data_bits_16_1(compute_io_wgt_rd_0_data_bits_16_1),
    .io_wgt_rd_0_data_bits_16_2(compute_io_wgt_rd_0_data_bits_16_2),
    .io_wgt_rd_0_data_bits_16_3(compute_io_wgt_rd_0_data_bits_16_3),
    .io_wgt_rd_0_data_bits_16_4(compute_io_wgt_rd_0_data_bits_16_4),
    .io_wgt_rd_0_data_bits_16_5(compute_io_wgt_rd_0_data_bits_16_5),
    .io_wgt_rd_0_data_bits_16_6(compute_io_wgt_rd_0_data_bits_16_6),
    .io_wgt_rd_0_data_bits_16_7(compute_io_wgt_rd_0_data_bits_16_7),
    .io_wgt_rd_0_data_bits_16_8(compute_io_wgt_rd_0_data_bits_16_8),
    .io_wgt_rd_0_data_bits_16_9(compute_io_wgt_rd_0_data_bits_16_9),
    .io_wgt_rd_0_data_bits_16_10(compute_io_wgt_rd_0_data_bits_16_10),
    .io_wgt_rd_0_data_bits_16_11(compute_io_wgt_rd_0_data_bits_16_11),
    .io_wgt_rd_0_data_bits_16_12(compute_io_wgt_rd_0_data_bits_16_12),
    .io_wgt_rd_0_data_bits_16_13(compute_io_wgt_rd_0_data_bits_16_13),
    .io_wgt_rd_0_data_bits_16_14(compute_io_wgt_rd_0_data_bits_16_14),
    .io_wgt_rd_0_data_bits_16_15(compute_io_wgt_rd_0_data_bits_16_15),
    .io_wgt_rd_0_data_bits_17_0(compute_io_wgt_rd_0_data_bits_17_0),
    .io_wgt_rd_0_data_bits_17_1(compute_io_wgt_rd_0_data_bits_17_1),
    .io_wgt_rd_0_data_bits_17_2(compute_io_wgt_rd_0_data_bits_17_2),
    .io_wgt_rd_0_data_bits_17_3(compute_io_wgt_rd_0_data_bits_17_3),
    .io_wgt_rd_0_data_bits_17_4(compute_io_wgt_rd_0_data_bits_17_4),
    .io_wgt_rd_0_data_bits_17_5(compute_io_wgt_rd_0_data_bits_17_5),
    .io_wgt_rd_0_data_bits_17_6(compute_io_wgt_rd_0_data_bits_17_6),
    .io_wgt_rd_0_data_bits_17_7(compute_io_wgt_rd_0_data_bits_17_7),
    .io_wgt_rd_0_data_bits_17_8(compute_io_wgt_rd_0_data_bits_17_8),
    .io_wgt_rd_0_data_bits_17_9(compute_io_wgt_rd_0_data_bits_17_9),
    .io_wgt_rd_0_data_bits_17_10(compute_io_wgt_rd_0_data_bits_17_10),
    .io_wgt_rd_0_data_bits_17_11(compute_io_wgt_rd_0_data_bits_17_11),
    .io_wgt_rd_0_data_bits_17_12(compute_io_wgt_rd_0_data_bits_17_12),
    .io_wgt_rd_0_data_bits_17_13(compute_io_wgt_rd_0_data_bits_17_13),
    .io_wgt_rd_0_data_bits_17_14(compute_io_wgt_rd_0_data_bits_17_14),
    .io_wgt_rd_0_data_bits_17_15(compute_io_wgt_rd_0_data_bits_17_15),
    .io_wgt_rd_0_data_bits_18_0(compute_io_wgt_rd_0_data_bits_18_0),
    .io_wgt_rd_0_data_bits_18_1(compute_io_wgt_rd_0_data_bits_18_1),
    .io_wgt_rd_0_data_bits_18_2(compute_io_wgt_rd_0_data_bits_18_2),
    .io_wgt_rd_0_data_bits_18_3(compute_io_wgt_rd_0_data_bits_18_3),
    .io_wgt_rd_0_data_bits_18_4(compute_io_wgt_rd_0_data_bits_18_4),
    .io_wgt_rd_0_data_bits_18_5(compute_io_wgt_rd_0_data_bits_18_5),
    .io_wgt_rd_0_data_bits_18_6(compute_io_wgt_rd_0_data_bits_18_6),
    .io_wgt_rd_0_data_bits_18_7(compute_io_wgt_rd_0_data_bits_18_7),
    .io_wgt_rd_0_data_bits_18_8(compute_io_wgt_rd_0_data_bits_18_8),
    .io_wgt_rd_0_data_bits_18_9(compute_io_wgt_rd_0_data_bits_18_9),
    .io_wgt_rd_0_data_bits_18_10(compute_io_wgt_rd_0_data_bits_18_10),
    .io_wgt_rd_0_data_bits_18_11(compute_io_wgt_rd_0_data_bits_18_11),
    .io_wgt_rd_0_data_bits_18_12(compute_io_wgt_rd_0_data_bits_18_12),
    .io_wgt_rd_0_data_bits_18_13(compute_io_wgt_rd_0_data_bits_18_13),
    .io_wgt_rd_0_data_bits_18_14(compute_io_wgt_rd_0_data_bits_18_14),
    .io_wgt_rd_0_data_bits_18_15(compute_io_wgt_rd_0_data_bits_18_15),
    .io_wgt_rd_0_data_bits_19_0(compute_io_wgt_rd_0_data_bits_19_0),
    .io_wgt_rd_0_data_bits_19_1(compute_io_wgt_rd_0_data_bits_19_1),
    .io_wgt_rd_0_data_bits_19_2(compute_io_wgt_rd_0_data_bits_19_2),
    .io_wgt_rd_0_data_bits_19_3(compute_io_wgt_rd_0_data_bits_19_3),
    .io_wgt_rd_0_data_bits_19_4(compute_io_wgt_rd_0_data_bits_19_4),
    .io_wgt_rd_0_data_bits_19_5(compute_io_wgt_rd_0_data_bits_19_5),
    .io_wgt_rd_0_data_bits_19_6(compute_io_wgt_rd_0_data_bits_19_6),
    .io_wgt_rd_0_data_bits_19_7(compute_io_wgt_rd_0_data_bits_19_7),
    .io_wgt_rd_0_data_bits_19_8(compute_io_wgt_rd_0_data_bits_19_8),
    .io_wgt_rd_0_data_bits_19_9(compute_io_wgt_rd_0_data_bits_19_9),
    .io_wgt_rd_0_data_bits_19_10(compute_io_wgt_rd_0_data_bits_19_10),
    .io_wgt_rd_0_data_bits_19_11(compute_io_wgt_rd_0_data_bits_19_11),
    .io_wgt_rd_0_data_bits_19_12(compute_io_wgt_rd_0_data_bits_19_12),
    .io_wgt_rd_0_data_bits_19_13(compute_io_wgt_rd_0_data_bits_19_13),
    .io_wgt_rd_0_data_bits_19_14(compute_io_wgt_rd_0_data_bits_19_14),
    .io_wgt_rd_0_data_bits_19_15(compute_io_wgt_rd_0_data_bits_19_15),
    .io_wgt_rd_0_data_bits_20_0(compute_io_wgt_rd_0_data_bits_20_0),
    .io_wgt_rd_0_data_bits_20_1(compute_io_wgt_rd_0_data_bits_20_1),
    .io_wgt_rd_0_data_bits_20_2(compute_io_wgt_rd_0_data_bits_20_2),
    .io_wgt_rd_0_data_bits_20_3(compute_io_wgt_rd_0_data_bits_20_3),
    .io_wgt_rd_0_data_bits_20_4(compute_io_wgt_rd_0_data_bits_20_4),
    .io_wgt_rd_0_data_bits_20_5(compute_io_wgt_rd_0_data_bits_20_5),
    .io_wgt_rd_0_data_bits_20_6(compute_io_wgt_rd_0_data_bits_20_6),
    .io_wgt_rd_0_data_bits_20_7(compute_io_wgt_rd_0_data_bits_20_7),
    .io_wgt_rd_0_data_bits_20_8(compute_io_wgt_rd_0_data_bits_20_8),
    .io_wgt_rd_0_data_bits_20_9(compute_io_wgt_rd_0_data_bits_20_9),
    .io_wgt_rd_0_data_bits_20_10(compute_io_wgt_rd_0_data_bits_20_10),
    .io_wgt_rd_0_data_bits_20_11(compute_io_wgt_rd_0_data_bits_20_11),
    .io_wgt_rd_0_data_bits_20_12(compute_io_wgt_rd_0_data_bits_20_12),
    .io_wgt_rd_0_data_bits_20_13(compute_io_wgt_rd_0_data_bits_20_13),
    .io_wgt_rd_0_data_bits_20_14(compute_io_wgt_rd_0_data_bits_20_14),
    .io_wgt_rd_0_data_bits_20_15(compute_io_wgt_rd_0_data_bits_20_15),
    .io_wgt_rd_0_data_bits_21_0(compute_io_wgt_rd_0_data_bits_21_0),
    .io_wgt_rd_0_data_bits_21_1(compute_io_wgt_rd_0_data_bits_21_1),
    .io_wgt_rd_0_data_bits_21_2(compute_io_wgt_rd_0_data_bits_21_2),
    .io_wgt_rd_0_data_bits_21_3(compute_io_wgt_rd_0_data_bits_21_3),
    .io_wgt_rd_0_data_bits_21_4(compute_io_wgt_rd_0_data_bits_21_4),
    .io_wgt_rd_0_data_bits_21_5(compute_io_wgt_rd_0_data_bits_21_5),
    .io_wgt_rd_0_data_bits_21_6(compute_io_wgt_rd_0_data_bits_21_6),
    .io_wgt_rd_0_data_bits_21_7(compute_io_wgt_rd_0_data_bits_21_7),
    .io_wgt_rd_0_data_bits_21_8(compute_io_wgt_rd_0_data_bits_21_8),
    .io_wgt_rd_0_data_bits_21_9(compute_io_wgt_rd_0_data_bits_21_9),
    .io_wgt_rd_0_data_bits_21_10(compute_io_wgt_rd_0_data_bits_21_10),
    .io_wgt_rd_0_data_bits_21_11(compute_io_wgt_rd_0_data_bits_21_11),
    .io_wgt_rd_0_data_bits_21_12(compute_io_wgt_rd_0_data_bits_21_12),
    .io_wgt_rd_0_data_bits_21_13(compute_io_wgt_rd_0_data_bits_21_13),
    .io_wgt_rd_0_data_bits_21_14(compute_io_wgt_rd_0_data_bits_21_14),
    .io_wgt_rd_0_data_bits_21_15(compute_io_wgt_rd_0_data_bits_21_15),
    .io_wgt_rd_0_data_bits_22_0(compute_io_wgt_rd_0_data_bits_22_0),
    .io_wgt_rd_0_data_bits_22_1(compute_io_wgt_rd_0_data_bits_22_1),
    .io_wgt_rd_0_data_bits_22_2(compute_io_wgt_rd_0_data_bits_22_2),
    .io_wgt_rd_0_data_bits_22_3(compute_io_wgt_rd_0_data_bits_22_3),
    .io_wgt_rd_0_data_bits_22_4(compute_io_wgt_rd_0_data_bits_22_4),
    .io_wgt_rd_0_data_bits_22_5(compute_io_wgt_rd_0_data_bits_22_5),
    .io_wgt_rd_0_data_bits_22_6(compute_io_wgt_rd_0_data_bits_22_6),
    .io_wgt_rd_0_data_bits_22_7(compute_io_wgt_rd_0_data_bits_22_7),
    .io_wgt_rd_0_data_bits_22_8(compute_io_wgt_rd_0_data_bits_22_8),
    .io_wgt_rd_0_data_bits_22_9(compute_io_wgt_rd_0_data_bits_22_9),
    .io_wgt_rd_0_data_bits_22_10(compute_io_wgt_rd_0_data_bits_22_10),
    .io_wgt_rd_0_data_bits_22_11(compute_io_wgt_rd_0_data_bits_22_11),
    .io_wgt_rd_0_data_bits_22_12(compute_io_wgt_rd_0_data_bits_22_12),
    .io_wgt_rd_0_data_bits_22_13(compute_io_wgt_rd_0_data_bits_22_13),
    .io_wgt_rd_0_data_bits_22_14(compute_io_wgt_rd_0_data_bits_22_14),
    .io_wgt_rd_0_data_bits_22_15(compute_io_wgt_rd_0_data_bits_22_15),
    .io_wgt_rd_0_data_bits_23_0(compute_io_wgt_rd_0_data_bits_23_0),
    .io_wgt_rd_0_data_bits_23_1(compute_io_wgt_rd_0_data_bits_23_1),
    .io_wgt_rd_0_data_bits_23_2(compute_io_wgt_rd_0_data_bits_23_2),
    .io_wgt_rd_0_data_bits_23_3(compute_io_wgt_rd_0_data_bits_23_3),
    .io_wgt_rd_0_data_bits_23_4(compute_io_wgt_rd_0_data_bits_23_4),
    .io_wgt_rd_0_data_bits_23_5(compute_io_wgt_rd_0_data_bits_23_5),
    .io_wgt_rd_0_data_bits_23_6(compute_io_wgt_rd_0_data_bits_23_6),
    .io_wgt_rd_0_data_bits_23_7(compute_io_wgt_rd_0_data_bits_23_7),
    .io_wgt_rd_0_data_bits_23_8(compute_io_wgt_rd_0_data_bits_23_8),
    .io_wgt_rd_0_data_bits_23_9(compute_io_wgt_rd_0_data_bits_23_9),
    .io_wgt_rd_0_data_bits_23_10(compute_io_wgt_rd_0_data_bits_23_10),
    .io_wgt_rd_0_data_bits_23_11(compute_io_wgt_rd_0_data_bits_23_11),
    .io_wgt_rd_0_data_bits_23_12(compute_io_wgt_rd_0_data_bits_23_12),
    .io_wgt_rd_0_data_bits_23_13(compute_io_wgt_rd_0_data_bits_23_13),
    .io_wgt_rd_0_data_bits_23_14(compute_io_wgt_rd_0_data_bits_23_14),
    .io_wgt_rd_0_data_bits_23_15(compute_io_wgt_rd_0_data_bits_23_15),
    .io_wgt_rd_0_data_bits_24_0(compute_io_wgt_rd_0_data_bits_24_0),
    .io_wgt_rd_0_data_bits_24_1(compute_io_wgt_rd_0_data_bits_24_1),
    .io_wgt_rd_0_data_bits_24_2(compute_io_wgt_rd_0_data_bits_24_2),
    .io_wgt_rd_0_data_bits_24_3(compute_io_wgt_rd_0_data_bits_24_3),
    .io_wgt_rd_0_data_bits_24_4(compute_io_wgt_rd_0_data_bits_24_4),
    .io_wgt_rd_0_data_bits_24_5(compute_io_wgt_rd_0_data_bits_24_5),
    .io_wgt_rd_0_data_bits_24_6(compute_io_wgt_rd_0_data_bits_24_6),
    .io_wgt_rd_0_data_bits_24_7(compute_io_wgt_rd_0_data_bits_24_7),
    .io_wgt_rd_0_data_bits_24_8(compute_io_wgt_rd_0_data_bits_24_8),
    .io_wgt_rd_0_data_bits_24_9(compute_io_wgt_rd_0_data_bits_24_9),
    .io_wgt_rd_0_data_bits_24_10(compute_io_wgt_rd_0_data_bits_24_10),
    .io_wgt_rd_0_data_bits_24_11(compute_io_wgt_rd_0_data_bits_24_11),
    .io_wgt_rd_0_data_bits_24_12(compute_io_wgt_rd_0_data_bits_24_12),
    .io_wgt_rd_0_data_bits_24_13(compute_io_wgt_rd_0_data_bits_24_13),
    .io_wgt_rd_0_data_bits_24_14(compute_io_wgt_rd_0_data_bits_24_14),
    .io_wgt_rd_0_data_bits_24_15(compute_io_wgt_rd_0_data_bits_24_15),
    .io_wgt_rd_0_data_bits_25_0(compute_io_wgt_rd_0_data_bits_25_0),
    .io_wgt_rd_0_data_bits_25_1(compute_io_wgt_rd_0_data_bits_25_1),
    .io_wgt_rd_0_data_bits_25_2(compute_io_wgt_rd_0_data_bits_25_2),
    .io_wgt_rd_0_data_bits_25_3(compute_io_wgt_rd_0_data_bits_25_3),
    .io_wgt_rd_0_data_bits_25_4(compute_io_wgt_rd_0_data_bits_25_4),
    .io_wgt_rd_0_data_bits_25_5(compute_io_wgt_rd_0_data_bits_25_5),
    .io_wgt_rd_0_data_bits_25_6(compute_io_wgt_rd_0_data_bits_25_6),
    .io_wgt_rd_0_data_bits_25_7(compute_io_wgt_rd_0_data_bits_25_7),
    .io_wgt_rd_0_data_bits_25_8(compute_io_wgt_rd_0_data_bits_25_8),
    .io_wgt_rd_0_data_bits_25_9(compute_io_wgt_rd_0_data_bits_25_9),
    .io_wgt_rd_0_data_bits_25_10(compute_io_wgt_rd_0_data_bits_25_10),
    .io_wgt_rd_0_data_bits_25_11(compute_io_wgt_rd_0_data_bits_25_11),
    .io_wgt_rd_0_data_bits_25_12(compute_io_wgt_rd_0_data_bits_25_12),
    .io_wgt_rd_0_data_bits_25_13(compute_io_wgt_rd_0_data_bits_25_13),
    .io_wgt_rd_0_data_bits_25_14(compute_io_wgt_rd_0_data_bits_25_14),
    .io_wgt_rd_0_data_bits_25_15(compute_io_wgt_rd_0_data_bits_25_15),
    .io_wgt_rd_0_data_bits_26_0(compute_io_wgt_rd_0_data_bits_26_0),
    .io_wgt_rd_0_data_bits_26_1(compute_io_wgt_rd_0_data_bits_26_1),
    .io_wgt_rd_0_data_bits_26_2(compute_io_wgt_rd_0_data_bits_26_2),
    .io_wgt_rd_0_data_bits_26_3(compute_io_wgt_rd_0_data_bits_26_3),
    .io_wgt_rd_0_data_bits_26_4(compute_io_wgt_rd_0_data_bits_26_4),
    .io_wgt_rd_0_data_bits_26_5(compute_io_wgt_rd_0_data_bits_26_5),
    .io_wgt_rd_0_data_bits_26_6(compute_io_wgt_rd_0_data_bits_26_6),
    .io_wgt_rd_0_data_bits_26_7(compute_io_wgt_rd_0_data_bits_26_7),
    .io_wgt_rd_0_data_bits_26_8(compute_io_wgt_rd_0_data_bits_26_8),
    .io_wgt_rd_0_data_bits_26_9(compute_io_wgt_rd_0_data_bits_26_9),
    .io_wgt_rd_0_data_bits_26_10(compute_io_wgt_rd_0_data_bits_26_10),
    .io_wgt_rd_0_data_bits_26_11(compute_io_wgt_rd_0_data_bits_26_11),
    .io_wgt_rd_0_data_bits_26_12(compute_io_wgt_rd_0_data_bits_26_12),
    .io_wgt_rd_0_data_bits_26_13(compute_io_wgt_rd_0_data_bits_26_13),
    .io_wgt_rd_0_data_bits_26_14(compute_io_wgt_rd_0_data_bits_26_14),
    .io_wgt_rd_0_data_bits_26_15(compute_io_wgt_rd_0_data_bits_26_15),
    .io_wgt_rd_0_data_bits_27_0(compute_io_wgt_rd_0_data_bits_27_0),
    .io_wgt_rd_0_data_bits_27_1(compute_io_wgt_rd_0_data_bits_27_1),
    .io_wgt_rd_0_data_bits_27_2(compute_io_wgt_rd_0_data_bits_27_2),
    .io_wgt_rd_0_data_bits_27_3(compute_io_wgt_rd_0_data_bits_27_3),
    .io_wgt_rd_0_data_bits_27_4(compute_io_wgt_rd_0_data_bits_27_4),
    .io_wgt_rd_0_data_bits_27_5(compute_io_wgt_rd_0_data_bits_27_5),
    .io_wgt_rd_0_data_bits_27_6(compute_io_wgt_rd_0_data_bits_27_6),
    .io_wgt_rd_0_data_bits_27_7(compute_io_wgt_rd_0_data_bits_27_7),
    .io_wgt_rd_0_data_bits_27_8(compute_io_wgt_rd_0_data_bits_27_8),
    .io_wgt_rd_0_data_bits_27_9(compute_io_wgt_rd_0_data_bits_27_9),
    .io_wgt_rd_0_data_bits_27_10(compute_io_wgt_rd_0_data_bits_27_10),
    .io_wgt_rd_0_data_bits_27_11(compute_io_wgt_rd_0_data_bits_27_11),
    .io_wgt_rd_0_data_bits_27_12(compute_io_wgt_rd_0_data_bits_27_12),
    .io_wgt_rd_0_data_bits_27_13(compute_io_wgt_rd_0_data_bits_27_13),
    .io_wgt_rd_0_data_bits_27_14(compute_io_wgt_rd_0_data_bits_27_14),
    .io_wgt_rd_0_data_bits_27_15(compute_io_wgt_rd_0_data_bits_27_15),
    .io_wgt_rd_0_data_bits_28_0(compute_io_wgt_rd_0_data_bits_28_0),
    .io_wgt_rd_0_data_bits_28_1(compute_io_wgt_rd_0_data_bits_28_1),
    .io_wgt_rd_0_data_bits_28_2(compute_io_wgt_rd_0_data_bits_28_2),
    .io_wgt_rd_0_data_bits_28_3(compute_io_wgt_rd_0_data_bits_28_3),
    .io_wgt_rd_0_data_bits_28_4(compute_io_wgt_rd_0_data_bits_28_4),
    .io_wgt_rd_0_data_bits_28_5(compute_io_wgt_rd_0_data_bits_28_5),
    .io_wgt_rd_0_data_bits_28_6(compute_io_wgt_rd_0_data_bits_28_6),
    .io_wgt_rd_0_data_bits_28_7(compute_io_wgt_rd_0_data_bits_28_7),
    .io_wgt_rd_0_data_bits_28_8(compute_io_wgt_rd_0_data_bits_28_8),
    .io_wgt_rd_0_data_bits_28_9(compute_io_wgt_rd_0_data_bits_28_9),
    .io_wgt_rd_0_data_bits_28_10(compute_io_wgt_rd_0_data_bits_28_10),
    .io_wgt_rd_0_data_bits_28_11(compute_io_wgt_rd_0_data_bits_28_11),
    .io_wgt_rd_0_data_bits_28_12(compute_io_wgt_rd_0_data_bits_28_12),
    .io_wgt_rd_0_data_bits_28_13(compute_io_wgt_rd_0_data_bits_28_13),
    .io_wgt_rd_0_data_bits_28_14(compute_io_wgt_rd_0_data_bits_28_14),
    .io_wgt_rd_0_data_bits_28_15(compute_io_wgt_rd_0_data_bits_28_15),
    .io_wgt_rd_0_data_bits_29_0(compute_io_wgt_rd_0_data_bits_29_0),
    .io_wgt_rd_0_data_bits_29_1(compute_io_wgt_rd_0_data_bits_29_1),
    .io_wgt_rd_0_data_bits_29_2(compute_io_wgt_rd_0_data_bits_29_2),
    .io_wgt_rd_0_data_bits_29_3(compute_io_wgt_rd_0_data_bits_29_3),
    .io_wgt_rd_0_data_bits_29_4(compute_io_wgt_rd_0_data_bits_29_4),
    .io_wgt_rd_0_data_bits_29_5(compute_io_wgt_rd_0_data_bits_29_5),
    .io_wgt_rd_0_data_bits_29_6(compute_io_wgt_rd_0_data_bits_29_6),
    .io_wgt_rd_0_data_bits_29_7(compute_io_wgt_rd_0_data_bits_29_7),
    .io_wgt_rd_0_data_bits_29_8(compute_io_wgt_rd_0_data_bits_29_8),
    .io_wgt_rd_0_data_bits_29_9(compute_io_wgt_rd_0_data_bits_29_9),
    .io_wgt_rd_0_data_bits_29_10(compute_io_wgt_rd_0_data_bits_29_10),
    .io_wgt_rd_0_data_bits_29_11(compute_io_wgt_rd_0_data_bits_29_11),
    .io_wgt_rd_0_data_bits_29_12(compute_io_wgt_rd_0_data_bits_29_12),
    .io_wgt_rd_0_data_bits_29_13(compute_io_wgt_rd_0_data_bits_29_13),
    .io_wgt_rd_0_data_bits_29_14(compute_io_wgt_rd_0_data_bits_29_14),
    .io_wgt_rd_0_data_bits_29_15(compute_io_wgt_rd_0_data_bits_29_15),
    .io_wgt_rd_0_data_bits_30_0(compute_io_wgt_rd_0_data_bits_30_0),
    .io_wgt_rd_0_data_bits_30_1(compute_io_wgt_rd_0_data_bits_30_1),
    .io_wgt_rd_0_data_bits_30_2(compute_io_wgt_rd_0_data_bits_30_2),
    .io_wgt_rd_0_data_bits_30_3(compute_io_wgt_rd_0_data_bits_30_3),
    .io_wgt_rd_0_data_bits_30_4(compute_io_wgt_rd_0_data_bits_30_4),
    .io_wgt_rd_0_data_bits_30_5(compute_io_wgt_rd_0_data_bits_30_5),
    .io_wgt_rd_0_data_bits_30_6(compute_io_wgt_rd_0_data_bits_30_6),
    .io_wgt_rd_0_data_bits_30_7(compute_io_wgt_rd_0_data_bits_30_7),
    .io_wgt_rd_0_data_bits_30_8(compute_io_wgt_rd_0_data_bits_30_8),
    .io_wgt_rd_0_data_bits_30_9(compute_io_wgt_rd_0_data_bits_30_9),
    .io_wgt_rd_0_data_bits_30_10(compute_io_wgt_rd_0_data_bits_30_10),
    .io_wgt_rd_0_data_bits_30_11(compute_io_wgt_rd_0_data_bits_30_11),
    .io_wgt_rd_0_data_bits_30_12(compute_io_wgt_rd_0_data_bits_30_12),
    .io_wgt_rd_0_data_bits_30_13(compute_io_wgt_rd_0_data_bits_30_13),
    .io_wgt_rd_0_data_bits_30_14(compute_io_wgt_rd_0_data_bits_30_14),
    .io_wgt_rd_0_data_bits_30_15(compute_io_wgt_rd_0_data_bits_30_15),
    .io_wgt_rd_0_data_bits_31_0(compute_io_wgt_rd_0_data_bits_31_0),
    .io_wgt_rd_0_data_bits_31_1(compute_io_wgt_rd_0_data_bits_31_1),
    .io_wgt_rd_0_data_bits_31_2(compute_io_wgt_rd_0_data_bits_31_2),
    .io_wgt_rd_0_data_bits_31_3(compute_io_wgt_rd_0_data_bits_31_3),
    .io_wgt_rd_0_data_bits_31_4(compute_io_wgt_rd_0_data_bits_31_4),
    .io_wgt_rd_0_data_bits_31_5(compute_io_wgt_rd_0_data_bits_31_5),
    .io_wgt_rd_0_data_bits_31_6(compute_io_wgt_rd_0_data_bits_31_6),
    .io_wgt_rd_0_data_bits_31_7(compute_io_wgt_rd_0_data_bits_31_7),
    .io_wgt_rd_0_data_bits_31_8(compute_io_wgt_rd_0_data_bits_31_8),
    .io_wgt_rd_0_data_bits_31_9(compute_io_wgt_rd_0_data_bits_31_9),
    .io_wgt_rd_0_data_bits_31_10(compute_io_wgt_rd_0_data_bits_31_10),
    .io_wgt_rd_0_data_bits_31_11(compute_io_wgt_rd_0_data_bits_31_11),
    .io_wgt_rd_0_data_bits_31_12(compute_io_wgt_rd_0_data_bits_31_12),
    .io_wgt_rd_0_data_bits_31_13(compute_io_wgt_rd_0_data_bits_31_13),
    .io_wgt_rd_0_data_bits_31_14(compute_io_wgt_rd_0_data_bits_31_14),
    .io_wgt_rd_0_data_bits_31_15(compute_io_wgt_rd_0_data_bits_31_15),
    .io_out_wr_0_valid(compute_io_out_wr_0_valid),
    .io_out_wr_0_bits_idx(compute_io_out_wr_0_bits_idx),
    .io_out_wr_0_bits_data_0_0(compute_io_out_wr_0_bits_data_0_0),
    .io_out_wr_0_bits_data_0_1(compute_io_out_wr_0_bits_data_0_1),
    .io_out_wr_0_bits_data_0_2(compute_io_out_wr_0_bits_data_0_2),
    .io_out_wr_0_bits_data_0_3(compute_io_out_wr_0_bits_data_0_3),
    .io_out_wr_0_bits_data_0_4(compute_io_out_wr_0_bits_data_0_4),
    .io_out_wr_0_bits_data_0_5(compute_io_out_wr_0_bits_data_0_5),
    .io_out_wr_0_bits_data_0_6(compute_io_out_wr_0_bits_data_0_6),
    .io_out_wr_0_bits_data_0_7(compute_io_out_wr_0_bits_data_0_7),
    .io_out_wr_0_bits_data_0_8(compute_io_out_wr_0_bits_data_0_8),
    .io_out_wr_0_bits_data_0_9(compute_io_out_wr_0_bits_data_0_9),
    .io_out_wr_0_bits_data_0_10(compute_io_out_wr_0_bits_data_0_10),
    .io_out_wr_0_bits_data_0_11(compute_io_out_wr_0_bits_data_0_11),
    .io_out_wr_0_bits_data_0_12(compute_io_out_wr_0_bits_data_0_12),
    .io_out_wr_0_bits_data_0_13(compute_io_out_wr_0_bits_data_0_13),
    .io_out_wr_0_bits_data_0_14(compute_io_out_wr_0_bits_data_0_14),
    .io_out_wr_0_bits_data_0_15(compute_io_out_wr_0_bits_data_0_15),
    .io_out_wr_0_bits_data_0_16(compute_io_out_wr_0_bits_data_0_16),
    .io_out_wr_0_bits_data_0_17(compute_io_out_wr_0_bits_data_0_17),
    .io_out_wr_0_bits_data_0_18(compute_io_out_wr_0_bits_data_0_18),
    .io_out_wr_0_bits_data_0_19(compute_io_out_wr_0_bits_data_0_19),
    .io_out_wr_0_bits_data_0_20(compute_io_out_wr_0_bits_data_0_20),
    .io_out_wr_0_bits_data_0_21(compute_io_out_wr_0_bits_data_0_21),
    .io_out_wr_0_bits_data_0_22(compute_io_out_wr_0_bits_data_0_22),
    .io_out_wr_0_bits_data_0_23(compute_io_out_wr_0_bits_data_0_23),
    .io_out_wr_0_bits_data_0_24(compute_io_out_wr_0_bits_data_0_24),
    .io_out_wr_0_bits_data_0_25(compute_io_out_wr_0_bits_data_0_25),
    .io_out_wr_0_bits_data_0_26(compute_io_out_wr_0_bits_data_0_26),
    .io_out_wr_0_bits_data_0_27(compute_io_out_wr_0_bits_data_0_27),
    .io_out_wr_0_bits_data_0_28(compute_io_out_wr_0_bits_data_0_28),
    .io_out_wr_0_bits_data_0_29(compute_io_out_wr_0_bits_data_0_29),
    .io_out_wr_0_bits_data_0_30(compute_io_out_wr_0_bits_data_0_30),
    .io_out_wr_0_bits_data_0_31(compute_io_out_wr_0_bits_data_0_31),
    .io_finish(compute_io_finish),
    .io_acc_wr_event(compute_io_acc_wr_event)
  );
  Store store ( // @[Core.scala 70:21]
    .clock(store_clock),
    .reset(store_reset),
    .io_i_post(store_io_i_post),
    .io_o_post(store_io_o_post),
    .io_inst_ready(store_io_inst_ready),
    .io_inst_valid(store_io_inst_valid),
    .io_inst_bits(store_io_inst_bits),
    .io_out_baddr(store_io_out_baddr),
    .io_vme_wr_cmd_ready(store_io_vme_wr_cmd_ready),
    .io_vme_wr_cmd_valid(store_io_vme_wr_cmd_valid),
    .io_vme_wr_cmd_bits_addr(store_io_vme_wr_cmd_bits_addr),
    .io_vme_wr_cmd_bits_len(store_io_vme_wr_cmd_bits_len),
    .io_vme_wr_data_ready(store_io_vme_wr_data_ready),
    .io_vme_wr_data_valid(store_io_vme_wr_data_valid),
    .io_vme_wr_data_bits_data(store_io_vme_wr_data_bits_data),
    .io_vme_wr_ack(store_io_vme_wr_ack),
    .io_out_wr_0_valid(store_io_out_wr_0_valid),
    .io_out_wr_0_bits_idx(store_io_out_wr_0_bits_idx),
    .io_out_wr_0_bits_data_0_0(store_io_out_wr_0_bits_data_0_0),
    .io_out_wr_0_bits_data_0_1(store_io_out_wr_0_bits_data_0_1),
    .io_out_wr_0_bits_data_0_2(store_io_out_wr_0_bits_data_0_2),
    .io_out_wr_0_bits_data_0_3(store_io_out_wr_0_bits_data_0_3),
    .io_out_wr_0_bits_data_0_4(store_io_out_wr_0_bits_data_0_4),
    .io_out_wr_0_bits_data_0_5(store_io_out_wr_0_bits_data_0_5),
    .io_out_wr_0_bits_data_0_6(store_io_out_wr_0_bits_data_0_6),
    .io_out_wr_0_bits_data_0_7(store_io_out_wr_0_bits_data_0_7),
    .io_out_wr_0_bits_data_0_8(store_io_out_wr_0_bits_data_0_8),
    .io_out_wr_0_bits_data_0_9(store_io_out_wr_0_bits_data_0_9),
    .io_out_wr_0_bits_data_0_10(store_io_out_wr_0_bits_data_0_10),
    .io_out_wr_0_bits_data_0_11(store_io_out_wr_0_bits_data_0_11),
    .io_out_wr_0_bits_data_0_12(store_io_out_wr_0_bits_data_0_12),
    .io_out_wr_0_bits_data_0_13(store_io_out_wr_0_bits_data_0_13),
    .io_out_wr_0_bits_data_0_14(store_io_out_wr_0_bits_data_0_14),
    .io_out_wr_0_bits_data_0_15(store_io_out_wr_0_bits_data_0_15),
    .io_out_wr_0_bits_data_0_16(store_io_out_wr_0_bits_data_0_16),
    .io_out_wr_0_bits_data_0_17(store_io_out_wr_0_bits_data_0_17),
    .io_out_wr_0_bits_data_0_18(store_io_out_wr_0_bits_data_0_18),
    .io_out_wr_0_bits_data_0_19(store_io_out_wr_0_bits_data_0_19),
    .io_out_wr_0_bits_data_0_20(store_io_out_wr_0_bits_data_0_20),
    .io_out_wr_0_bits_data_0_21(store_io_out_wr_0_bits_data_0_21),
    .io_out_wr_0_bits_data_0_22(store_io_out_wr_0_bits_data_0_22),
    .io_out_wr_0_bits_data_0_23(store_io_out_wr_0_bits_data_0_23),
    .io_out_wr_0_bits_data_0_24(store_io_out_wr_0_bits_data_0_24),
    .io_out_wr_0_bits_data_0_25(store_io_out_wr_0_bits_data_0_25),
    .io_out_wr_0_bits_data_0_26(store_io_out_wr_0_bits_data_0_26),
    .io_out_wr_0_bits_data_0_27(store_io_out_wr_0_bits_data_0_27),
    .io_out_wr_0_bits_data_0_28(store_io_out_wr_0_bits_data_0_28),
    .io_out_wr_0_bits_data_0_29(store_io_out_wr_0_bits_data_0_29),
    .io_out_wr_0_bits_data_0_30(store_io_out_wr_0_bits_data_0_30),
    .io_out_wr_0_bits_data_0_31(store_io_out_wr_0_bits_data_0_31)
  );
  EventCounters ecounters ( // @[Core.scala 71:25]
    .clock(ecounters_clock),
    .reset(ecounters_reset),
    .io_launch(ecounters_io_launch),
    .io_finish(ecounters_io_finish),
    .io_ecnt_0_valid(ecounters_io_ecnt_0_valid),
    .io_ecnt_0_bits(ecounters_io_ecnt_0_bits),
    .io_ucnt_0_valid(ecounters_io_ucnt_0_valid),
    .io_ucnt_0_bits(ecounters_io_ucnt_0_bits),
    .io_acc_wr_event(ecounters_io_acc_wr_event)
  );
  assign io_vcr_finish = finish; // @[Core.scala 120:17]
  assign io_vcr_ecnt_0_valid = ecounters_io_ecnt_0_valid; // @[Core.scala 114:15]
  assign io_vcr_ecnt_0_bits = ecounters_io_ecnt_0_bits; // @[Core.scala 114:15]
  assign io_vcr_ucnt_0_valid = ecounters_io_ucnt_0_valid; // @[Core.scala 115:15]
  assign io_vcr_ucnt_0_bits = ecounters_io_ucnt_0_bits; // @[Core.scala 115:15]
  assign io_vme_rd_0_cmd_valid = fetch_io_vme_rd_cmd_valid; // @[Core.scala 74:16]
  assign io_vme_rd_0_cmd_bits_addr = fetch_io_vme_rd_cmd_bits_addr; // @[Core.scala 74:16]
  assign io_vme_rd_0_cmd_bits_len = fetch_io_vme_rd_cmd_bits_len; // @[Core.scala 74:16]
  assign io_vme_rd_0_data_ready = fetch_io_vme_rd_data_ready; // @[Core.scala 74:16]
  assign io_vme_rd_1_cmd_valid = compute_io_vme_rd_0_cmd_valid; // @[Core.scala 75:16]
  assign io_vme_rd_1_cmd_bits_addr = compute_io_vme_rd_0_cmd_bits_addr; // @[Core.scala 75:16]
  assign io_vme_rd_1_cmd_bits_len = compute_io_vme_rd_0_cmd_bits_len; // @[Core.scala 75:16]
  assign io_vme_rd_1_cmd_bits_tag = compute_io_vme_rd_0_cmd_bits_tag; // @[Core.scala 75:16]
  assign io_vme_rd_2_cmd_valid = load_io_vme_rd_0_cmd_valid; // @[Core.scala 76:16]
  assign io_vme_rd_2_cmd_bits_addr = load_io_vme_rd_0_cmd_bits_addr; // @[Core.scala 76:16]
  assign io_vme_rd_2_cmd_bits_len = load_io_vme_rd_0_cmd_bits_len; // @[Core.scala 76:16]
  assign io_vme_rd_2_cmd_bits_tag = load_io_vme_rd_0_cmd_bits_tag; // @[Core.scala 76:16]
  assign io_vme_rd_3_cmd_valid = load_io_vme_rd_1_cmd_valid; // @[Core.scala 77:16]
  assign io_vme_rd_3_cmd_bits_addr = load_io_vme_rd_1_cmd_bits_addr; // @[Core.scala 77:16]
  assign io_vme_rd_3_cmd_bits_len = load_io_vme_rd_1_cmd_bits_len; // @[Core.scala 77:16]
  assign io_vme_rd_3_cmd_bits_tag = load_io_vme_rd_1_cmd_bits_tag; // @[Core.scala 77:16]
  assign io_vme_rd_4_cmd_valid = compute_io_vme_rd_1_cmd_valid; // @[Core.scala 78:16]
  assign io_vme_rd_4_cmd_bits_addr = compute_io_vme_rd_1_cmd_bits_addr; // @[Core.scala 78:16]
  assign io_vme_rd_4_cmd_bits_len = compute_io_vme_rd_1_cmd_bits_len; // @[Core.scala 78:16]
  assign io_vme_rd_4_cmd_bits_tag = compute_io_vme_rd_1_cmd_bits_tag; // @[Core.scala 78:16]
  assign io_vme_wr_0_cmd_valid = store_io_vme_wr_cmd_valid; // @[Core.scala 79:16]
  assign io_vme_wr_0_cmd_bits_addr = store_io_vme_wr_cmd_bits_addr; // @[Core.scala 79:16]
  assign io_vme_wr_0_cmd_bits_len = store_io_vme_wr_cmd_bits_len; // @[Core.scala 79:16]
  assign io_vme_wr_0_data_valid = store_io_vme_wr_data_valid; // @[Core.scala 79:16]
  assign io_vme_wr_0_data_bits_data = store_io_vme_wr_data_bits_data; // @[Core.scala 79:16]
  assign fetch_clock = clock;
  assign fetch_reset = reset;
  assign fetch_io_launch = io_vcr_launch; // @[Core.scala 82:19]
  assign fetch_io_ins_baddr = io_vcr_ptrs_0; // @[Core.scala 83:22]
  assign fetch_io_ins_count = io_vcr_vals_0; // @[Core.scala 84:22]
  assign fetch_io_vme_rd_cmd_ready = io_vme_rd_0_cmd_ready; // @[Core.scala 74:16]
  assign fetch_io_vme_rd_data_valid = io_vme_rd_0_data_valid; // @[Core.scala 74:16]
  assign fetch_io_vme_rd_data_bits_data = io_vme_rd_0_data_bits_data; // @[Core.scala 74:16]
  assign fetch_io_inst_ld_ready = load_io_inst_ready; // @[Core.scala 88:16]
  assign fetch_io_inst_co_ready = compute_io_inst_ready; // @[Core.scala 97:19]
  assign fetch_io_inst_st_ready = store_io_inst_ready; // @[Core.scala 107:17]
  assign load_clock = clock;
  assign load_reset = reset;
  assign load_io_i_post = compute_io_o_post_0; // @[Core.scala 87:18]
  assign load_io_inst_valid = fetch_io_inst_ld_valid; // @[Core.scala 88:16]
  assign load_io_inst_bits = fetch_io_inst_ld_bits; // @[Core.scala 88:16]
  assign load_io_inp_baddr = io_vcr_ptrs_2; // @[Core.scala 89:21]
  assign load_io_wgt_baddr = io_vcr_ptrs_3; // @[Core.scala 90:21]
  assign load_io_vme_rd_0_cmd_ready = io_vme_rd_2_cmd_ready; // @[Core.scala 76:16]
  assign load_io_vme_rd_0_data_valid = io_vme_rd_2_data_valid; // @[Core.scala 76:16]
  assign load_io_vme_rd_0_data_bits_data = io_vme_rd_2_data_bits_data; // @[Core.scala 76:16]
  assign load_io_vme_rd_0_data_bits_tag = io_vme_rd_2_data_bits_tag; // @[Core.scala 76:16]
  assign load_io_vme_rd_1_cmd_ready = io_vme_rd_3_cmd_ready; // @[Core.scala 77:16]
  assign load_io_vme_rd_1_data_valid = io_vme_rd_3_data_valid; // @[Core.scala 77:16]
  assign load_io_vme_rd_1_data_bits_data = io_vme_rd_3_data_bits_data; // @[Core.scala 77:16]
  assign load_io_vme_rd_1_data_bits_tag = io_vme_rd_3_data_bits_tag; // @[Core.scala 77:16]
  assign load_io_inp_rd_0_idx_valid = compute_io_inp_rd_0_idx_valid; // @[Core.scala 100:18]
  assign load_io_inp_rd_0_idx_bits = compute_io_inp_rd_0_idx_bits; // @[Core.scala 100:18]
  assign load_io_wgt_rd_0_idx_valid = compute_io_wgt_rd_0_idx_valid; // @[Core.scala 101:18]
  assign load_io_wgt_rd_0_idx_bits = compute_io_wgt_rd_0_idx_bits; // @[Core.scala 101:18]
  assign compute_clock = clock;
  assign compute_reset = reset;
  assign compute_io_i_post_0 = load_io_o_post; // @[Core.scala 95:24]
  assign compute_io_i_post_1 = store_io_o_post; // @[Core.scala 96:24]
  assign compute_io_inst_valid = fetch_io_inst_co_valid; // @[Core.scala 97:19]
  assign compute_io_inst_bits = fetch_io_inst_co_bits; // @[Core.scala 97:19]
  assign compute_io_uop_baddr = io_vcr_ptrs_1; // @[Core.scala 98:24]
  assign compute_io_acc_baddr = io_vcr_ptrs_4; // @[Core.scala 99:24]
  assign compute_io_vme_rd_0_cmd_ready = io_vme_rd_1_cmd_ready; // @[Core.scala 75:16]
  assign compute_io_vme_rd_0_data_valid = io_vme_rd_1_data_valid; // @[Core.scala 75:16]
  assign compute_io_vme_rd_0_data_bits_data = io_vme_rd_1_data_bits_data; // @[Core.scala 75:16]
  assign compute_io_vme_rd_0_data_bits_tag = io_vme_rd_1_data_bits_tag; // @[Core.scala 75:16]
  assign compute_io_vme_rd_0_data_bits_last = io_vme_rd_1_data_bits_last; // @[Core.scala 75:16]
  assign compute_io_vme_rd_1_cmd_ready = io_vme_rd_4_cmd_ready; // @[Core.scala 78:16]
  assign compute_io_vme_rd_1_data_valid = io_vme_rd_4_data_valid; // @[Core.scala 78:16]
  assign compute_io_vme_rd_1_data_bits_data = io_vme_rd_4_data_bits_data; // @[Core.scala 78:16]
  assign compute_io_vme_rd_1_data_bits_tag = io_vme_rd_4_data_bits_tag; // @[Core.scala 78:16]
  assign compute_io_inp_rd_0_data_valid = load_io_inp_rd_0_data_valid; // @[Core.scala 100:18]
  assign compute_io_inp_rd_0_data_bits_0_0 = load_io_inp_rd_0_data_bits_0_0; // @[Core.scala 100:18]
  assign compute_io_inp_rd_0_data_bits_0_1 = load_io_inp_rd_0_data_bits_0_1; // @[Core.scala 100:18]
  assign compute_io_inp_rd_0_data_bits_0_2 = load_io_inp_rd_0_data_bits_0_2; // @[Core.scala 100:18]
  assign compute_io_inp_rd_0_data_bits_0_3 = load_io_inp_rd_0_data_bits_0_3; // @[Core.scala 100:18]
  assign compute_io_inp_rd_0_data_bits_0_4 = load_io_inp_rd_0_data_bits_0_4; // @[Core.scala 100:18]
  assign compute_io_inp_rd_0_data_bits_0_5 = load_io_inp_rd_0_data_bits_0_5; // @[Core.scala 100:18]
  assign compute_io_inp_rd_0_data_bits_0_6 = load_io_inp_rd_0_data_bits_0_6; // @[Core.scala 100:18]
  assign compute_io_inp_rd_0_data_bits_0_7 = load_io_inp_rd_0_data_bits_0_7; // @[Core.scala 100:18]
  assign compute_io_inp_rd_0_data_bits_0_8 = load_io_inp_rd_0_data_bits_0_8; // @[Core.scala 100:18]
  assign compute_io_inp_rd_0_data_bits_0_9 = load_io_inp_rd_0_data_bits_0_9; // @[Core.scala 100:18]
  assign compute_io_inp_rd_0_data_bits_0_10 = load_io_inp_rd_0_data_bits_0_10; // @[Core.scala 100:18]
  assign compute_io_inp_rd_0_data_bits_0_11 = load_io_inp_rd_0_data_bits_0_11; // @[Core.scala 100:18]
  assign compute_io_inp_rd_0_data_bits_0_12 = load_io_inp_rd_0_data_bits_0_12; // @[Core.scala 100:18]
  assign compute_io_inp_rd_0_data_bits_0_13 = load_io_inp_rd_0_data_bits_0_13; // @[Core.scala 100:18]
  assign compute_io_inp_rd_0_data_bits_0_14 = load_io_inp_rd_0_data_bits_0_14; // @[Core.scala 100:18]
  assign compute_io_inp_rd_0_data_bits_0_15 = load_io_inp_rd_0_data_bits_0_15; // @[Core.scala 100:18]
  assign compute_io_wgt_rd_0_data_valid = load_io_wgt_rd_0_data_valid; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_0_0 = load_io_wgt_rd_0_data_bits_0_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_0_1 = load_io_wgt_rd_0_data_bits_0_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_0_2 = load_io_wgt_rd_0_data_bits_0_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_0_3 = load_io_wgt_rd_0_data_bits_0_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_0_4 = load_io_wgt_rd_0_data_bits_0_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_0_5 = load_io_wgt_rd_0_data_bits_0_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_0_6 = load_io_wgt_rd_0_data_bits_0_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_0_7 = load_io_wgt_rd_0_data_bits_0_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_0_8 = load_io_wgt_rd_0_data_bits_0_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_0_9 = load_io_wgt_rd_0_data_bits_0_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_0_10 = load_io_wgt_rd_0_data_bits_0_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_0_11 = load_io_wgt_rd_0_data_bits_0_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_0_12 = load_io_wgt_rd_0_data_bits_0_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_0_13 = load_io_wgt_rd_0_data_bits_0_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_0_14 = load_io_wgt_rd_0_data_bits_0_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_0_15 = load_io_wgt_rd_0_data_bits_0_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_1_0 = load_io_wgt_rd_0_data_bits_1_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_1_1 = load_io_wgt_rd_0_data_bits_1_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_1_2 = load_io_wgt_rd_0_data_bits_1_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_1_3 = load_io_wgt_rd_0_data_bits_1_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_1_4 = load_io_wgt_rd_0_data_bits_1_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_1_5 = load_io_wgt_rd_0_data_bits_1_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_1_6 = load_io_wgt_rd_0_data_bits_1_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_1_7 = load_io_wgt_rd_0_data_bits_1_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_1_8 = load_io_wgt_rd_0_data_bits_1_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_1_9 = load_io_wgt_rd_0_data_bits_1_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_1_10 = load_io_wgt_rd_0_data_bits_1_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_1_11 = load_io_wgt_rd_0_data_bits_1_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_1_12 = load_io_wgt_rd_0_data_bits_1_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_1_13 = load_io_wgt_rd_0_data_bits_1_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_1_14 = load_io_wgt_rd_0_data_bits_1_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_1_15 = load_io_wgt_rd_0_data_bits_1_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_2_0 = load_io_wgt_rd_0_data_bits_2_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_2_1 = load_io_wgt_rd_0_data_bits_2_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_2_2 = load_io_wgt_rd_0_data_bits_2_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_2_3 = load_io_wgt_rd_0_data_bits_2_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_2_4 = load_io_wgt_rd_0_data_bits_2_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_2_5 = load_io_wgt_rd_0_data_bits_2_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_2_6 = load_io_wgt_rd_0_data_bits_2_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_2_7 = load_io_wgt_rd_0_data_bits_2_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_2_8 = load_io_wgt_rd_0_data_bits_2_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_2_9 = load_io_wgt_rd_0_data_bits_2_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_2_10 = load_io_wgt_rd_0_data_bits_2_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_2_11 = load_io_wgt_rd_0_data_bits_2_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_2_12 = load_io_wgt_rd_0_data_bits_2_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_2_13 = load_io_wgt_rd_0_data_bits_2_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_2_14 = load_io_wgt_rd_0_data_bits_2_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_2_15 = load_io_wgt_rd_0_data_bits_2_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_3_0 = load_io_wgt_rd_0_data_bits_3_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_3_1 = load_io_wgt_rd_0_data_bits_3_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_3_2 = load_io_wgt_rd_0_data_bits_3_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_3_3 = load_io_wgt_rd_0_data_bits_3_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_3_4 = load_io_wgt_rd_0_data_bits_3_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_3_5 = load_io_wgt_rd_0_data_bits_3_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_3_6 = load_io_wgt_rd_0_data_bits_3_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_3_7 = load_io_wgt_rd_0_data_bits_3_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_3_8 = load_io_wgt_rd_0_data_bits_3_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_3_9 = load_io_wgt_rd_0_data_bits_3_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_3_10 = load_io_wgt_rd_0_data_bits_3_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_3_11 = load_io_wgt_rd_0_data_bits_3_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_3_12 = load_io_wgt_rd_0_data_bits_3_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_3_13 = load_io_wgt_rd_0_data_bits_3_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_3_14 = load_io_wgt_rd_0_data_bits_3_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_3_15 = load_io_wgt_rd_0_data_bits_3_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_4_0 = load_io_wgt_rd_0_data_bits_4_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_4_1 = load_io_wgt_rd_0_data_bits_4_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_4_2 = load_io_wgt_rd_0_data_bits_4_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_4_3 = load_io_wgt_rd_0_data_bits_4_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_4_4 = load_io_wgt_rd_0_data_bits_4_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_4_5 = load_io_wgt_rd_0_data_bits_4_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_4_6 = load_io_wgt_rd_0_data_bits_4_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_4_7 = load_io_wgt_rd_0_data_bits_4_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_4_8 = load_io_wgt_rd_0_data_bits_4_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_4_9 = load_io_wgt_rd_0_data_bits_4_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_4_10 = load_io_wgt_rd_0_data_bits_4_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_4_11 = load_io_wgt_rd_0_data_bits_4_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_4_12 = load_io_wgt_rd_0_data_bits_4_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_4_13 = load_io_wgt_rd_0_data_bits_4_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_4_14 = load_io_wgt_rd_0_data_bits_4_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_4_15 = load_io_wgt_rd_0_data_bits_4_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_5_0 = load_io_wgt_rd_0_data_bits_5_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_5_1 = load_io_wgt_rd_0_data_bits_5_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_5_2 = load_io_wgt_rd_0_data_bits_5_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_5_3 = load_io_wgt_rd_0_data_bits_5_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_5_4 = load_io_wgt_rd_0_data_bits_5_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_5_5 = load_io_wgt_rd_0_data_bits_5_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_5_6 = load_io_wgt_rd_0_data_bits_5_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_5_7 = load_io_wgt_rd_0_data_bits_5_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_5_8 = load_io_wgt_rd_0_data_bits_5_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_5_9 = load_io_wgt_rd_0_data_bits_5_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_5_10 = load_io_wgt_rd_0_data_bits_5_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_5_11 = load_io_wgt_rd_0_data_bits_5_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_5_12 = load_io_wgt_rd_0_data_bits_5_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_5_13 = load_io_wgt_rd_0_data_bits_5_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_5_14 = load_io_wgt_rd_0_data_bits_5_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_5_15 = load_io_wgt_rd_0_data_bits_5_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_6_0 = load_io_wgt_rd_0_data_bits_6_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_6_1 = load_io_wgt_rd_0_data_bits_6_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_6_2 = load_io_wgt_rd_0_data_bits_6_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_6_3 = load_io_wgt_rd_0_data_bits_6_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_6_4 = load_io_wgt_rd_0_data_bits_6_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_6_5 = load_io_wgt_rd_0_data_bits_6_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_6_6 = load_io_wgt_rd_0_data_bits_6_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_6_7 = load_io_wgt_rd_0_data_bits_6_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_6_8 = load_io_wgt_rd_0_data_bits_6_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_6_9 = load_io_wgt_rd_0_data_bits_6_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_6_10 = load_io_wgt_rd_0_data_bits_6_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_6_11 = load_io_wgt_rd_0_data_bits_6_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_6_12 = load_io_wgt_rd_0_data_bits_6_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_6_13 = load_io_wgt_rd_0_data_bits_6_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_6_14 = load_io_wgt_rd_0_data_bits_6_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_6_15 = load_io_wgt_rd_0_data_bits_6_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_7_0 = load_io_wgt_rd_0_data_bits_7_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_7_1 = load_io_wgt_rd_0_data_bits_7_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_7_2 = load_io_wgt_rd_0_data_bits_7_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_7_3 = load_io_wgt_rd_0_data_bits_7_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_7_4 = load_io_wgt_rd_0_data_bits_7_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_7_5 = load_io_wgt_rd_0_data_bits_7_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_7_6 = load_io_wgt_rd_0_data_bits_7_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_7_7 = load_io_wgt_rd_0_data_bits_7_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_7_8 = load_io_wgt_rd_0_data_bits_7_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_7_9 = load_io_wgt_rd_0_data_bits_7_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_7_10 = load_io_wgt_rd_0_data_bits_7_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_7_11 = load_io_wgt_rd_0_data_bits_7_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_7_12 = load_io_wgt_rd_0_data_bits_7_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_7_13 = load_io_wgt_rd_0_data_bits_7_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_7_14 = load_io_wgt_rd_0_data_bits_7_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_7_15 = load_io_wgt_rd_0_data_bits_7_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_8_0 = load_io_wgt_rd_0_data_bits_8_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_8_1 = load_io_wgt_rd_0_data_bits_8_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_8_2 = load_io_wgt_rd_0_data_bits_8_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_8_3 = load_io_wgt_rd_0_data_bits_8_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_8_4 = load_io_wgt_rd_0_data_bits_8_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_8_5 = load_io_wgt_rd_0_data_bits_8_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_8_6 = load_io_wgt_rd_0_data_bits_8_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_8_7 = load_io_wgt_rd_0_data_bits_8_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_8_8 = load_io_wgt_rd_0_data_bits_8_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_8_9 = load_io_wgt_rd_0_data_bits_8_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_8_10 = load_io_wgt_rd_0_data_bits_8_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_8_11 = load_io_wgt_rd_0_data_bits_8_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_8_12 = load_io_wgt_rd_0_data_bits_8_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_8_13 = load_io_wgt_rd_0_data_bits_8_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_8_14 = load_io_wgt_rd_0_data_bits_8_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_8_15 = load_io_wgt_rd_0_data_bits_8_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_9_0 = load_io_wgt_rd_0_data_bits_9_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_9_1 = load_io_wgt_rd_0_data_bits_9_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_9_2 = load_io_wgt_rd_0_data_bits_9_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_9_3 = load_io_wgt_rd_0_data_bits_9_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_9_4 = load_io_wgt_rd_0_data_bits_9_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_9_5 = load_io_wgt_rd_0_data_bits_9_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_9_6 = load_io_wgt_rd_0_data_bits_9_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_9_7 = load_io_wgt_rd_0_data_bits_9_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_9_8 = load_io_wgt_rd_0_data_bits_9_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_9_9 = load_io_wgt_rd_0_data_bits_9_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_9_10 = load_io_wgt_rd_0_data_bits_9_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_9_11 = load_io_wgt_rd_0_data_bits_9_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_9_12 = load_io_wgt_rd_0_data_bits_9_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_9_13 = load_io_wgt_rd_0_data_bits_9_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_9_14 = load_io_wgt_rd_0_data_bits_9_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_9_15 = load_io_wgt_rd_0_data_bits_9_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_10_0 = load_io_wgt_rd_0_data_bits_10_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_10_1 = load_io_wgt_rd_0_data_bits_10_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_10_2 = load_io_wgt_rd_0_data_bits_10_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_10_3 = load_io_wgt_rd_0_data_bits_10_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_10_4 = load_io_wgt_rd_0_data_bits_10_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_10_5 = load_io_wgt_rd_0_data_bits_10_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_10_6 = load_io_wgt_rd_0_data_bits_10_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_10_7 = load_io_wgt_rd_0_data_bits_10_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_10_8 = load_io_wgt_rd_0_data_bits_10_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_10_9 = load_io_wgt_rd_0_data_bits_10_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_10_10 = load_io_wgt_rd_0_data_bits_10_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_10_11 = load_io_wgt_rd_0_data_bits_10_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_10_12 = load_io_wgt_rd_0_data_bits_10_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_10_13 = load_io_wgt_rd_0_data_bits_10_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_10_14 = load_io_wgt_rd_0_data_bits_10_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_10_15 = load_io_wgt_rd_0_data_bits_10_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_11_0 = load_io_wgt_rd_0_data_bits_11_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_11_1 = load_io_wgt_rd_0_data_bits_11_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_11_2 = load_io_wgt_rd_0_data_bits_11_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_11_3 = load_io_wgt_rd_0_data_bits_11_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_11_4 = load_io_wgt_rd_0_data_bits_11_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_11_5 = load_io_wgt_rd_0_data_bits_11_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_11_6 = load_io_wgt_rd_0_data_bits_11_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_11_7 = load_io_wgt_rd_0_data_bits_11_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_11_8 = load_io_wgt_rd_0_data_bits_11_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_11_9 = load_io_wgt_rd_0_data_bits_11_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_11_10 = load_io_wgt_rd_0_data_bits_11_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_11_11 = load_io_wgt_rd_0_data_bits_11_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_11_12 = load_io_wgt_rd_0_data_bits_11_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_11_13 = load_io_wgt_rd_0_data_bits_11_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_11_14 = load_io_wgt_rd_0_data_bits_11_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_11_15 = load_io_wgt_rd_0_data_bits_11_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_12_0 = load_io_wgt_rd_0_data_bits_12_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_12_1 = load_io_wgt_rd_0_data_bits_12_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_12_2 = load_io_wgt_rd_0_data_bits_12_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_12_3 = load_io_wgt_rd_0_data_bits_12_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_12_4 = load_io_wgt_rd_0_data_bits_12_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_12_5 = load_io_wgt_rd_0_data_bits_12_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_12_6 = load_io_wgt_rd_0_data_bits_12_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_12_7 = load_io_wgt_rd_0_data_bits_12_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_12_8 = load_io_wgt_rd_0_data_bits_12_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_12_9 = load_io_wgt_rd_0_data_bits_12_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_12_10 = load_io_wgt_rd_0_data_bits_12_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_12_11 = load_io_wgt_rd_0_data_bits_12_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_12_12 = load_io_wgt_rd_0_data_bits_12_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_12_13 = load_io_wgt_rd_0_data_bits_12_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_12_14 = load_io_wgt_rd_0_data_bits_12_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_12_15 = load_io_wgt_rd_0_data_bits_12_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_13_0 = load_io_wgt_rd_0_data_bits_13_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_13_1 = load_io_wgt_rd_0_data_bits_13_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_13_2 = load_io_wgt_rd_0_data_bits_13_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_13_3 = load_io_wgt_rd_0_data_bits_13_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_13_4 = load_io_wgt_rd_0_data_bits_13_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_13_5 = load_io_wgt_rd_0_data_bits_13_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_13_6 = load_io_wgt_rd_0_data_bits_13_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_13_7 = load_io_wgt_rd_0_data_bits_13_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_13_8 = load_io_wgt_rd_0_data_bits_13_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_13_9 = load_io_wgt_rd_0_data_bits_13_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_13_10 = load_io_wgt_rd_0_data_bits_13_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_13_11 = load_io_wgt_rd_0_data_bits_13_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_13_12 = load_io_wgt_rd_0_data_bits_13_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_13_13 = load_io_wgt_rd_0_data_bits_13_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_13_14 = load_io_wgt_rd_0_data_bits_13_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_13_15 = load_io_wgt_rd_0_data_bits_13_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_14_0 = load_io_wgt_rd_0_data_bits_14_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_14_1 = load_io_wgt_rd_0_data_bits_14_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_14_2 = load_io_wgt_rd_0_data_bits_14_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_14_3 = load_io_wgt_rd_0_data_bits_14_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_14_4 = load_io_wgt_rd_0_data_bits_14_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_14_5 = load_io_wgt_rd_0_data_bits_14_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_14_6 = load_io_wgt_rd_0_data_bits_14_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_14_7 = load_io_wgt_rd_0_data_bits_14_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_14_8 = load_io_wgt_rd_0_data_bits_14_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_14_9 = load_io_wgt_rd_0_data_bits_14_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_14_10 = load_io_wgt_rd_0_data_bits_14_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_14_11 = load_io_wgt_rd_0_data_bits_14_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_14_12 = load_io_wgt_rd_0_data_bits_14_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_14_13 = load_io_wgt_rd_0_data_bits_14_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_14_14 = load_io_wgt_rd_0_data_bits_14_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_14_15 = load_io_wgt_rd_0_data_bits_14_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_15_0 = load_io_wgt_rd_0_data_bits_15_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_15_1 = load_io_wgt_rd_0_data_bits_15_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_15_2 = load_io_wgt_rd_0_data_bits_15_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_15_3 = load_io_wgt_rd_0_data_bits_15_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_15_4 = load_io_wgt_rd_0_data_bits_15_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_15_5 = load_io_wgt_rd_0_data_bits_15_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_15_6 = load_io_wgt_rd_0_data_bits_15_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_15_7 = load_io_wgt_rd_0_data_bits_15_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_15_8 = load_io_wgt_rd_0_data_bits_15_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_15_9 = load_io_wgt_rd_0_data_bits_15_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_15_10 = load_io_wgt_rd_0_data_bits_15_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_15_11 = load_io_wgt_rd_0_data_bits_15_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_15_12 = load_io_wgt_rd_0_data_bits_15_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_15_13 = load_io_wgt_rd_0_data_bits_15_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_15_14 = load_io_wgt_rd_0_data_bits_15_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_15_15 = load_io_wgt_rd_0_data_bits_15_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_16_0 = load_io_wgt_rd_0_data_bits_16_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_16_1 = load_io_wgt_rd_0_data_bits_16_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_16_2 = load_io_wgt_rd_0_data_bits_16_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_16_3 = load_io_wgt_rd_0_data_bits_16_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_16_4 = load_io_wgt_rd_0_data_bits_16_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_16_5 = load_io_wgt_rd_0_data_bits_16_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_16_6 = load_io_wgt_rd_0_data_bits_16_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_16_7 = load_io_wgt_rd_0_data_bits_16_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_16_8 = load_io_wgt_rd_0_data_bits_16_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_16_9 = load_io_wgt_rd_0_data_bits_16_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_16_10 = load_io_wgt_rd_0_data_bits_16_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_16_11 = load_io_wgt_rd_0_data_bits_16_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_16_12 = load_io_wgt_rd_0_data_bits_16_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_16_13 = load_io_wgt_rd_0_data_bits_16_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_16_14 = load_io_wgt_rd_0_data_bits_16_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_16_15 = load_io_wgt_rd_0_data_bits_16_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_17_0 = load_io_wgt_rd_0_data_bits_17_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_17_1 = load_io_wgt_rd_0_data_bits_17_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_17_2 = load_io_wgt_rd_0_data_bits_17_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_17_3 = load_io_wgt_rd_0_data_bits_17_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_17_4 = load_io_wgt_rd_0_data_bits_17_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_17_5 = load_io_wgt_rd_0_data_bits_17_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_17_6 = load_io_wgt_rd_0_data_bits_17_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_17_7 = load_io_wgt_rd_0_data_bits_17_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_17_8 = load_io_wgt_rd_0_data_bits_17_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_17_9 = load_io_wgt_rd_0_data_bits_17_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_17_10 = load_io_wgt_rd_0_data_bits_17_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_17_11 = load_io_wgt_rd_0_data_bits_17_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_17_12 = load_io_wgt_rd_0_data_bits_17_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_17_13 = load_io_wgt_rd_0_data_bits_17_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_17_14 = load_io_wgt_rd_0_data_bits_17_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_17_15 = load_io_wgt_rd_0_data_bits_17_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_18_0 = load_io_wgt_rd_0_data_bits_18_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_18_1 = load_io_wgt_rd_0_data_bits_18_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_18_2 = load_io_wgt_rd_0_data_bits_18_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_18_3 = load_io_wgt_rd_0_data_bits_18_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_18_4 = load_io_wgt_rd_0_data_bits_18_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_18_5 = load_io_wgt_rd_0_data_bits_18_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_18_6 = load_io_wgt_rd_0_data_bits_18_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_18_7 = load_io_wgt_rd_0_data_bits_18_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_18_8 = load_io_wgt_rd_0_data_bits_18_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_18_9 = load_io_wgt_rd_0_data_bits_18_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_18_10 = load_io_wgt_rd_0_data_bits_18_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_18_11 = load_io_wgt_rd_0_data_bits_18_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_18_12 = load_io_wgt_rd_0_data_bits_18_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_18_13 = load_io_wgt_rd_0_data_bits_18_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_18_14 = load_io_wgt_rd_0_data_bits_18_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_18_15 = load_io_wgt_rd_0_data_bits_18_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_19_0 = load_io_wgt_rd_0_data_bits_19_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_19_1 = load_io_wgt_rd_0_data_bits_19_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_19_2 = load_io_wgt_rd_0_data_bits_19_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_19_3 = load_io_wgt_rd_0_data_bits_19_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_19_4 = load_io_wgt_rd_0_data_bits_19_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_19_5 = load_io_wgt_rd_0_data_bits_19_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_19_6 = load_io_wgt_rd_0_data_bits_19_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_19_7 = load_io_wgt_rd_0_data_bits_19_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_19_8 = load_io_wgt_rd_0_data_bits_19_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_19_9 = load_io_wgt_rd_0_data_bits_19_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_19_10 = load_io_wgt_rd_0_data_bits_19_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_19_11 = load_io_wgt_rd_0_data_bits_19_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_19_12 = load_io_wgt_rd_0_data_bits_19_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_19_13 = load_io_wgt_rd_0_data_bits_19_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_19_14 = load_io_wgt_rd_0_data_bits_19_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_19_15 = load_io_wgt_rd_0_data_bits_19_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_20_0 = load_io_wgt_rd_0_data_bits_20_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_20_1 = load_io_wgt_rd_0_data_bits_20_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_20_2 = load_io_wgt_rd_0_data_bits_20_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_20_3 = load_io_wgt_rd_0_data_bits_20_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_20_4 = load_io_wgt_rd_0_data_bits_20_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_20_5 = load_io_wgt_rd_0_data_bits_20_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_20_6 = load_io_wgt_rd_0_data_bits_20_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_20_7 = load_io_wgt_rd_0_data_bits_20_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_20_8 = load_io_wgt_rd_0_data_bits_20_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_20_9 = load_io_wgt_rd_0_data_bits_20_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_20_10 = load_io_wgt_rd_0_data_bits_20_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_20_11 = load_io_wgt_rd_0_data_bits_20_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_20_12 = load_io_wgt_rd_0_data_bits_20_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_20_13 = load_io_wgt_rd_0_data_bits_20_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_20_14 = load_io_wgt_rd_0_data_bits_20_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_20_15 = load_io_wgt_rd_0_data_bits_20_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_21_0 = load_io_wgt_rd_0_data_bits_21_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_21_1 = load_io_wgt_rd_0_data_bits_21_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_21_2 = load_io_wgt_rd_0_data_bits_21_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_21_3 = load_io_wgt_rd_0_data_bits_21_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_21_4 = load_io_wgt_rd_0_data_bits_21_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_21_5 = load_io_wgt_rd_0_data_bits_21_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_21_6 = load_io_wgt_rd_0_data_bits_21_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_21_7 = load_io_wgt_rd_0_data_bits_21_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_21_8 = load_io_wgt_rd_0_data_bits_21_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_21_9 = load_io_wgt_rd_0_data_bits_21_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_21_10 = load_io_wgt_rd_0_data_bits_21_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_21_11 = load_io_wgt_rd_0_data_bits_21_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_21_12 = load_io_wgt_rd_0_data_bits_21_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_21_13 = load_io_wgt_rd_0_data_bits_21_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_21_14 = load_io_wgt_rd_0_data_bits_21_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_21_15 = load_io_wgt_rd_0_data_bits_21_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_22_0 = load_io_wgt_rd_0_data_bits_22_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_22_1 = load_io_wgt_rd_0_data_bits_22_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_22_2 = load_io_wgt_rd_0_data_bits_22_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_22_3 = load_io_wgt_rd_0_data_bits_22_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_22_4 = load_io_wgt_rd_0_data_bits_22_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_22_5 = load_io_wgt_rd_0_data_bits_22_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_22_6 = load_io_wgt_rd_0_data_bits_22_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_22_7 = load_io_wgt_rd_0_data_bits_22_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_22_8 = load_io_wgt_rd_0_data_bits_22_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_22_9 = load_io_wgt_rd_0_data_bits_22_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_22_10 = load_io_wgt_rd_0_data_bits_22_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_22_11 = load_io_wgt_rd_0_data_bits_22_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_22_12 = load_io_wgt_rd_0_data_bits_22_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_22_13 = load_io_wgt_rd_0_data_bits_22_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_22_14 = load_io_wgt_rd_0_data_bits_22_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_22_15 = load_io_wgt_rd_0_data_bits_22_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_23_0 = load_io_wgt_rd_0_data_bits_23_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_23_1 = load_io_wgt_rd_0_data_bits_23_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_23_2 = load_io_wgt_rd_0_data_bits_23_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_23_3 = load_io_wgt_rd_0_data_bits_23_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_23_4 = load_io_wgt_rd_0_data_bits_23_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_23_5 = load_io_wgt_rd_0_data_bits_23_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_23_6 = load_io_wgt_rd_0_data_bits_23_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_23_7 = load_io_wgt_rd_0_data_bits_23_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_23_8 = load_io_wgt_rd_0_data_bits_23_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_23_9 = load_io_wgt_rd_0_data_bits_23_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_23_10 = load_io_wgt_rd_0_data_bits_23_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_23_11 = load_io_wgt_rd_0_data_bits_23_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_23_12 = load_io_wgt_rd_0_data_bits_23_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_23_13 = load_io_wgt_rd_0_data_bits_23_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_23_14 = load_io_wgt_rd_0_data_bits_23_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_23_15 = load_io_wgt_rd_0_data_bits_23_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_24_0 = load_io_wgt_rd_0_data_bits_24_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_24_1 = load_io_wgt_rd_0_data_bits_24_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_24_2 = load_io_wgt_rd_0_data_bits_24_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_24_3 = load_io_wgt_rd_0_data_bits_24_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_24_4 = load_io_wgt_rd_0_data_bits_24_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_24_5 = load_io_wgt_rd_0_data_bits_24_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_24_6 = load_io_wgt_rd_0_data_bits_24_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_24_7 = load_io_wgt_rd_0_data_bits_24_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_24_8 = load_io_wgt_rd_0_data_bits_24_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_24_9 = load_io_wgt_rd_0_data_bits_24_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_24_10 = load_io_wgt_rd_0_data_bits_24_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_24_11 = load_io_wgt_rd_0_data_bits_24_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_24_12 = load_io_wgt_rd_0_data_bits_24_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_24_13 = load_io_wgt_rd_0_data_bits_24_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_24_14 = load_io_wgt_rd_0_data_bits_24_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_24_15 = load_io_wgt_rd_0_data_bits_24_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_25_0 = load_io_wgt_rd_0_data_bits_25_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_25_1 = load_io_wgt_rd_0_data_bits_25_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_25_2 = load_io_wgt_rd_0_data_bits_25_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_25_3 = load_io_wgt_rd_0_data_bits_25_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_25_4 = load_io_wgt_rd_0_data_bits_25_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_25_5 = load_io_wgt_rd_0_data_bits_25_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_25_6 = load_io_wgt_rd_0_data_bits_25_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_25_7 = load_io_wgt_rd_0_data_bits_25_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_25_8 = load_io_wgt_rd_0_data_bits_25_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_25_9 = load_io_wgt_rd_0_data_bits_25_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_25_10 = load_io_wgt_rd_0_data_bits_25_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_25_11 = load_io_wgt_rd_0_data_bits_25_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_25_12 = load_io_wgt_rd_0_data_bits_25_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_25_13 = load_io_wgt_rd_0_data_bits_25_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_25_14 = load_io_wgt_rd_0_data_bits_25_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_25_15 = load_io_wgt_rd_0_data_bits_25_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_26_0 = load_io_wgt_rd_0_data_bits_26_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_26_1 = load_io_wgt_rd_0_data_bits_26_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_26_2 = load_io_wgt_rd_0_data_bits_26_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_26_3 = load_io_wgt_rd_0_data_bits_26_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_26_4 = load_io_wgt_rd_0_data_bits_26_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_26_5 = load_io_wgt_rd_0_data_bits_26_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_26_6 = load_io_wgt_rd_0_data_bits_26_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_26_7 = load_io_wgt_rd_0_data_bits_26_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_26_8 = load_io_wgt_rd_0_data_bits_26_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_26_9 = load_io_wgt_rd_0_data_bits_26_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_26_10 = load_io_wgt_rd_0_data_bits_26_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_26_11 = load_io_wgt_rd_0_data_bits_26_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_26_12 = load_io_wgt_rd_0_data_bits_26_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_26_13 = load_io_wgt_rd_0_data_bits_26_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_26_14 = load_io_wgt_rd_0_data_bits_26_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_26_15 = load_io_wgt_rd_0_data_bits_26_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_27_0 = load_io_wgt_rd_0_data_bits_27_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_27_1 = load_io_wgt_rd_0_data_bits_27_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_27_2 = load_io_wgt_rd_0_data_bits_27_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_27_3 = load_io_wgt_rd_0_data_bits_27_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_27_4 = load_io_wgt_rd_0_data_bits_27_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_27_5 = load_io_wgt_rd_0_data_bits_27_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_27_6 = load_io_wgt_rd_0_data_bits_27_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_27_7 = load_io_wgt_rd_0_data_bits_27_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_27_8 = load_io_wgt_rd_0_data_bits_27_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_27_9 = load_io_wgt_rd_0_data_bits_27_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_27_10 = load_io_wgt_rd_0_data_bits_27_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_27_11 = load_io_wgt_rd_0_data_bits_27_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_27_12 = load_io_wgt_rd_0_data_bits_27_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_27_13 = load_io_wgt_rd_0_data_bits_27_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_27_14 = load_io_wgt_rd_0_data_bits_27_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_27_15 = load_io_wgt_rd_0_data_bits_27_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_28_0 = load_io_wgt_rd_0_data_bits_28_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_28_1 = load_io_wgt_rd_0_data_bits_28_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_28_2 = load_io_wgt_rd_0_data_bits_28_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_28_3 = load_io_wgt_rd_0_data_bits_28_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_28_4 = load_io_wgt_rd_0_data_bits_28_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_28_5 = load_io_wgt_rd_0_data_bits_28_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_28_6 = load_io_wgt_rd_0_data_bits_28_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_28_7 = load_io_wgt_rd_0_data_bits_28_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_28_8 = load_io_wgt_rd_0_data_bits_28_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_28_9 = load_io_wgt_rd_0_data_bits_28_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_28_10 = load_io_wgt_rd_0_data_bits_28_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_28_11 = load_io_wgt_rd_0_data_bits_28_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_28_12 = load_io_wgt_rd_0_data_bits_28_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_28_13 = load_io_wgt_rd_0_data_bits_28_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_28_14 = load_io_wgt_rd_0_data_bits_28_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_28_15 = load_io_wgt_rd_0_data_bits_28_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_29_0 = load_io_wgt_rd_0_data_bits_29_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_29_1 = load_io_wgt_rd_0_data_bits_29_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_29_2 = load_io_wgt_rd_0_data_bits_29_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_29_3 = load_io_wgt_rd_0_data_bits_29_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_29_4 = load_io_wgt_rd_0_data_bits_29_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_29_5 = load_io_wgt_rd_0_data_bits_29_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_29_6 = load_io_wgt_rd_0_data_bits_29_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_29_7 = load_io_wgt_rd_0_data_bits_29_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_29_8 = load_io_wgt_rd_0_data_bits_29_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_29_9 = load_io_wgt_rd_0_data_bits_29_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_29_10 = load_io_wgt_rd_0_data_bits_29_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_29_11 = load_io_wgt_rd_0_data_bits_29_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_29_12 = load_io_wgt_rd_0_data_bits_29_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_29_13 = load_io_wgt_rd_0_data_bits_29_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_29_14 = load_io_wgt_rd_0_data_bits_29_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_29_15 = load_io_wgt_rd_0_data_bits_29_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_30_0 = load_io_wgt_rd_0_data_bits_30_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_30_1 = load_io_wgt_rd_0_data_bits_30_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_30_2 = load_io_wgt_rd_0_data_bits_30_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_30_3 = load_io_wgt_rd_0_data_bits_30_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_30_4 = load_io_wgt_rd_0_data_bits_30_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_30_5 = load_io_wgt_rd_0_data_bits_30_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_30_6 = load_io_wgt_rd_0_data_bits_30_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_30_7 = load_io_wgt_rd_0_data_bits_30_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_30_8 = load_io_wgt_rd_0_data_bits_30_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_30_9 = load_io_wgt_rd_0_data_bits_30_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_30_10 = load_io_wgt_rd_0_data_bits_30_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_30_11 = load_io_wgt_rd_0_data_bits_30_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_30_12 = load_io_wgt_rd_0_data_bits_30_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_30_13 = load_io_wgt_rd_0_data_bits_30_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_30_14 = load_io_wgt_rd_0_data_bits_30_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_30_15 = load_io_wgt_rd_0_data_bits_30_15; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_31_0 = load_io_wgt_rd_0_data_bits_31_0; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_31_1 = load_io_wgt_rd_0_data_bits_31_1; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_31_2 = load_io_wgt_rd_0_data_bits_31_2; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_31_3 = load_io_wgt_rd_0_data_bits_31_3; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_31_4 = load_io_wgt_rd_0_data_bits_31_4; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_31_5 = load_io_wgt_rd_0_data_bits_31_5; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_31_6 = load_io_wgt_rd_0_data_bits_31_6; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_31_7 = load_io_wgt_rd_0_data_bits_31_7; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_31_8 = load_io_wgt_rd_0_data_bits_31_8; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_31_9 = load_io_wgt_rd_0_data_bits_31_9; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_31_10 = load_io_wgt_rd_0_data_bits_31_10; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_31_11 = load_io_wgt_rd_0_data_bits_31_11; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_31_12 = load_io_wgt_rd_0_data_bits_31_12; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_31_13 = load_io_wgt_rd_0_data_bits_31_13; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_31_14 = load_io_wgt_rd_0_data_bits_31_14; // @[Core.scala 101:18]
  assign compute_io_wgt_rd_0_data_bits_31_15 = load_io_wgt_rd_0_data_bits_31_15; // @[Core.scala 101:18]
  assign store_clock = clock;
  assign store_reset = reset;
  assign store_io_i_post = compute_io_o_post_1; // @[Core.scala 106:19]
  assign store_io_inst_valid = fetch_io_inst_st_valid; // @[Core.scala 107:17]
  assign store_io_inst_bits = fetch_io_inst_st_bits; // @[Core.scala 107:17]
  assign store_io_out_baddr = io_vcr_ptrs_5; // @[Core.scala 108:22]
  assign store_io_vme_wr_cmd_ready = io_vme_wr_0_cmd_ready; // @[Core.scala 79:16]
  assign store_io_vme_wr_data_ready = io_vme_wr_0_data_ready; // @[Core.scala 79:16]
  assign store_io_vme_wr_ack = io_vme_wr_0_ack; // @[Core.scala 79:16]
  assign store_io_out_wr_0_valid = compute_io_out_wr_0_valid; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_idx = compute_io_out_wr_0_bits_idx; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_0 = compute_io_out_wr_0_bits_data_0_0; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_1 = compute_io_out_wr_0_bits_data_0_1; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_2 = compute_io_out_wr_0_bits_data_0_2; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_3 = compute_io_out_wr_0_bits_data_0_3; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_4 = compute_io_out_wr_0_bits_data_0_4; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_5 = compute_io_out_wr_0_bits_data_0_5; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_6 = compute_io_out_wr_0_bits_data_0_6; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_7 = compute_io_out_wr_0_bits_data_0_7; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_8 = compute_io_out_wr_0_bits_data_0_8; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_9 = compute_io_out_wr_0_bits_data_0_9; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_10 = compute_io_out_wr_0_bits_data_0_10; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_11 = compute_io_out_wr_0_bits_data_0_11; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_12 = compute_io_out_wr_0_bits_data_0_12; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_13 = compute_io_out_wr_0_bits_data_0_13; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_14 = compute_io_out_wr_0_bits_data_0_14; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_15 = compute_io_out_wr_0_bits_data_0_15; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_16 = compute_io_out_wr_0_bits_data_0_16; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_17 = compute_io_out_wr_0_bits_data_0_17; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_18 = compute_io_out_wr_0_bits_data_0_18; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_19 = compute_io_out_wr_0_bits_data_0_19; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_20 = compute_io_out_wr_0_bits_data_0_20; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_21 = compute_io_out_wr_0_bits_data_0_21; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_22 = compute_io_out_wr_0_bits_data_0_22; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_23 = compute_io_out_wr_0_bits_data_0_23; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_24 = compute_io_out_wr_0_bits_data_0_24; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_25 = compute_io_out_wr_0_bits_data_0_25; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_26 = compute_io_out_wr_0_bits_data_0_26; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_27 = compute_io_out_wr_0_bits_data_0_27; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_28 = compute_io_out_wr_0_bits_data_0_28; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_29 = compute_io_out_wr_0_bits_data_0_29; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_30 = compute_io_out_wr_0_bits_data_0_30; // @[Core.scala 109:16]
  assign store_io_out_wr_0_bits_data_0_31 = compute_io_out_wr_0_bits_data_0_31; // @[Core.scala 109:16]
  assign ecounters_clock = clock;
  assign ecounters_reset = reset;
  assign ecounters_io_launch = io_vcr_launch; // @[Core.scala 112:23]
  assign ecounters_io_finish = compute_io_finish; // @[Core.scala 113:23]
  assign ecounters_io_acc_wr_event = compute_io_acc_wr_event; // @[Core.scala 116:29]
  always @(posedge clock) begin
    finish <= compute_io_finish; // @[Core.scala 119:23]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  finish = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module IntelShell(
  input         clock,
  input         reset,
  output        io_host_aw_ready,
  input         io_host_aw_valid,
  input  [15:0] io_host_aw_bits_addr,
  input  [12:0] io_host_aw_bits_id,
  input         io_host_aw_bits_user,
  input  [3:0]  io_host_aw_bits_len,
  input  [2:0]  io_host_aw_bits_size,
  input  [1:0]  io_host_aw_bits_burst,
  input  [1:0]  io_host_aw_bits_lock,
  input  [3:0]  io_host_aw_bits_cache,
  input  [2:0]  io_host_aw_bits_prot,
  input  [3:0]  io_host_aw_bits_qos,
  input  [3:0]  io_host_aw_bits_region,
  output        io_host_w_ready,
  input         io_host_w_valid,
  input  [31:0] io_host_w_bits_data,
  input  [3:0]  io_host_w_bits_strb,
  input         io_host_w_bits_last,
  input  [12:0] io_host_w_bits_id,
  input         io_host_w_bits_user,
  input         io_host_b_ready,
  output        io_host_b_valid,
  output [1:0]  io_host_b_bits_resp,
  output [12:0] io_host_b_bits_id,
  output        io_host_b_bits_user,
  output        io_host_ar_ready,
  input         io_host_ar_valid,
  input  [15:0] io_host_ar_bits_addr,
  input  [12:0] io_host_ar_bits_id,
  input         io_host_ar_bits_user,
  input  [3:0]  io_host_ar_bits_len,
  input  [2:0]  io_host_ar_bits_size,
  input  [1:0]  io_host_ar_bits_burst,
  input  [1:0]  io_host_ar_bits_lock,
  input  [3:0]  io_host_ar_bits_cache,
  input  [2:0]  io_host_ar_bits_prot,
  input  [3:0]  io_host_ar_bits_qos,
  input  [3:0]  io_host_ar_bits_region,
  input         io_host_r_ready,
  output        io_host_r_valid,
  output [31:0] io_host_r_bits_data,
  output [1:0]  io_host_r_bits_resp,
  output        io_host_r_bits_last,
  output [12:0] io_host_r_bits_id,
  output        io_host_r_bits_user,
  input         io_mem_aw_ready,
  output        io_mem_aw_valid,
  output [31:0] io_mem_aw_bits_addr,
  output [7:0]  io_mem_aw_bits_id,
  output [4:0]  io_mem_aw_bits_user,
  output [3:0]  io_mem_aw_bits_len,
  output [2:0]  io_mem_aw_bits_size,
  output [1:0]  io_mem_aw_bits_burst,
  output [1:0]  io_mem_aw_bits_lock,
  output [3:0]  io_mem_aw_bits_cache,
  output [2:0]  io_mem_aw_bits_prot,
  output [3:0]  io_mem_aw_bits_qos,
  output [3:0]  io_mem_aw_bits_region,
  input         io_mem_w_ready,
  output        io_mem_w_valid,
  output [63:0] io_mem_w_bits_data,
  output [7:0]  io_mem_w_bits_strb,
  output        io_mem_w_bits_last,
  output [7:0]  io_mem_w_bits_id,
  output [4:0]  io_mem_w_bits_user,
  output        io_mem_b_ready,
  input         io_mem_b_valid,
  input  [1:0]  io_mem_b_bits_resp,
  input  [7:0]  io_mem_b_bits_id,
  input  [4:0]  io_mem_b_bits_user,
  input         io_mem_ar_ready,
  output        io_mem_ar_valid,
  output [31:0] io_mem_ar_bits_addr,
  output [7:0]  io_mem_ar_bits_id,
  output [4:0]  io_mem_ar_bits_user,
  output [3:0]  io_mem_ar_bits_len,
  output [2:0]  io_mem_ar_bits_size,
  output [1:0]  io_mem_ar_bits_burst,
  output [1:0]  io_mem_ar_bits_lock,
  output [3:0]  io_mem_ar_bits_cache,
  output [2:0]  io_mem_ar_bits_prot,
  output [3:0]  io_mem_ar_bits_qos,
  output [3:0]  io_mem_ar_bits_region,
  output        io_mem_r_ready,
  input         io_mem_r_valid,
  input  [63:0] io_mem_r_bits_data,
  input  [1:0]  io_mem_r_bits_resp,
  input         io_mem_r_bits_last,
  input  [7:0]  io_mem_r_bits_id,
  input  [4:0]  io_mem_r_bits_user
);
  wire  vcr_clock; // @[IntelShell.scala 38:19]
  wire  vcr_reset; // @[IntelShell.scala 38:19]
  wire  vcr_io_host_aw_ready; // @[IntelShell.scala 38:19]
  wire  vcr_io_host_aw_valid; // @[IntelShell.scala 38:19]
  wire [15:0] vcr_io_host_aw_bits_addr; // @[IntelShell.scala 38:19]
  wire  vcr_io_host_w_ready; // @[IntelShell.scala 38:19]
  wire  vcr_io_host_w_valid; // @[IntelShell.scala 38:19]
  wire [31:0] vcr_io_host_w_bits_data; // @[IntelShell.scala 38:19]
  wire  vcr_io_host_b_ready; // @[IntelShell.scala 38:19]
  wire  vcr_io_host_b_valid; // @[IntelShell.scala 38:19]
  wire  vcr_io_host_ar_ready; // @[IntelShell.scala 38:19]
  wire  vcr_io_host_ar_valid; // @[IntelShell.scala 38:19]
  wire [15:0] vcr_io_host_ar_bits_addr; // @[IntelShell.scala 38:19]
  wire  vcr_io_host_r_ready; // @[IntelShell.scala 38:19]
  wire  vcr_io_host_r_valid; // @[IntelShell.scala 38:19]
  wire [31:0] vcr_io_host_r_bits_data; // @[IntelShell.scala 38:19]
  wire  vcr_io_vcr_launch; // @[IntelShell.scala 38:19]
  wire  vcr_io_vcr_finish; // @[IntelShell.scala 38:19]
  wire  vcr_io_vcr_ecnt_0_valid; // @[IntelShell.scala 38:19]
  wire [31:0] vcr_io_vcr_ecnt_0_bits; // @[IntelShell.scala 38:19]
  wire [31:0] vcr_io_vcr_vals_0; // @[IntelShell.scala 38:19]
  wire [31:0] vcr_io_vcr_ptrs_0; // @[IntelShell.scala 38:19]
  wire [31:0] vcr_io_vcr_ptrs_1; // @[IntelShell.scala 38:19]
  wire [31:0] vcr_io_vcr_ptrs_2; // @[IntelShell.scala 38:19]
  wire [31:0] vcr_io_vcr_ptrs_3; // @[IntelShell.scala 38:19]
  wire [31:0] vcr_io_vcr_ptrs_4; // @[IntelShell.scala 38:19]
  wire [31:0] vcr_io_vcr_ptrs_5; // @[IntelShell.scala 38:19]
  wire  vcr_io_vcr_ucnt_0_valid; // @[IntelShell.scala 38:19]
  wire [31:0] vcr_io_vcr_ucnt_0_bits; // @[IntelShell.scala 38:19]
  wire  vme_clock; // @[IntelShell.scala 39:19]
  wire  vme_reset; // @[IntelShell.scala 39:19]
  wire  vme_io_mem_aw_ready; // @[IntelShell.scala 39:19]
  wire  vme_io_mem_aw_valid; // @[IntelShell.scala 39:19]
  wire [31:0] vme_io_mem_aw_bits_addr; // @[IntelShell.scala 39:19]
  wire [3:0] vme_io_mem_aw_bits_len; // @[IntelShell.scala 39:19]
  wire  vme_io_mem_w_ready; // @[IntelShell.scala 39:19]
  wire  vme_io_mem_w_valid; // @[IntelShell.scala 39:19]
  wire [63:0] vme_io_mem_w_bits_data; // @[IntelShell.scala 39:19]
  wire  vme_io_mem_w_bits_last; // @[IntelShell.scala 39:19]
  wire  vme_io_mem_b_ready; // @[IntelShell.scala 39:19]
  wire  vme_io_mem_b_valid; // @[IntelShell.scala 39:19]
  wire  vme_io_mem_ar_ready; // @[IntelShell.scala 39:19]
  wire  vme_io_mem_ar_valid; // @[IntelShell.scala 39:19]
  wire [31:0] vme_io_mem_ar_bits_addr; // @[IntelShell.scala 39:19]
  wire [7:0] vme_io_mem_ar_bits_id; // @[IntelShell.scala 39:19]
  wire [3:0] vme_io_mem_ar_bits_len; // @[IntelShell.scala 39:19]
  wire  vme_io_mem_r_valid; // @[IntelShell.scala 39:19]
  wire [63:0] vme_io_mem_r_bits_data; // @[IntelShell.scala 39:19]
  wire  vme_io_mem_r_bits_last; // @[IntelShell.scala 39:19]
  wire [7:0] vme_io_mem_r_bits_id; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_0_cmd_ready; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_0_cmd_valid; // @[IntelShell.scala 39:19]
  wire [31:0] vme_io_vme_rd_0_cmd_bits_addr; // @[IntelShell.scala 39:19]
  wire [3:0] vme_io_vme_rd_0_cmd_bits_len; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_0_data_ready; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_0_data_valid; // @[IntelShell.scala 39:19]
  wire [63:0] vme_io_vme_rd_0_data_bits_data; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_1_cmd_ready; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_1_cmd_valid; // @[IntelShell.scala 39:19]
  wire [31:0] vme_io_vme_rd_1_cmd_bits_addr; // @[IntelShell.scala 39:19]
  wire [3:0] vme_io_vme_rd_1_cmd_bits_len; // @[IntelShell.scala 39:19]
  wire [20:0] vme_io_vme_rd_1_cmd_bits_tag; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_1_data_valid; // @[IntelShell.scala 39:19]
  wire [63:0] vme_io_vme_rd_1_data_bits_data; // @[IntelShell.scala 39:19]
  wire [20:0] vme_io_vme_rd_1_data_bits_tag; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_1_data_bits_last; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_2_cmd_ready; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_2_cmd_valid; // @[IntelShell.scala 39:19]
  wire [31:0] vme_io_vme_rd_2_cmd_bits_addr; // @[IntelShell.scala 39:19]
  wire [3:0] vme_io_vme_rd_2_cmd_bits_len; // @[IntelShell.scala 39:19]
  wire [20:0] vme_io_vme_rd_2_cmd_bits_tag; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_2_data_valid; // @[IntelShell.scala 39:19]
  wire [63:0] vme_io_vme_rd_2_data_bits_data; // @[IntelShell.scala 39:19]
  wire [20:0] vme_io_vme_rd_2_data_bits_tag; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_3_cmd_ready; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_3_cmd_valid; // @[IntelShell.scala 39:19]
  wire [31:0] vme_io_vme_rd_3_cmd_bits_addr; // @[IntelShell.scala 39:19]
  wire [3:0] vme_io_vme_rd_3_cmd_bits_len; // @[IntelShell.scala 39:19]
  wire [20:0] vme_io_vme_rd_3_cmd_bits_tag; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_3_data_valid; // @[IntelShell.scala 39:19]
  wire [63:0] vme_io_vme_rd_3_data_bits_data; // @[IntelShell.scala 39:19]
  wire [20:0] vme_io_vme_rd_3_data_bits_tag; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_4_cmd_ready; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_4_cmd_valid; // @[IntelShell.scala 39:19]
  wire [31:0] vme_io_vme_rd_4_cmd_bits_addr; // @[IntelShell.scala 39:19]
  wire [3:0] vme_io_vme_rd_4_cmd_bits_len; // @[IntelShell.scala 39:19]
  wire [20:0] vme_io_vme_rd_4_cmd_bits_tag; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_rd_4_data_valid; // @[IntelShell.scala 39:19]
  wire [63:0] vme_io_vme_rd_4_data_bits_data; // @[IntelShell.scala 39:19]
  wire [20:0] vme_io_vme_rd_4_data_bits_tag; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_wr_0_cmd_ready; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_wr_0_cmd_valid; // @[IntelShell.scala 39:19]
  wire [31:0] vme_io_vme_wr_0_cmd_bits_addr; // @[IntelShell.scala 39:19]
  wire [3:0] vme_io_vme_wr_0_cmd_bits_len; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_wr_0_data_ready; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_wr_0_data_valid; // @[IntelShell.scala 39:19]
  wire [63:0] vme_io_vme_wr_0_data_bits_data; // @[IntelShell.scala 39:19]
  wire  vme_io_vme_wr_0_ack; // @[IntelShell.scala 39:19]
  wire  core_clock; // @[IntelShell.scala 40:20]
  wire  core_reset; // @[IntelShell.scala 40:20]
  wire  core_io_vcr_launch; // @[IntelShell.scala 40:20]
  wire  core_io_vcr_finish; // @[IntelShell.scala 40:20]
  wire  core_io_vcr_ecnt_0_valid; // @[IntelShell.scala 40:20]
  wire [31:0] core_io_vcr_ecnt_0_bits; // @[IntelShell.scala 40:20]
  wire [31:0] core_io_vcr_vals_0; // @[IntelShell.scala 40:20]
  wire [31:0] core_io_vcr_ptrs_0; // @[IntelShell.scala 40:20]
  wire [31:0] core_io_vcr_ptrs_1; // @[IntelShell.scala 40:20]
  wire [31:0] core_io_vcr_ptrs_2; // @[IntelShell.scala 40:20]
  wire [31:0] core_io_vcr_ptrs_3; // @[IntelShell.scala 40:20]
  wire [31:0] core_io_vcr_ptrs_4; // @[IntelShell.scala 40:20]
  wire [31:0] core_io_vcr_ptrs_5; // @[IntelShell.scala 40:20]
  wire  core_io_vcr_ucnt_0_valid; // @[IntelShell.scala 40:20]
  wire [31:0] core_io_vcr_ucnt_0_bits; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_0_cmd_ready; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_0_cmd_valid; // @[IntelShell.scala 40:20]
  wire [31:0] core_io_vme_rd_0_cmd_bits_addr; // @[IntelShell.scala 40:20]
  wire [3:0] core_io_vme_rd_0_cmd_bits_len; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_0_data_ready; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_0_data_valid; // @[IntelShell.scala 40:20]
  wire [63:0] core_io_vme_rd_0_data_bits_data; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_1_cmd_ready; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_1_cmd_valid; // @[IntelShell.scala 40:20]
  wire [31:0] core_io_vme_rd_1_cmd_bits_addr; // @[IntelShell.scala 40:20]
  wire [3:0] core_io_vme_rd_1_cmd_bits_len; // @[IntelShell.scala 40:20]
  wire [20:0] core_io_vme_rd_1_cmd_bits_tag; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_1_data_valid; // @[IntelShell.scala 40:20]
  wire [63:0] core_io_vme_rd_1_data_bits_data; // @[IntelShell.scala 40:20]
  wire [20:0] core_io_vme_rd_1_data_bits_tag; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_1_data_bits_last; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_2_cmd_ready; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_2_cmd_valid; // @[IntelShell.scala 40:20]
  wire [31:0] core_io_vme_rd_2_cmd_bits_addr; // @[IntelShell.scala 40:20]
  wire [3:0] core_io_vme_rd_2_cmd_bits_len; // @[IntelShell.scala 40:20]
  wire [20:0] core_io_vme_rd_2_cmd_bits_tag; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_2_data_valid; // @[IntelShell.scala 40:20]
  wire [63:0] core_io_vme_rd_2_data_bits_data; // @[IntelShell.scala 40:20]
  wire [20:0] core_io_vme_rd_2_data_bits_tag; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_3_cmd_ready; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_3_cmd_valid; // @[IntelShell.scala 40:20]
  wire [31:0] core_io_vme_rd_3_cmd_bits_addr; // @[IntelShell.scala 40:20]
  wire [3:0] core_io_vme_rd_3_cmd_bits_len; // @[IntelShell.scala 40:20]
  wire [20:0] core_io_vme_rd_3_cmd_bits_tag; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_3_data_valid; // @[IntelShell.scala 40:20]
  wire [63:0] core_io_vme_rd_3_data_bits_data; // @[IntelShell.scala 40:20]
  wire [20:0] core_io_vme_rd_3_data_bits_tag; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_4_cmd_ready; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_4_cmd_valid; // @[IntelShell.scala 40:20]
  wire [31:0] core_io_vme_rd_4_cmd_bits_addr; // @[IntelShell.scala 40:20]
  wire [3:0] core_io_vme_rd_4_cmd_bits_len; // @[IntelShell.scala 40:20]
  wire [20:0] core_io_vme_rd_4_cmd_bits_tag; // @[IntelShell.scala 40:20]
  wire  core_io_vme_rd_4_data_valid; // @[IntelShell.scala 40:20]
  wire [63:0] core_io_vme_rd_4_data_bits_data; // @[IntelShell.scala 40:20]
  wire [20:0] core_io_vme_rd_4_data_bits_tag; // @[IntelShell.scala 40:20]
  wire  core_io_vme_wr_0_cmd_ready; // @[IntelShell.scala 40:20]
  wire  core_io_vme_wr_0_cmd_valid; // @[IntelShell.scala 40:20]
  wire [31:0] core_io_vme_wr_0_cmd_bits_addr; // @[IntelShell.scala 40:20]
  wire [3:0] core_io_vme_wr_0_cmd_bits_len; // @[IntelShell.scala 40:20]
  wire  core_io_vme_wr_0_data_ready; // @[IntelShell.scala 40:20]
  wire  core_io_vme_wr_0_data_valid; // @[IntelShell.scala 40:20]
  wire [63:0] core_io_vme_wr_0_data_bits_data; // @[IntelShell.scala 40:20]
  wire  core_io_vme_wr_0_ack; // @[IntelShell.scala 40:20]
  VCR vcr ( // @[IntelShell.scala 38:19]
    .clock(vcr_clock),
    .reset(vcr_reset),
    .io_host_aw_ready(vcr_io_host_aw_ready),
    .io_host_aw_valid(vcr_io_host_aw_valid),
    .io_host_aw_bits_addr(vcr_io_host_aw_bits_addr),
    .io_host_w_ready(vcr_io_host_w_ready),
    .io_host_w_valid(vcr_io_host_w_valid),
    .io_host_w_bits_data(vcr_io_host_w_bits_data),
    .io_host_b_ready(vcr_io_host_b_ready),
    .io_host_b_valid(vcr_io_host_b_valid),
    .io_host_ar_ready(vcr_io_host_ar_ready),
    .io_host_ar_valid(vcr_io_host_ar_valid),
    .io_host_ar_bits_addr(vcr_io_host_ar_bits_addr),
    .io_host_r_ready(vcr_io_host_r_ready),
    .io_host_r_valid(vcr_io_host_r_valid),
    .io_host_r_bits_data(vcr_io_host_r_bits_data),
    .io_vcr_launch(vcr_io_vcr_launch),
    .io_vcr_finish(vcr_io_vcr_finish),
    .io_vcr_ecnt_0_valid(vcr_io_vcr_ecnt_0_valid),
    .io_vcr_ecnt_0_bits(vcr_io_vcr_ecnt_0_bits),
    .io_vcr_vals_0(vcr_io_vcr_vals_0),
    .io_vcr_ptrs_0(vcr_io_vcr_ptrs_0),
    .io_vcr_ptrs_1(vcr_io_vcr_ptrs_1),
    .io_vcr_ptrs_2(vcr_io_vcr_ptrs_2),
    .io_vcr_ptrs_3(vcr_io_vcr_ptrs_3),
    .io_vcr_ptrs_4(vcr_io_vcr_ptrs_4),
    .io_vcr_ptrs_5(vcr_io_vcr_ptrs_5),
    .io_vcr_ucnt_0_valid(vcr_io_vcr_ucnt_0_valid),
    .io_vcr_ucnt_0_bits(vcr_io_vcr_ucnt_0_bits)
  );
  VME vme ( // @[IntelShell.scala 39:19]
    .clock(vme_clock),
    .reset(vme_reset),
    .io_mem_aw_ready(vme_io_mem_aw_ready),
    .io_mem_aw_valid(vme_io_mem_aw_valid),
    .io_mem_aw_bits_addr(vme_io_mem_aw_bits_addr),
    .io_mem_aw_bits_len(vme_io_mem_aw_bits_len),
    .io_mem_w_ready(vme_io_mem_w_ready),
    .io_mem_w_valid(vme_io_mem_w_valid),
    .io_mem_w_bits_data(vme_io_mem_w_bits_data),
    .io_mem_w_bits_last(vme_io_mem_w_bits_last),
    .io_mem_b_ready(vme_io_mem_b_ready),
    .io_mem_b_valid(vme_io_mem_b_valid),
    .io_mem_ar_ready(vme_io_mem_ar_ready),
    .io_mem_ar_valid(vme_io_mem_ar_valid),
    .io_mem_ar_bits_addr(vme_io_mem_ar_bits_addr),
    .io_mem_ar_bits_id(vme_io_mem_ar_bits_id),
    .io_mem_ar_bits_len(vme_io_mem_ar_bits_len),
    .io_mem_r_valid(vme_io_mem_r_valid),
    .io_mem_r_bits_data(vme_io_mem_r_bits_data),
    .io_mem_r_bits_last(vme_io_mem_r_bits_last),
    .io_mem_r_bits_id(vme_io_mem_r_bits_id),
    .io_vme_rd_0_cmd_ready(vme_io_vme_rd_0_cmd_ready),
    .io_vme_rd_0_cmd_valid(vme_io_vme_rd_0_cmd_valid),
    .io_vme_rd_0_cmd_bits_addr(vme_io_vme_rd_0_cmd_bits_addr),
    .io_vme_rd_0_cmd_bits_len(vme_io_vme_rd_0_cmd_bits_len),
    .io_vme_rd_0_data_ready(vme_io_vme_rd_0_data_ready),
    .io_vme_rd_0_data_valid(vme_io_vme_rd_0_data_valid),
    .io_vme_rd_0_data_bits_data(vme_io_vme_rd_0_data_bits_data),
    .io_vme_rd_1_cmd_ready(vme_io_vme_rd_1_cmd_ready),
    .io_vme_rd_1_cmd_valid(vme_io_vme_rd_1_cmd_valid),
    .io_vme_rd_1_cmd_bits_addr(vme_io_vme_rd_1_cmd_bits_addr),
    .io_vme_rd_1_cmd_bits_len(vme_io_vme_rd_1_cmd_bits_len),
    .io_vme_rd_1_cmd_bits_tag(vme_io_vme_rd_1_cmd_bits_tag),
    .io_vme_rd_1_data_valid(vme_io_vme_rd_1_data_valid),
    .io_vme_rd_1_data_bits_data(vme_io_vme_rd_1_data_bits_data),
    .io_vme_rd_1_data_bits_tag(vme_io_vme_rd_1_data_bits_tag),
    .io_vme_rd_1_data_bits_last(vme_io_vme_rd_1_data_bits_last),
    .io_vme_rd_2_cmd_ready(vme_io_vme_rd_2_cmd_ready),
    .io_vme_rd_2_cmd_valid(vme_io_vme_rd_2_cmd_valid),
    .io_vme_rd_2_cmd_bits_addr(vme_io_vme_rd_2_cmd_bits_addr),
    .io_vme_rd_2_cmd_bits_len(vme_io_vme_rd_2_cmd_bits_len),
    .io_vme_rd_2_cmd_bits_tag(vme_io_vme_rd_2_cmd_bits_tag),
    .io_vme_rd_2_data_valid(vme_io_vme_rd_2_data_valid),
    .io_vme_rd_2_data_bits_data(vme_io_vme_rd_2_data_bits_data),
    .io_vme_rd_2_data_bits_tag(vme_io_vme_rd_2_data_bits_tag),
    .io_vme_rd_3_cmd_ready(vme_io_vme_rd_3_cmd_ready),
    .io_vme_rd_3_cmd_valid(vme_io_vme_rd_3_cmd_valid),
    .io_vme_rd_3_cmd_bits_addr(vme_io_vme_rd_3_cmd_bits_addr),
    .io_vme_rd_3_cmd_bits_len(vme_io_vme_rd_3_cmd_bits_len),
    .io_vme_rd_3_cmd_bits_tag(vme_io_vme_rd_3_cmd_bits_tag),
    .io_vme_rd_3_data_valid(vme_io_vme_rd_3_data_valid),
    .io_vme_rd_3_data_bits_data(vme_io_vme_rd_3_data_bits_data),
    .io_vme_rd_3_data_bits_tag(vme_io_vme_rd_3_data_bits_tag),
    .io_vme_rd_4_cmd_ready(vme_io_vme_rd_4_cmd_ready),
    .io_vme_rd_4_cmd_valid(vme_io_vme_rd_4_cmd_valid),
    .io_vme_rd_4_cmd_bits_addr(vme_io_vme_rd_4_cmd_bits_addr),
    .io_vme_rd_4_cmd_bits_len(vme_io_vme_rd_4_cmd_bits_len),
    .io_vme_rd_4_cmd_bits_tag(vme_io_vme_rd_4_cmd_bits_tag),
    .io_vme_rd_4_data_valid(vme_io_vme_rd_4_data_valid),
    .io_vme_rd_4_data_bits_data(vme_io_vme_rd_4_data_bits_data),
    .io_vme_rd_4_data_bits_tag(vme_io_vme_rd_4_data_bits_tag),
    .io_vme_wr_0_cmd_ready(vme_io_vme_wr_0_cmd_ready),
    .io_vme_wr_0_cmd_valid(vme_io_vme_wr_0_cmd_valid),
    .io_vme_wr_0_cmd_bits_addr(vme_io_vme_wr_0_cmd_bits_addr),
    .io_vme_wr_0_cmd_bits_len(vme_io_vme_wr_0_cmd_bits_len),
    .io_vme_wr_0_data_ready(vme_io_vme_wr_0_data_ready),
    .io_vme_wr_0_data_valid(vme_io_vme_wr_0_data_valid),
    .io_vme_wr_0_data_bits_data(vme_io_vme_wr_0_data_bits_data),
    .io_vme_wr_0_ack(vme_io_vme_wr_0_ack)
  );
  Core core ( // @[IntelShell.scala 40:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_vcr_launch(core_io_vcr_launch),
    .io_vcr_finish(core_io_vcr_finish),
    .io_vcr_ecnt_0_valid(core_io_vcr_ecnt_0_valid),
    .io_vcr_ecnt_0_bits(core_io_vcr_ecnt_0_bits),
    .io_vcr_vals_0(core_io_vcr_vals_0),
    .io_vcr_ptrs_0(core_io_vcr_ptrs_0),
    .io_vcr_ptrs_1(core_io_vcr_ptrs_1),
    .io_vcr_ptrs_2(core_io_vcr_ptrs_2),
    .io_vcr_ptrs_3(core_io_vcr_ptrs_3),
    .io_vcr_ptrs_4(core_io_vcr_ptrs_4),
    .io_vcr_ptrs_5(core_io_vcr_ptrs_5),
    .io_vcr_ucnt_0_valid(core_io_vcr_ucnt_0_valid),
    .io_vcr_ucnt_0_bits(core_io_vcr_ucnt_0_bits),
    .io_vme_rd_0_cmd_ready(core_io_vme_rd_0_cmd_ready),
    .io_vme_rd_0_cmd_valid(core_io_vme_rd_0_cmd_valid),
    .io_vme_rd_0_cmd_bits_addr(core_io_vme_rd_0_cmd_bits_addr),
    .io_vme_rd_0_cmd_bits_len(core_io_vme_rd_0_cmd_bits_len),
    .io_vme_rd_0_data_ready(core_io_vme_rd_0_data_ready),
    .io_vme_rd_0_data_valid(core_io_vme_rd_0_data_valid),
    .io_vme_rd_0_data_bits_data(core_io_vme_rd_0_data_bits_data),
    .io_vme_rd_1_cmd_ready(core_io_vme_rd_1_cmd_ready),
    .io_vme_rd_1_cmd_valid(core_io_vme_rd_1_cmd_valid),
    .io_vme_rd_1_cmd_bits_addr(core_io_vme_rd_1_cmd_bits_addr),
    .io_vme_rd_1_cmd_bits_len(core_io_vme_rd_1_cmd_bits_len),
    .io_vme_rd_1_cmd_bits_tag(core_io_vme_rd_1_cmd_bits_tag),
    .io_vme_rd_1_data_valid(core_io_vme_rd_1_data_valid),
    .io_vme_rd_1_data_bits_data(core_io_vme_rd_1_data_bits_data),
    .io_vme_rd_1_data_bits_tag(core_io_vme_rd_1_data_bits_tag),
    .io_vme_rd_1_data_bits_last(core_io_vme_rd_1_data_bits_last),
    .io_vme_rd_2_cmd_ready(core_io_vme_rd_2_cmd_ready),
    .io_vme_rd_2_cmd_valid(core_io_vme_rd_2_cmd_valid),
    .io_vme_rd_2_cmd_bits_addr(core_io_vme_rd_2_cmd_bits_addr),
    .io_vme_rd_2_cmd_bits_len(core_io_vme_rd_2_cmd_bits_len),
    .io_vme_rd_2_cmd_bits_tag(core_io_vme_rd_2_cmd_bits_tag),
    .io_vme_rd_2_data_valid(core_io_vme_rd_2_data_valid),
    .io_vme_rd_2_data_bits_data(core_io_vme_rd_2_data_bits_data),
    .io_vme_rd_2_data_bits_tag(core_io_vme_rd_2_data_bits_tag),
    .io_vme_rd_3_cmd_ready(core_io_vme_rd_3_cmd_ready),
    .io_vme_rd_3_cmd_valid(core_io_vme_rd_3_cmd_valid),
    .io_vme_rd_3_cmd_bits_addr(core_io_vme_rd_3_cmd_bits_addr),
    .io_vme_rd_3_cmd_bits_len(core_io_vme_rd_3_cmd_bits_len),
    .io_vme_rd_3_cmd_bits_tag(core_io_vme_rd_3_cmd_bits_tag),
    .io_vme_rd_3_data_valid(core_io_vme_rd_3_data_valid),
    .io_vme_rd_3_data_bits_data(core_io_vme_rd_3_data_bits_data),
    .io_vme_rd_3_data_bits_tag(core_io_vme_rd_3_data_bits_tag),
    .io_vme_rd_4_cmd_ready(core_io_vme_rd_4_cmd_ready),
    .io_vme_rd_4_cmd_valid(core_io_vme_rd_4_cmd_valid),
    .io_vme_rd_4_cmd_bits_addr(core_io_vme_rd_4_cmd_bits_addr),
    .io_vme_rd_4_cmd_bits_len(core_io_vme_rd_4_cmd_bits_len),
    .io_vme_rd_4_cmd_bits_tag(core_io_vme_rd_4_cmd_bits_tag),
    .io_vme_rd_4_data_valid(core_io_vme_rd_4_data_valid),
    .io_vme_rd_4_data_bits_data(core_io_vme_rd_4_data_bits_data),
    .io_vme_rd_4_data_bits_tag(core_io_vme_rd_4_data_bits_tag),
    .io_vme_wr_0_cmd_ready(core_io_vme_wr_0_cmd_ready),
    .io_vme_wr_0_cmd_valid(core_io_vme_wr_0_cmd_valid),
    .io_vme_wr_0_cmd_bits_addr(core_io_vme_wr_0_cmd_bits_addr),
    .io_vme_wr_0_cmd_bits_len(core_io_vme_wr_0_cmd_bits_len),
    .io_vme_wr_0_data_ready(core_io_vme_wr_0_data_ready),
    .io_vme_wr_0_data_valid(core_io_vme_wr_0_data_valid),
    .io_vme_wr_0_data_bits_data(core_io_vme_wr_0_data_bits_data),
    .io_vme_wr_0_ack(core_io_vme_wr_0_ack)
  );
  assign io_host_aw_ready = vcr_io_host_aw_ready; // @[IntelShell.scala 46:20]
  assign io_host_w_ready = vcr_io_host_w_ready; // @[IntelShell.scala 49:19]
  assign io_host_b_valid = vcr_io_host_b_valid; // @[IntelShell.scala 54:19]
  assign io_host_b_bits_resp = 2'h0; // @[IntelShell.scala 55:23]
  assign io_host_b_bits_id = io_host_w_bits_id; // @[IntelShell.scala 56:21]
  assign io_host_b_bits_user = 1'h0;
  assign io_host_ar_ready = vcr_io_host_ar_ready; // @[IntelShell.scala 58:20]
  assign io_host_r_valid = vcr_io_host_r_valid; // @[IntelShell.scala 62:19]
  assign io_host_r_bits_data = vcr_io_host_r_bits_data; // @[IntelShell.scala 63:23]
  assign io_host_r_bits_resp = 2'h0; // @[IntelShell.scala 64:23]
  assign io_host_r_bits_last = 1'h1; // @[IntelShell.scala 69:23]
  assign io_host_r_bits_id = io_host_ar_bits_id; // @[IntelShell.scala 65:21]
  assign io_host_r_bits_user = 1'h0;
  assign io_mem_aw_valid = vme_io_mem_aw_valid; // @[IntelShell.scala 71:10]
  assign io_mem_aw_bits_addr = vme_io_mem_aw_bits_addr; // @[IntelShell.scala 71:10]
  assign io_mem_aw_bits_id = 8'h0; // @[IntelShell.scala 71:10]
  assign io_mem_aw_bits_user = 5'h1; // @[IntelShell.scala 71:10]
  assign io_mem_aw_bits_len = vme_io_mem_aw_bits_len; // @[IntelShell.scala 71:10]
  assign io_mem_aw_bits_size = 3'h3; // @[IntelShell.scala 71:10]
  assign io_mem_aw_bits_burst = 2'h1; // @[IntelShell.scala 71:10]
  assign io_mem_aw_bits_lock = 2'h0; // @[IntelShell.scala 71:10]
  assign io_mem_aw_bits_cache = 4'hf; // @[IntelShell.scala 71:10]
  assign io_mem_aw_bits_prot = 3'h4; // @[IntelShell.scala 71:10]
  assign io_mem_aw_bits_qos = 4'h0; // @[IntelShell.scala 71:10]
  assign io_mem_aw_bits_region = 4'h0; // @[IntelShell.scala 71:10]
  assign io_mem_w_valid = vme_io_mem_w_valid; // @[IntelShell.scala 71:10]
  assign io_mem_w_bits_data = vme_io_mem_w_bits_data; // @[IntelShell.scala 71:10]
  assign io_mem_w_bits_strb = 8'hff; // @[IntelShell.scala 71:10]
  assign io_mem_w_bits_last = vme_io_mem_w_bits_last; // @[IntelShell.scala 71:10]
  assign io_mem_w_bits_id = 8'h0; // @[IntelShell.scala 71:10]
  assign io_mem_w_bits_user = 5'h1; // @[IntelShell.scala 71:10]
  assign io_mem_b_ready = vme_io_mem_b_ready; // @[IntelShell.scala 71:10]
  assign io_mem_ar_valid = vme_io_mem_ar_valid; // @[IntelShell.scala 71:10]
  assign io_mem_ar_bits_addr = vme_io_mem_ar_bits_addr; // @[IntelShell.scala 71:10]
  assign io_mem_ar_bits_id = vme_io_mem_ar_bits_id; // @[IntelShell.scala 71:10]
  assign io_mem_ar_bits_user = 5'h1; // @[IntelShell.scala 71:10]
  assign io_mem_ar_bits_len = vme_io_mem_ar_bits_len; // @[IntelShell.scala 71:10]
  assign io_mem_ar_bits_size = 3'h3; // @[IntelShell.scala 71:10]
  assign io_mem_ar_bits_burst = 2'h1; // @[IntelShell.scala 71:10]
  assign io_mem_ar_bits_lock = 2'h0; // @[IntelShell.scala 71:10]
  assign io_mem_ar_bits_cache = 4'hf; // @[IntelShell.scala 71:10]
  assign io_mem_ar_bits_prot = 3'h4; // @[IntelShell.scala 71:10]
  assign io_mem_ar_bits_qos = 4'h0; // @[IntelShell.scala 71:10]
  assign io_mem_ar_bits_region = 4'h0; // @[IntelShell.scala 71:10]
  assign io_mem_r_ready = 1'h1; // @[IntelShell.scala 71:10]
  assign vcr_clock = clock;
  assign vcr_reset = reset;
  assign vcr_io_host_aw_valid = io_host_aw_valid; // @[IntelShell.scala 47:24]
  assign vcr_io_host_aw_bits_addr = io_host_aw_bits_addr; // @[IntelShell.scala 48:28]
  assign vcr_io_host_w_valid = io_host_w_valid; // @[IntelShell.scala 50:23]
  assign vcr_io_host_w_bits_data = io_host_w_bits_data; // @[IntelShell.scala 51:27]
  assign vcr_io_host_b_ready = io_host_b_ready; // @[IntelShell.scala 53:23]
  assign vcr_io_host_ar_valid = io_host_ar_valid; // @[IntelShell.scala 59:24]
  assign vcr_io_host_ar_bits_addr = io_host_ar_bits_addr; // @[IntelShell.scala 60:28]
  assign vcr_io_host_r_ready = io_host_r_ready; // @[IntelShell.scala 61:23]
  assign vcr_io_vcr_finish = core_io_vcr_finish; // @[IntelShell.scala 42:15]
  assign vcr_io_vcr_ecnt_0_valid = core_io_vcr_ecnt_0_valid; // @[IntelShell.scala 42:15]
  assign vcr_io_vcr_ecnt_0_bits = core_io_vcr_ecnt_0_bits; // @[IntelShell.scala 42:15]
  assign vcr_io_vcr_ucnt_0_valid = core_io_vcr_ucnt_0_valid; // @[IntelShell.scala 42:15]
  assign vcr_io_vcr_ucnt_0_bits = core_io_vcr_ucnt_0_bits; // @[IntelShell.scala 42:15]
  assign vme_clock = clock;
  assign vme_reset = reset;
  assign vme_io_mem_aw_ready = io_mem_aw_ready; // @[IntelShell.scala 71:10]
  assign vme_io_mem_w_ready = io_mem_w_ready; // @[IntelShell.scala 71:10]
  assign vme_io_mem_b_valid = io_mem_b_valid; // @[IntelShell.scala 71:10]
  assign vme_io_mem_ar_ready = io_mem_ar_ready; // @[IntelShell.scala 71:10]
  assign vme_io_mem_r_valid = io_mem_r_valid; // @[IntelShell.scala 71:10]
  assign vme_io_mem_r_bits_data = io_mem_r_bits_data; // @[IntelShell.scala 71:10]
  assign vme_io_mem_r_bits_last = io_mem_r_bits_last; // @[IntelShell.scala 71:10]
  assign vme_io_mem_r_bits_id = io_mem_r_bits_id; // @[IntelShell.scala 71:10]
  assign vme_io_vme_rd_0_cmd_valid = core_io_vme_rd_0_cmd_valid; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_0_cmd_bits_addr = core_io_vme_rd_0_cmd_bits_addr; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_0_cmd_bits_len = core_io_vme_rd_0_cmd_bits_len; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_0_data_ready = core_io_vme_rd_0_data_ready; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_1_cmd_valid = core_io_vme_rd_1_cmd_valid; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_1_cmd_bits_addr = core_io_vme_rd_1_cmd_bits_addr; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_1_cmd_bits_len = core_io_vme_rd_1_cmd_bits_len; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_1_cmd_bits_tag = core_io_vme_rd_1_cmd_bits_tag; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_2_cmd_valid = core_io_vme_rd_2_cmd_valid; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_2_cmd_bits_addr = core_io_vme_rd_2_cmd_bits_addr; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_2_cmd_bits_len = core_io_vme_rd_2_cmd_bits_len; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_2_cmd_bits_tag = core_io_vme_rd_2_cmd_bits_tag; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_3_cmd_valid = core_io_vme_rd_3_cmd_valid; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_3_cmd_bits_addr = core_io_vme_rd_3_cmd_bits_addr; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_3_cmd_bits_len = core_io_vme_rd_3_cmd_bits_len; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_3_cmd_bits_tag = core_io_vme_rd_3_cmd_bits_tag; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_4_cmd_valid = core_io_vme_rd_4_cmd_valid; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_4_cmd_bits_addr = core_io_vme_rd_4_cmd_bits_addr; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_4_cmd_bits_len = core_io_vme_rd_4_cmd_bits_len; // @[IntelShell.scala 43:14]
  assign vme_io_vme_rd_4_cmd_bits_tag = core_io_vme_rd_4_cmd_bits_tag; // @[IntelShell.scala 43:14]
  assign vme_io_vme_wr_0_cmd_valid = core_io_vme_wr_0_cmd_valid; // @[IntelShell.scala 43:14]
  assign vme_io_vme_wr_0_cmd_bits_addr = core_io_vme_wr_0_cmd_bits_addr; // @[IntelShell.scala 43:14]
  assign vme_io_vme_wr_0_cmd_bits_len = core_io_vme_wr_0_cmd_bits_len; // @[IntelShell.scala 43:14]
  assign vme_io_vme_wr_0_data_valid = core_io_vme_wr_0_data_valid; // @[IntelShell.scala 43:14]
  assign vme_io_vme_wr_0_data_bits_data = core_io_vme_wr_0_data_bits_data; // @[IntelShell.scala 43:14]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_vcr_launch = vcr_io_vcr_launch; // @[IntelShell.scala 42:15]
  assign core_io_vcr_vals_0 = vcr_io_vcr_vals_0; // @[IntelShell.scala 42:15]
  assign core_io_vcr_ptrs_0 = vcr_io_vcr_ptrs_0; // @[IntelShell.scala 42:15]
  assign core_io_vcr_ptrs_1 = vcr_io_vcr_ptrs_1; // @[IntelShell.scala 42:15]
  assign core_io_vcr_ptrs_2 = vcr_io_vcr_ptrs_2; // @[IntelShell.scala 42:15]
  assign core_io_vcr_ptrs_3 = vcr_io_vcr_ptrs_3; // @[IntelShell.scala 42:15]
  assign core_io_vcr_ptrs_4 = vcr_io_vcr_ptrs_4; // @[IntelShell.scala 42:15]
  assign core_io_vcr_ptrs_5 = vcr_io_vcr_ptrs_5; // @[IntelShell.scala 42:15]
  assign core_io_vme_rd_0_cmd_ready = vme_io_vme_rd_0_cmd_ready; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_0_data_valid = vme_io_vme_rd_0_data_valid; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_0_data_bits_data = vme_io_vme_rd_0_data_bits_data; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_1_cmd_ready = vme_io_vme_rd_1_cmd_ready; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_1_data_valid = vme_io_vme_rd_1_data_valid; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_1_data_bits_data = vme_io_vme_rd_1_data_bits_data; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_1_data_bits_tag = vme_io_vme_rd_1_data_bits_tag; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_1_data_bits_last = vme_io_vme_rd_1_data_bits_last; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_2_cmd_ready = vme_io_vme_rd_2_cmd_ready; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_2_data_valid = vme_io_vme_rd_2_data_valid; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_2_data_bits_data = vme_io_vme_rd_2_data_bits_data; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_2_data_bits_tag = vme_io_vme_rd_2_data_bits_tag; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_3_cmd_ready = vme_io_vme_rd_3_cmd_ready; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_3_data_valid = vme_io_vme_rd_3_data_valid; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_3_data_bits_data = vme_io_vme_rd_3_data_bits_data; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_3_data_bits_tag = vme_io_vme_rd_3_data_bits_tag; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_4_cmd_ready = vme_io_vme_rd_4_cmd_ready; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_4_data_valid = vme_io_vme_rd_4_data_valid; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_4_data_bits_data = vme_io_vme_rd_4_data_bits_data; // @[IntelShell.scala 43:14]
  assign core_io_vme_rd_4_data_bits_tag = vme_io_vme_rd_4_data_bits_tag; // @[IntelShell.scala 43:14]
  assign core_io_vme_wr_0_cmd_ready = vme_io_vme_wr_0_cmd_ready; // @[IntelShell.scala 43:14]
  assign core_io_vme_wr_0_data_ready = vme_io_vme_wr_0_data_ready; // @[IntelShell.scala 43:14]
  assign core_io_vme_wr_0_ack = vme_io_vme_wr_0_ack; // @[IntelShell.scala 43:14]
endmodule
