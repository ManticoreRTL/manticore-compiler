module ProcessingElement(
  input         clock,
  input         reset,
  output        io_left_in_ready,
  input         io_left_in_valid,
  input  [31:0] io_left_in_bits,
  output        io_top_in_ready,
  input         io_top_in_valid,
  input  [31:0] io_top_in_bits,
  input         io_sum_ready,
  output        io_sum_valid,
  output [31:0] io_sum_bits,
  input         io_right_out_ready,
  output        io_right_out_valid,
  output [31:0] io_right_out_bits,
  input         io_bottom_out_ready,
  output        io_bottom_out_valid,
  output [31:0] io_bottom_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [15:0] value; // @[Counter.scala 62:40]
  reg [31:0] acc; // @[Stab.scala 24:20]
  reg [1:0] state; // @[Stab.scala 27:50]
  wire [63:0] mul = io_left_in_bits * io_top_in_bits; // @[Stab.scala 28:71]
  wire  _T_1 = io_left_in_valid & io_top_in_valid; // @[Stab.scala 45:29]
  wire  _T_5 = _T_1 & io_right_out_ready & io_bottom_out_ready; // @[Stab.scala 50:70]
  wire [63:0] _GEN_31 = {{32'd0}, acc}; // @[Stab.scala 51:36]
  wire [63:0] _acc_T_1 = _GEN_31 + mul; // @[Stab.scala 51:36]
  wire  wrap = value == 16'hfffe; // @[Counter.scala 74:24]
  wire [15:0] _value_T_1 = value + 16'h1; // @[Counter.scala 78:24]
  wire [15:0] _GEN_2 = wrap ? 16'h0 : _value_T_1; // @[Counter.scala 78:15 88:{20,28}]
  wire [15:0] _T_7 = 16'h10 - 16'h1; // @[Stab.scala 55:48]
  wire [1:0] _GEN_3 = value == _T_7 ? 2'h2 : state; // @[Stab.scala 55:56 56:17 27:50]
  wire [63:0] _GEN_4 = _T_1 & io_right_out_ready & io_bottom_out_ready ? _acc_T_1 : {{32'd0}, acc}; // @[Stab.scala 24:20 50:94 51:29]
  wire [31:0] _GEN_10 = io_sum_ready ? 32'h0 : acc; // @[Stab.scala 24:20 61:26 64:22]
  wire [1:0] _GEN_11 = io_sum_ready ? 2'h0 : state; // @[Stab.scala 61:26 65:22 27:50]
  wire [15:0] _GEN_12 = io_sum_ready ? 16'h0 : value; // @[Stab.scala 61:26 Counter.scala 99:11 62:40]
  wire [31:0] _GEN_15 = 2'h2 == state ? _GEN_10 : acc; // @[Stab.scala 40:17 24:20]
  wire [63:0] _GEN_18 = 2'h1 == state ? _GEN_4 : {{32'd0}, _GEN_15}; // @[Stab.scala 40:17]
  wire  _GEN_22 = 2'h1 == state ? 1'h0 : 2'h2 == state & io_sum_ready; // @[Stab.scala 38:16 40:17]
  wire [63:0] _GEN_26 = 2'h0 == state ? {{32'd0}, acc} : _GEN_18; // @[Stab.scala 40:17 24:20]
  wire [63:0] _GEN_32 = reset ? 64'h0 : _GEN_26; // @[Stab.scala 24:{20,20}]
  assign io_left_in_ready = state == 2'h1; // @[Stab.scala 30:33]
  assign io_top_in_ready = state == 2'h1; // @[Stab.scala 31:33]
  assign io_sum_valid = 2'h0 == state ? 1'h0 : _GEN_22; // @[Stab.scala 38:16 40:17]
  assign io_sum_bits = acc; // @[Stab.scala 39:16 40:17]
  assign io_right_out_valid = 2'h0 == state ? 1'h0 : 2'h1 == state & _T_5; // @[Stab.scala 40:17 33:23]
  assign io_right_out_bits = io_left_in_bits; // @[Stab.scala 36:22]
  assign io_bottom_out_valid = 2'h0 == state ? 1'h0 : 2'h1 == state & _T_5; // @[Stab.scala 40:17 33:23]
  assign io_bottom_out_bits = io_top_in_bits; // @[Stab.scala 35:22]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 62:40]
      value <= 16'h0; // @[Counter.scala 62:40]
    end else if (!(2'h0 == state)) begin // @[Stab.scala 40:17]
      if (2'h1 == state) begin // @[Stab.scala 40:17]
        if (_T_1 & io_right_out_ready & io_bottom_out_ready) begin // @[Stab.scala 50:94]
          value <= _GEN_2;
        end
      end else if (2'h2 == state) begin // @[Stab.scala 40:17]
        value <= _GEN_12;
      end
    end
    acc <= _GEN_32[31:0]; // @[Stab.scala 24:{20,20}]
    if (reset) begin // @[Stab.scala 27:50]
      state <= 2'h0; // @[Stab.scala 27:50]
    end else if (2'h0 == state) begin // @[Stab.scala 40:17]
      if (io_left_in_valid & io_top_in_valid) begin // @[Stab.scala 45:49]
        state <= 2'h1; // @[Stab.scala 46:15]
      end
    end else if (2'h1 == state) begin // @[Stab.scala 40:17]
      if (_T_1 & io_right_out_ready & io_bottom_out_ready) begin // @[Stab.scala 50:94]
        state <= _GEN_3;
      end
    end else if (2'h2 == state) begin // @[Stab.scala 40:17]
      state <= _GEN_11;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[15:0];
  _RAND_1 = {1{`RANDOM}};
  acc = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Queue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] ram [0:3]; // @[Decoupled.scala 259:44]
  wire  ram_io_deq_bits_MPORT_en; // @[Decoupled.scala 259:44]
  wire [1:0] ram_io_deq_bits_MPORT_addr; // @[Decoupled.scala 259:44]
  wire [31:0] ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 259:44]
  wire [31:0] ram_MPORT_data; // @[Decoupled.scala 259:44]
  wire [1:0] ram_MPORT_addr; // @[Decoupled.scala 259:44]
  wire  ram_MPORT_mask; // @[Decoupled.scala 259:44]
  wire  ram_MPORT_en; // @[Decoupled.scala 259:44]
  reg  ram_io_deq_bits_MPORT_en_pipe_0;
  reg [1:0] ram_io_deq_bits_MPORT_addr_pipe_0;
  reg [1:0] value; // @[Counter.scala 62:40]
  reg [1:0] value_1; // @[Counter.scala 62:40]
  reg  maybe_full; // @[Decoupled.scala 262:27]
  wire  ptr_match = value == value_1; // @[Decoupled.scala 263:33]
  wire  empty = ptr_match & ~maybe_full; // @[Decoupled.scala 264:25]
  wire  full = ptr_match & maybe_full; // @[Decoupled.scala 265:24]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _value_T_1 = value + 2'h1; // @[Counter.scala 78:24]
  wire [1:0] _value_T_3 = value_1 + 2'h1; // @[Counter.scala 78:24]
  wire [2:0] _deq_ptr_next_T_1 = 3'h4 - 3'h1; // @[Decoupled.scala 292:57]
  wire [2:0] _GEN_15 = {{1'd0}, value_1}; // @[Decoupled.scala 292:42]
  assign ram_io_deq_bits_MPORT_en = ram_io_deq_bits_MPORT_en_pipe_0;
  assign ram_io_deq_bits_MPORT_addr = ram_io_deq_bits_MPORT_addr_pipe_0;
  assign ram_io_deq_bits_MPORT_data = ram[ram_io_deq_bits_MPORT_addr]; // @[Decoupled.scala 259:44]
  assign ram_MPORT_data = io_enq_bits;
  assign ram_MPORT_addr = value;
  assign ram_MPORT_mask = 1'h1;
  assign ram_MPORT_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~full; // @[Decoupled.scala 289:19]
  assign io_deq_valid = ~empty; // @[Decoupled.scala 288:19]
  assign io_deq_bits = ram_io_deq_bits_MPORT_data; // @[Decoupled.scala 294:17]
  always @(posedge clock) begin
    if (ram_MPORT_en & ram_MPORT_mask) begin
      ram[ram_MPORT_addr] <= ram_MPORT_data; // @[Decoupled.scala 259:44]
    end
    ram_io_deq_bits_MPORT_en_pipe_0 <= 1'h1;
    if (1'h1) begin
      if (do_deq) begin
        if (_GEN_15 == _deq_ptr_next_T_1) begin // @[Decoupled.scala 292:27]
          ram_io_deq_bits_MPORT_addr_pipe_0 <= 2'h0;
        end else begin
          ram_io_deq_bits_MPORT_addr_pipe_0 <= _value_T_3;
        end
      end else begin
        ram_io_deq_bits_MPORT_addr_pipe_0 <= value_1;
      end
    end
    if (reset) begin // @[Counter.scala 62:40]
      value <= 2'h0; // @[Counter.scala 62:40]
    end else if (do_enq) begin // @[Decoupled.scala 272:16]
      value <= _value_T_1; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Counter.scala 62:40]
      value_1 <= 2'h0; // @[Counter.scala 62:40]
    end else if (do_deq) begin // @[Decoupled.scala 276:16]
      value_1 <= _value_T_3; // @[Counter.scala 78:15]
    end
    if (reset) begin // @[Decoupled.scala 262:27]
      maybe_full <= 1'h0; // @[Decoupled.scala 262:27]
    end else if (do_enq != do_deq) begin // @[Decoupled.scala 279:27]
      maybe_full <= do_enq; // @[Decoupled.scala 280:16]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_io_deq_bits_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_io_deq_bits_MPORT_addr_pipe_0 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  value = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  value_1 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  maybe_full = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BareMatrixMultiplier(
  input         clock,
  input         reset,
  output        io_weight_in_0_ready,
  input         io_weight_in_0_valid,
  input  [31:0] io_weight_in_0_bits,
  output        io_weight_in_1_ready,
  input         io_weight_in_1_valid,
  input  [31:0] io_weight_in_1_bits,
  output        io_weight_in_2_ready,
  input         io_weight_in_2_valid,
  input  [31:0] io_weight_in_2_bits,
  output        io_weight_in_3_ready,
  input         io_weight_in_3_valid,
  input  [31:0] io_weight_in_3_bits,
  output        io_weight_in_4_ready,
  input         io_weight_in_4_valid,
  input  [31:0] io_weight_in_4_bits,
  output        io_weight_in_5_ready,
  input         io_weight_in_5_valid,
  input  [31:0] io_weight_in_5_bits,
  output        io_weight_in_6_ready,
  input         io_weight_in_6_valid,
  input  [31:0] io_weight_in_6_bits,
  output        io_weight_in_7_ready,
  input         io_weight_in_7_valid,
  input  [31:0] io_weight_in_7_bits,
  output        io_weight_in_8_ready,
  input         io_weight_in_8_valid,
  input  [31:0] io_weight_in_8_bits,
  output        io_weight_in_9_ready,
  input         io_weight_in_9_valid,
  input  [31:0] io_weight_in_9_bits,
  output        io_weight_in_10_ready,
  input         io_weight_in_10_valid,
  input  [31:0] io_weight_in_10_bits,
  output        io_weight_in_11_ready,
  input         io_weight_in_11_valid,
  input  [31:0] io_weight_in_11_bits,
  output        io_weight_in_12_ready,
  input         io_weight_in_12_valid,
  input  [31:0] io_weight_in_12_bits,
  output        io_weight_in_13_ready,
  input         io_weight_in_13_valid,
  input  [31:0] io_weight_in_13_bits,
  output        io_weight_in_14_ready,
  input         io_weight_in_14_valid,
  input  [31:0] io_weight_in_14_bits,
  output        io_weight_in_15_ready,
  input         io_weight_in_15_valid,
  input  [31:0] io_weight_in_15_bits,
  output        io_value_in_0_ready,
  input         io_value_in_0_valid,
  input  [31:0] io_value_in_0_bits,
  output        io_value_in_1_ready,
  input         io_value_in_1_valid,
  input  [31:0] io_value_in_1_bits,
  output        io_value_in_2_ready,
  input         io_value_in_2_valid,
  input  [31:0] io_value_in_2_bits,
  output        io_value_in_3_ready,
  input         io_value_in_3_valid,
  input  [31:0] io_value_in_3_bits,
  output        io_value_in_4_ready,
  input         io_value_in_4_valid,
  input  [31:0] io_value_in_4_bits,
  output        io_value_in_5_ready,
  input         io_value_in_5_valid,
  input  [31:0] io_value_in_5_bits,
  output        io_value_in_6_ready,
  input         io_value_in_6_valid,
  input  [31:0] io_value_in_6_bits,
  output        io_value_in_7_ready,
  input         io_value_in_7_valid,
  input  [31:0] io_value_in_7_bits,
  output        io_value_in_8_ready,
  input         io_value_in_8_valid,
  input  [31:0] io_value_in_8_bits,
  output        io_value_in_9_ready,
  input         io_value_in_9_valid,
  input  [31:0] io_value_in_9_bits,
  output        io_value_in_10_ready,
  input         io_value_in_10_valid,
  input  [31:0] io_value_in_10_bits,
  output        io_value_in_11_ready,
  input         io_value_in_11_valid,
  input  [31:0] io_value_in_11_bits,
  output        io_value_in_12_ready,
  input         io_value_in_12_valid,
  input  [31:0] io_value_in_12_bits,
  output        io_value_in_13_ready,
  input         io_value_in_13_valid,
  input  [31:0] io_value_in_13_bits,
  output        io_value_in_14_ready,
  input         io_value_in_14_valid,
  input  [31:0] io_value_in_14_bits,
  output        io_value_in_15_ready,
  input         io_value_in_15_valid,
  input  [31:0] io_value_in_15_bits,
  input         io_value_out_0_0_ready,
  output        io_value_out_0_0_valid,
  output [31:0] io_value_out_0_0_bits,
  input         io_value_out_0_1_ready,
  output        io_value_out_0_1_valid,
  output [31:0] io_value_out_0_1_bits,
  input         io_value_out_0_2_ready,
  output        io_value_out_0_2_valid,
  output [31:0] io_value_out_0_2_bits,
  input         io_value_out_0_3_ready,
  output        io_value_out_0_3_valid,
  output [31:0] io_value_out_0_3_bits,
  input         io_value_out_0_4_ready,
  output        io_value_out_0_4_valid,
  output [31:0] io_value_out_0_4_bits,
  input         io_value_out_0_5_ready,
  output        io_value_out_0_5_valid,
  output [31:0] io_value_out_0_5_bits,
  input         io_value_out_0_6_ready,
  output        io_value_out_0_6_valid,
  output [31:0] io_value_out_0_6_bits,
  input         io_value_out_0_7_ready,
  output        io_value_out_0_7_valid,
  output [31:0] io_value_out_0_7_bits,
  input         io_value_out_0_8_ready,
  output        io_value_out_0_8_valid,
  output [31:0] io_value_out_0_8_bits,
  input         io_value_out_0_9_ready,
  output        io_value_out_0_9_valid,
  output [31:0] io_value_out_0_9_bits,
  input         io_value_out_0_10_ready,
  output        io_value_out_0_10_valid,
  output [31:0] io_value_out_0_10_bits,
  input         io_value_out_0_11_ready,
  output        io_value_out_0_11_valid,
  output [31:0] io_value_out_0_11_bits,
  input         io_value_out_0_12_ready,
  output        io_value_out_0_12_valid,
  output [31:0] io_value_out_0_12_bits,
  input         io_value_out_0_13_ready,
  output        io_value_out_0_13_valid,
  output [31:0] io_value_out_0_13_bits,
  input         io_value_out_0_14_ready,
  output        io_value_out_0_14_valid,
  output [31:0] io_value_out_0_14_bits,
  input         io_value_out_0_15_ready,
  output        io_value_out_0_15_valid,
  output [31:0] io_value_out_0_15_bits,
  input         io_value_out_1_0_ready,
  output        io_value_out_1_0_valid,
  output [31:0] io_value_out_1_0_bits,
  input         io_value_out_1_1_ready,
  output        io_value_out_1_1_valid,
  output [31:0] io_value_out_1_1_bits,
  input         io_value_out_1_2_ready,
  output        io_value_out_1_2_valid,
  output [31:0] io_value_out_1_2_bits,
  input         io_value_out_1_3_ready,
  output        io_value_out_1_3_valid,
  output [31:0] io_value_out_1_3_bits,
  input         io_value_out_1_4_ready,
  output        io_value_out_1_4_valid,
  output [31:0] io_value_out_1_4_bits,
  input         io_value_out_1_5_ready,
  output        io_value_out_1_5_valid,
  output [31:0] io_value_out_1_5_bits,
  input         io_value_out_1_6_ready,
  output        io_value_out_1_6_valid,
  output [31:0] io_value_out_1_6_bits,
  input         io_value_out_1_7_ready,
  output        io_value_out_1_7_valid,
  output [31:0] io_value_out_1_7_bits,
  input         io_value_out_1_8_ready,
  output        io_value_out_1_8_valid,
  output [31:0] io_value_out_1_8_bits,
  input         io_value_out_1_9_ready,
  output        io_value_out_1_9_valid,
  output [31:0] io_value_out_1_9_bits,
  input         io_value_out_1_10_ready,
  output        io_value_out_1_10_valid,
  output [31:0] io_value_out_1_10_bits,
  input         io_value_out_1_11_ready,
  output        io_value_out_1_11_valid,
  output [31:0] io_value_out_1_11_bits,
  input         io_value_out_1_12_ready,
  output        io_value_out_1_12_valid,
  output [31:0] io_value_out_1_12_bits,
  input         io_value_out_1_13_ready,
  output        io_value_out_1_13_valid,
  output [31:0] io_value_out_1_13_bits,
  input         io_value_out_1_14_ready,
  output        io_value_out_1_14_valid,
  output [31:0] io_value_out_1_14_bits,
  input         io_value_out_1_15_ready,
  output        io_value_out_1_15_valid,
  output [31:0] io_value_out_1_15_bits,
  input         io_value_out_2_0_ready,
  output        io_value_out_2_0_valid,
  output [31:0] io_value_out_2_0_bits,
  input         io_value_out_2_1_ready,
  output        io_value_out_2_1_valid,
  output [31:0] io_value_out_2_1_bits,
  input         io_value_out_2_2_ready,
  output        io_value_out_2_2_valid,
  output [31:0] io_value_out_2_2_bits,
  input         io_value_out_2_3_ready,
  output        io_value_out_2_3_valid,
  output [31:0] io_value_out_2_3_bits,
  input         io_value_out_2_4_ready,
  output        io_value_out_2_4_valid,
  output [31:0] io_value_out_2_4_bits,
  input         io_value_out_2_5_ready,
  output        io_value_out_2_5_valid,
  output [31:0] io_value_out_2_5_bits,
  input         io_value_out_2_6_ready,
  output        io_value_out_2_6_valid,
  output [31:0] io_value_out_2_6_bits,
  input         io_value_out_2_7_ready,
  output        io_value_out_2_7_valid,
  output [31:0] io_value_out_2_7_bits,
  input         io_value_out_2_8_ready,
  output        io_value_out_2_8_valid,
  output [31:0] io_value_out_2_8_bits,
  input         io_value_out_2_9_ready,
  output        io_value_out_2_9_valid,
  output [31:0] io_value_out_2_9_bits,
  input         io_value_out_2_10_ready,
  output        io_value_out_2_10_valid,
  output [31:0] io_value_out_2_10_bits,
  input         io_value_out_2_11_ready,
  output        io_value_out_2_11_valid,
  output [31:0] io_value_out_2_11_bits,
  input         io_value_out_2_12_ready,
  output        io_value_out_2_12_valid,
  output [31:0] io_value_out_2_12_bits,
  input         io_value_out_2_13_ready,
  output        io_value_out_2_13_valid,
  output [31:0] io_value_out_2_13_bits,
  input         io_value_out_2_14_ready,
  output        io_value_out_2_14_valid,
  output [31:0] io_value_out_2_14_bits,
  input         io_value_out_2_15_ready,
  output        io_value_out_2_15_valid,
  output [31:0] io_value_out_2_15_bits,
  input         io_value_out_3_0_ready,
  output        io_value_out_3_0_valid,
  output [31:0] io_value_out_3_0_bits,
  input         io_value_out_3_1_ready,
  output        io_value_out_3_1_valid,
  output [31:0] io_value_out_3_1_bits,
  input         io_value_out_3_2_ready,
  output        io_value_out_3_2_valid,
  output [31:0] io_value_out_3_2_bits,
  input         io_value_out_3_3_ready,
  output        io_value_out_3_3_valid,
  output [31:0] io_value_out_3_3_bits,
  input         io_value_out_3_4_ready,
  output        io_value_out_3_4_valid,
  output [31:0] io_value_out_3_4_bits,
  input         io_value_out_3_5_ready,
  output        io_value_out_3_5_valid,
  output [31:0] io_value_out_3_5_bits,
  input         io_value_out_3_6_ready,
  output        io_value_out_3_6_valid,
  output [31:0] io_value_out_3_6_bits,
  input         io_value_out_3_7_ready,
  output        io_value_out_3_7_valid,
  output [31:0] io_value_out_3_7_bits,
  input         io_value_out_3_8_ready,
  output        io_value_out_3_8_valid,
  output [31:0] io_value_out_3_8_bits,
  input         io_value_out_3_9_ready,
  output        io_value_out_3_9_valid,
  output [31:0] io_value_out_3_9_bits,
  input         io_value_out_3_10_ready,
  output        io_value_out_3_10_valid,
  output [31:0] io_value_out_3_10_bits,
  input         io_value_out_3_11_ready,
  output        io_value_out_3_11_valid,
  output [31:0] io_value_out_3_11_bits,
  input         io_value_out_3_12_ready,
  output        io_value_out_3_12_valid,
  output [31:0] io_value_out_3_12_bits,
  input         io_value_out_3_13_ready,
  output        io_value_out_3_13_valid,
  output [31:0] io_value_out_3_13_bits,
  input         io_value_out_3_14_ready,
  output        io_value_out_3_14_valid,
  output [31:0] io_value_out_3_14_bits,
  input         io_value_out_3_15_ready,
  output        io_value_out_3_15_valid,
  output [31:0] io_value_out_3_15_bits,
  input         io_value_out_4_0_ready,
  output        io_value_out_4_0_valid,
  output [31:0] io_value_out_4_0_bits,
  input         io_value_out_4_1_ready,
  output        io_value_out_4_1_valid,
  output [31:0] io_value_out_4_1_bits,
  input         io_value_out_4_2_ready,
  output        io_value_out_4_2_valid,
  output [31:0] io_value_out_4_2_bits,
  input         io_value_out_4_3_ready,
  output        io_value_out_4_3_valid,
  output [31:0] io_value_out_4_3_bits,
  input         io_value_out_4_4_ready,
  output        io_value_out_4_4_valid,
  output [31:0] io_value_out_4_4_bits,
  input         io_value_out_4_5_ready,
  output        io_value_out_4_5_valid,
  output [31:0] io_value_out_4_5_bits,
  input         io_value_out_4_6_ready,
  output        io_value_out_4_6_valid,
  output [31:0] io_value_out_4_6_bits,
  input         io_value_out_4_7_ready,
  output        io_value_out_4_7_valid,
  output [31:0] io_value_out_4_7_bits,
  input         io_value_out_4_8_ready,
  output        io_value_out_4_8_valid,
  output [31:0] io_value_out_4_8_bits,
  input         io_value_out_4_9_ready,
  output        io_value_out_4_9_valid,
  output [31:0] io_value_out_4_9_bits,
  input         io_value_out_4_10_ready,
  output        io_value_out_4_10_valid,
  output [31:0] io_value_out_4_10_bits,
  input         io_value_out_4_11_ready,
  output        io_value_out_4_11_valid,
  output [31:0] io_value_out_4_11_bits,
  input         io_value_out_4_12_ready,
  output        io_value_out_4_12_valid,
  output [31:0] io_value_out_4_12_bits,
  input         io_value_out_4_13_ready,
  output        io_value_out_4_13_valid,
  output [31:0] io_value_out_4_13_bits,
  input         io_value_out_4_14_ready,
  output        io_value_out_4_14_valid,
  output [31:0] io_value_out_4_14_bits,
  input         io_value_out_4_15_ready,
  output        io_value_out_4_15_valid,
  output [31:0] io_value_out_4_15_bits,
  input         io_value_out_5_0_ready,
  output        io_value_out_5_0_valid,
  output [31:0] io_value_out_5_0_bits,
  input         io_value_out_5_1_ready,
  output        io_value_out_5_1_valid,
  output [31:0] io_value_out_5_1_bits,
  input         io_value_out_5_2_ready,
  output        io_value_out_5_2_valid,
  output [31:0] io_value_out_5_2_bits,
  input         io_value_out_5_3_ready,
  output        io_value_out_5_3_valid,
  output [31:0] io_value_out_5_3_bits,
  input         io_value_out_5_4_ready,
  output        io_value_out_5_4_valid,
  output [31:0] io_value_out_5_4_bits,
  input         io_value_out_5_5_ready,
  output        io_value_out_5_5_valid,
  output [31:0] io_value_out_5_5_bits,
  input         io_value_out_5_6_ready,
  output        io_value_out_5_6_valid,
  output [31:0] io_value_out_5_6_bits,
  input         io_value_out_5_7_ready,
  output        io_value_out_5_7_valid,
  output [31:0] io_value_out_5_7_bits,
  input         io_value_out_5_8_ready,
  output        io_value_out_5_8_valid,
  output [31:0] io_value_out_5_8_bits,
  input         io_value_out_5_9_ready,
  output        io_value_out_5_9_valid,
  output [31:0] io_value_out_5_9_bits,
  input         io_value_out_5_10_ready,
  output        io_value_out_5_10_valid,
  output [31:0] io_value_out_5_10_bits,
  input         io_value_out_5_11_ready,
  output        io_value_out_5_11_valid,
  output [31:0] io_value_out_5_11_bits,
  input         io_value_out_5_12_ready,
  output        io_value_out_5_12_valid,
  output [31:0] io_value_out_5_12_bits,
  input         io_value_out_5_13_ready,
  output        io_value_out_5_13_valid,
  output [31:0] io_value_out_5_13_bits,
  input         io_value_out_5_14_ready,
  output        io_value_out_5_14_valid,
  output [31:0] io_value_out_5_14_bits,
  input         io_value_out_5_15_ready,
  output        io_value_out_5_15_valid,
  output [31:0] io_value_out_5_15_bits,
  input         io_value_out_6_0_ready,
  output        io_value_out_6_0_valid,
  output [31:0] io_value_out_6_0_bits,
  input         io_value_out_6_1_ready,
  output        io_value_out_6_1_valid,
  output [31:0] io_value_out_6_1_bits,
  input         io_value_out_6_2_ready,
  output        io_value_out_6_2_valid,
  output [31:0] io_value_out_6_2_bits,
  input         io_value_out_6_3_ready,
  output        io_value_out_6_3_valid,
  output [31:0] io_value_out_6_3_bits,
  input         io_value_out_6_4_ready,
  output        io_value_out_6_4_valid,
  output [31:0] io_value_out_6_4_bits,
  input         io_value_out_6_5_ready,
  output        io_value_out_6_5_valid,
  output [31:0] io_value_out_6_5_bits,
  input         io_value_out_6_6_ready,
  output        io_value_out_6_6_valid,
  output [31:0] io_value_out_6_6_bits,
  input         io_value_out_6_7_ready,
  output        io_value_out_6_7_valid,
  output [31:0] io_value_out_6_7_bits,
  input         io_value_out_6_8_ready,
  output        io_value_out_6_8_valid,
  output [31:0] io_value_out_6_8_bits,
  input         io_value_out_6_9_ready,
  output        io_value_out_6_9_valid,
  output [31:0] io_value_out_6_9_bits,
  input         io_value_out_6_10_ready,
  output        io_value_out_6_10_valid,
  output [31:0] io_value_out_6_10_bits,
  input         io_value_out_6_11_ready,
  output        io_value_out_6_11_valid,
  output [31:0] io_value_out_6_11_bits,
  input         io_value_out_6_12_ready,
  output        io_value_out_6_12_valid,
  output [31:0] io_value_out_6_12_bits,
  input         io_value_out_6_13_ready,
  output        io_value_out_6_13_valid,
  output [31:0] io_value_out_6_13_bits,
  input         io_value_out_6_14_ready,
  output        io_value_out_6_14_valid,
  output [31:0] io_value_out_6_14_bits,
  input         io_value_out_6_15_ready,
  output        io_value_out_6_15_valid,
  output [31:0] io_value_out_6_15_bits,
  input         io_value_out_7_0_ready,
  output        io_value_out_7_0_valid,
  output [31:0] io_value_out_7_0_bits,
  input         io_value_out_7_1_ready,
  output        io_value_out_7_1_valid,
  output [31:0] io_value_out_7_1_bits,
  input         io_value_out_7_2_ready,
  output        io_value_out_7_2_valid,
  output [31:0] io_value_out_7_2_bits,
  input         io_value_out_7_3_ready,
  output        io_value_out_7_3_valid,
  output [31:0] io_value_out_7_3_bits,
  input         io_value_out_7_4_ready,
  output        io_value_out_7_4_valid,
  output [31:0] io_value_out_7_4_bits,
  input         io_value_out_7_5_ready,
  output        io_value_out_7_5_valid,
  output [31:0] io_value_out_7_5_bits,
  input         io_value_out_7_6_ready,
  output        io_value_out_7_6_valid,
  output [31:0] io_value_out_7_6_bits,
  input         io_value_out_7_7_ready,
  output        io_value_out_7_7_valid,
  output [31:0] io_value_out_7_7_bits,
  input         io_value_out_7_8_ready,
  output        io_value_out_7_8_valid,
  output [31:0] io_value_out_7_8_bits,
  input         io_value_out_7_9_ready,
  output        io_value_out_7_9_valid,
  output [31:0] io_value_out_7_9_bits,
  input         io_value_out_7_10_ready,
  output        io_value_out_7_10_valid,
  output [31:0] io_value_out_7_10_bits,
  input         io_value_out_7_11_ready,
  output        io_value_out_7_11_valid,
  output [31:0] io_value_out_7_11_bits,
  input         io_value_out_7_12_ready,
  output        io_value_out_7_12_valid,
  output [31:0] io_value_out_7_12_bits,
  input         io_value_out_7_13_ready,
  output        io_value_out_7_13_valid,
  output [31:0] io_value_out_7_13_bits,
  input         io_value_out_7_14_ready,
  output        io_value_out_7_14_valid,
  output [31:0] io_value_out_7_14_bits,
  input         io_value_out_7_15_ready,
  output        io_value_out_7_15_valid,
  output [31:0] io_value_out_7_15_bits,
  input         io_value_out_8_0_ready,
  output        io_value_out_8_0_valid,
  output [31:0] io_value_out_8_0_bits,
  input         io_value_out_8_1_ready,
  output        io_value_out_8_1_valid,
  output [31:0] io_value_out_8_1_bits,
  input         io_value_out_8_2_ready,
  output        io_value_out_8_2_valid,
  output [31:0] io_value_out_8_2_bits,
  input         io_value_out_8_3_ready,
  output        io_value_out_8_3_valid,
  output [31:0] io_value_out_8_3_bits,
  input         io_value_out_8_4_ready,
  output        io_value_out_8_4_valid,
  output [31:0] io_value_out_8_4_bits,
  input         io_value_out_8_5_ready,
  output        io_value_out_8_5_valid,
  output [31:0] io_value_out_8_5_bits,
  input         io_value_out_8_6_ready,
  output        io_value_out_8_6_valid,
  output [31:0] io_value_out_8_6_bits,
  input         io_value_out_8_7_ready,
  output        io_value_out_8_7_valid,
  output [31:0] io_value_out_8_7_bits,
  input         io_value_out_8_8_ready,
  output        io_value_out_8_8_valid,
  output [31:0] io_value_out_8_8_bits,
  input         io_value_out_8_9_ready,
  output        io_value_out_8_9_valid,
  output [31:0] io_value_out_8_9_bits,
  input         io_value_out_8_10_ready,
  output        io_value_out_8_10_valid,
  output [31:0] io_value_out_8_10_bits,
  input         io_value_out_8_11_ready,
  output        io_value_out_8_11_valid,
  output [31:0] io_value_out_8_11_bits,
  input         io_value_out_8_12_ready,
  output        io_value_out_8_12_valid,
  output [31:0] io_value_out_8_12_bits,
  input         io_value_out_8_13_ready,
  output        io_value_out_8_13_valid,
  output [31:0] io_value_out_8_13_bits,
  input         io_value_out_8_14_ready,
  output        io_value_out_8_14_valid,
  output [31:0] io_value_out_8_14_bits,
  input         io_value_out_8_15_ready,
  output        io_value_out_8_15_valid,
  output [31:0] io_value_out_8_15_bits,
  input         io_value_out_9_0_ready,
  output        io_value_out_9_0_valid,
  output [31:0] io_value_out_9_0_bits,
  input         io_value_out_9_1_ready,
  output        io_value_out_9_1_valid,
  output [31:0] io_value_out_9_1_bits,
  input         io_value_out_9_2_ready,
  output        io_value_out_9_2_valid,
  output [31:0] io_value_out_9_2_bits,
  input         io_value_out_9_3_ready,
  output        io_value_out_9_3_valid,
  output [31:0] io_value_out_9_3_bits,
  input         io_value_out_9_4_ready,
  output        io_value_out_9_4_valid,
  output [31:0] io_value_out_9_4_bits,
  input         io_value_out_9_5_ready,
  output        io_value_out_9_5_valid,
  output [31:0] io_value_out_9_5_bits,
  input         io_value_out_9_6_ready,
  output        io_value_out_9_6_valid,
  output [31:0] io_value_out_9_6_bits,
  input         io_value_out_9_7_ready,
  output        io_value_out_9_7_valid,
  output [31:0] io_value_out_9_7_bits,
  input         io_value_out_9_8_ready,
  output        io_value_out_9_8_valid,
  output [31:0] io_value_out_9_8_bits,
  input         io_value_out_9_9_ready,
  output        io_value_out_9_9_valid,
  output [31:0] io_value_out_9_9_bits,
  input         io_value_out_9_10_ready,
  output        io_value_out_9_10_valid,
  output [31:0] io_value_out_9_10_bits,
  input         io_value_out_9_11_ready,
  output        io_value_out_9_11_valid,
  output [31:0] io_value_out_9_11_bits,
  input         io_value_out_9_12_ready,
  output        io_value_out_9_12_valid,
  output [31:0] io_value_out_9_12_bits,
  input         io_value_out_9_13_ready,
  output        io_value_out_9_13_valid,
  output [31:0] io_value_out_9_13_bits,
  input         io_value_out_9_14_ready,
  output        io_value_out_9_14_valid,
  output [31:0] io_value_out_9_14_bits,
  input         io_value_out_9_15_ready,
  output        io_value_out_9_15_valid,
  output [31:0] io_value_out_9_15_bits,
  input         io_value_out_10_0_ready,
  output        io_value_out_10_0_valid,
  output [31:0] io_value_out_10_0_bits,
  input         io_value_out_10_1_ready,
  output        io_value_out_10_1_valid,
  output [31:0] io_value_out_10_1_bits,
  input         io_value_out_10_2_ready,
  output        io_value_out_10_2_valid,
  output [31:0] io_value_out_10_2_bits,
  input         io_value_out_10_3_ready,
  output        io_value_out_10_3_valid,
  output [31:0] io_value_out_10_3_bits,
  input         io_value_out_10_4_ready,
  output        io_value_out_10_4_valid,
  output [31:0] io_value_out_10_4_bits,
  input         io_value_out_10_5_ready,
  output        io_value_out_10_5_valid,
  output [31:0] io_value_out_10_5_bits,
  input         io_value_out_10_6_ready,
  output        io_value_out_10_6_valid,
  output [31:0] io_value_out_10_6_bits,
  input         io_value_out_10_7_ready,
  output        io_value_out_10_7_valid,
  output [31:0] io_value_out_10_7_bits,
  input         io_value_out_10_8_ready,
  output        io_value_out_10_8_valid,
  output [31:0] io_value_out_10_8_bits,
  input         io_value_out_10_9_ready,
  output        io_value_out_10_9_valid,
  output [31:0] io_value_out_10_9_bits,
  input         io_value_out_10_10_ready,
  output        io_value_out_10_10_valid,
  output [31:0] io_value_out_10_10_bits,
  input         io_value_out_10_11_ready,
  output        io_value_out_10_11_valid,
  output [31:0] io_value_out_10_11_bits,
  input         io_value_out_10_12_ready,
  output        io_value_out_10_12_valid,
  output [31:0] io_value_out_10_12_bits,
  input         io_value_out_10_13_ready,
  output        io_value_out_10_13_valid,
  output [31:0] io_value_out_10_13_bits,
  input         io_value_out_10_14_ready,
  output        io_value_out_10_14_valid,
  output [31:0] io_value_out_10_14_bits,
  input         io_value_out_10_15_ready,
  output        io_value_out_10_15_valid,
  output [31:0] io_value_out_10_15_bits,
  input         io_value_out_11_0_ready,
  output        io_value_out_11_0_valid,
  output [31:0] io_value_out_11_0_bits,
  input         io_value_out_11_1_ready,
  output        io_value_out_11_1_valid,
  output [31:0] io_value_out_11_1_bits,
  input         io_value_out_11_2_ready,
  output        io_value_out_11_2_valid,
  output [31:0] io_value_out_11_2_bits,
  input         io_value_out_11_3_ready,
  output        io_value_out_11_3_valid,
  output [31:0] io_value_out_11_3_bits,
  input         io_value_out_11_4_ready,
  output        io_value_out_11_4_valid,
  output [31:0] io_value_out_11_4_bits,
  input         io_value_out_11_5_ready,
  output        io_value_out_11_5_valid,
  output [31:0] io_value_out_11_5_bits,
  input         io_value_out_11_6_ready,
  output        io_value_out_11_6_valid,
  output [31:0] io_value_out_11_6_bits,
  input         io_value_out_11_7_ready,
  output        io_value_out_11_7_valid,
  output [31:0] io_value_out_11_7_bits,
  input         io_value_out_11_8_ready,
  output        io_value_out_11_8_valid,
  output [31:0] io_value_out_11_8_bits,
  input         io_value_out_11_9_ready,
  output        io_value_out_11_9_valid,
  output [31:0] io_value_out_11_9_bits,
  input         io_value_out_11_10_ready,
  output        io_value_out_11_10_valid,
  output [31:0] io_value_out_11_10_bits,
  input         io_value_out_11_11_ready,
  output        io_value_out_11_11_valid,
  output [31:0] io_value_out_11_11_bits,
  input         io_value_out_11_12_ready,
  output        io_value_out_11_12_valid,
  output [31:0] io_value_out_11_12_bits,
  input         io_value_out_11_13_ready,
  output        io_value_out_11_13_valid,
  output [31:0] io_value_out_11_13_bits,
  input         io_value_out_11_14_ready,
  output        io_value_out_11_14_valid,
  output [31:0] io_value_out_11_14_bits,
  input         io_value_out_11_15_ready,
  output        io_value_out_11_15_valid,
  output [31:0] io_value_out_11_15_bits,
  input         io_value_out_12_0_ready,
  output        io_value_out_12_0_valid,
  output [31:0] io_value_out_12_0_bits,
  input         io_value_out_12_1_ready,
  output        io_value_out_12_1_valid,
  output [31:0] io_value_out_12_1_bits,
  input         io_value_out_12_2_ready,
  output        io_value_out_12_2_valid,
  output [31:0] io_value_out_12_2_bits,
  input         io_value_out_12_3_ready,
  output        io_value_out_12_3_valid,
  output [31:0] io_value_out_12_3_bits,
  input         io_value_out_12_4_ready,
  output        io_value_out_12_4_valid,
  output [31:0] io_value_out_12_4_bits,
  input         io_value_out_12_5_ready,
  output        io_value_out_12_5_valid,
  output [31:0] io_value_out_12_5_bits,
  input         io_value_out_12_6_ready,
  output        io_value_out_12_6_valid,
  output [31:0] io_value_out_12_6_bits,
  input         io_value_out_12_7_ready,
  output        io_value_out_12_7_valid,
  output [31:0] io_value_out_12_7_bits,
  input         io_value_out_12_8_ready,
  output        io_value_out_12_8_valid,
  output [31:0] io_value_out_12_8_bits,
  input         io_value_out_12_9_ready,
  output        io_value_out_12_9_valid,
  output [31:0] io_value_out_12_9_bits,
  input         io_value_out_12_10_ready,
  output        io_value_out_12_10_valid,
  output [31:0] io_value_out_12_10_bits,
  input         io_value_out_12_11_ready,
  output        io_value_out_12_11_valid,
  output [31:0] io_value_out_12_11_bits,
  input         io_value_out_12_12_ready,
  output        io_value_out_12_12_valid,
  output [31:0] io_value_out_12_12_bits,
  input         io_value_out_12_13_ready,
  output        io_value_out_12_13_valid,
  output [31:0] io_value_out_12_13_bits,
  input         io_value_out_12_14_ready,
  output        io_value_out_12_14_valid,
  output [31:0] io_value_out_12_14_bits,
  input         io_value_out_12_15_ready,
  output        io_value_out_12_15_valid,
  output [31:0] io_value_out_12_15_bits,
  input         io_value_out_13_0_ready,
  output        io_value_out_13_0_valid,
  output [31:0] io_value_out_13_0_bits,
  input         io_value_out_13_1_ready,
  output        io_value_out_13_1_valid,
  output [31:0] io_value_out_13_1_bits,
  input         io_value_out_13_2_ready,
  output        io_value_out_13_2_valid,
  output [31:0] io_value_out_13_2_bits,
  input         io_value_out_13_3_ready,
  output        io_value_out_13_3_valid,
  output [31:0] io_value_out_13_3_bits,
  input         io_value_out_13_4_ready,
  output        io_value_out_13_4_valid,
  output [31:0] io_value_out_13_4_bits,
  input         io_value_out_13_5_ready,
  output        io_value_out_13_5_valid,
  output [31:0] io_value_out_13_5_bits,
  input         io_value_out_13_6_ready,
  output        io_value_out_13_6_valid,
  output [31:0] io_value_out_13_6_bits,
  input         io_value_out_13_7_ready,
  output        io_value_out_13_7_valid,
  output [31:0] io_value_out_13_7_bits,
  input         io_value_out_13_8_ready,
  output        io_value_out_13_8_valid,
  output [31:0] io_value_out_13_8_bits,
  input         io_value_out_13_9_ready,
  output        io_value_out_13_9_valid,
  output [31:0] io_value_out_13_9_bits,
  input         io_value_out_13_10_ready,
  output        io_value_out_13_10_valid,
  output [31:0] io_value_out_13_10_bits,
  input         io_value_out_13_11_ready,
  output        io_value_out_13_11_valid,
  output [31:0] io_value_out_13_11_bits,
  input         io_value_out_13_12_ready,
  output        io_value_out_13_12_valid,
  output [31:0] io_value_out_13_12_bits,
  input         io_value_out_13_13_ready,
  output        io_value_out_13_13_valid,
  output [31:0] io_value_out_13_13_bits,
  input         io_value_out_13_14_ready,
  output        io_value_out_13_14_valid,
  output [31:0] io_value_out_13_14_bits,
  input         io_value_out_13_15_ready,
  output        io_value_out_13_15_valid,
  output [31:0] io_value_out_13_15_bits,
  input         io_value_out_14_0_ready,
  output        io_value_out_14_0_valid,
  output [31:0] io_value_out_14_0_bits,
  input         io_value_out_14_1_ready,
  output        io_value_out_14_1_valid,
  output [31:0] io_value_out_14_1_bits,
  input         io_value_out_14_2_ready,
  output        io_value_out_14_2_valid,
  output [31:0] io_value_out_14_2_bits,
  input         io_value_out_14_3_ready,
  output        io_value_out_14_3_valid,
  output [31:0] io_value_out_14_3_bits,
  input         io_value_out_14_4_ready,
  output        io_value_out_14_4_valid,
  output [31:0] io_value_out_14_4_bits,
  input         io_value_out_14_5_ready,
  output        io_value_out_14_5_valid,
  output [31:0] io_value_out_14_5_bits,
  input         io_value_out_14_6_ready,
  output        io_value_out_14_6_valid,
  output [31:0] io_value_out_14_6_bits,
  input         io_value_out_14_7_ready,
  output        io_value_out_14_7_valid,
  output [31:0] io_value_out_14_7_bits,
  input         io_value_out_14_8_ready,
  output        io_value_out_14_8_valid,
  output [31:0] io_value_out_14_8_bits,
  input         io_value_out_14_9_ready,
  output        io_value_out_14_9_valid,
  output [31:0] io_value_out_14_9_bits,
  input         io_value_out_14_10_ready,
  output        io_value_out_14_10_valid,
  output [31:0] io_value_out_14_10_bits,
  input         io_value_out_14_11_ready,
  output        io_value_out_14_11_valid,
  output [31:0] io_value_out_14_11_bits,
  input         io_value_out_14_12_ready,
  output        io_value_out_14_12_valid,
  output [31:0] io_value_out_14_12_bits,
  input         io_value_out_14_13_ready,
  output        io_value_out_14_13_valid,
  output [31:0] io_value_out_14_13_bits,
  input         io_value_out_14_14_ready,
  output        io_value_out_14_14_valid,
  output [31:0] io_value_out_14_14_bits,
  input         io_value_out_14_15_ready,
  output        io_value_out_14_15_valid,
  output [31:0] io_value_out_14_15_bits,
  input         io_value_out_15_0_ready,
  output        io_value_out_15_0_valid,
  output [31:0] io_value_out_15_0_bits,
  input         io_value_out_15_1_ready,
  output        io_value_out_15_1_valid,
  output [31:0] io_value_out_15_1_bits,
  input         io_value_out_15_2_ready,
  output        io_value_out_15_2_valid,
  output [31:0] io_value_out_15_2_bits,
  input         io_value_out_15_3_ready,
  output        io_value_out_15_3_valid,
  output [31:0] io_value_out_15_3_bits,
  input         io_value_out_15_4_ready,
  output        io_value_out_15_4_valid,
  output [31:0] io_value_out_15_4_bits,
  input         io_value_out_15_5_ready,
  output        io_value_out_15_5_valid,
  output [31:0] io_value_out_15_5_bits,
  input         io_value_out_15_6_ready,
  output        io_value_out_15_6_valid,
  output [31:0] io_value_out_15_6_bits,
  input         io_value_out_15_7_ready,
  output        io_value_out_15_7_valid,
  output [31:0] io_value_out_15_7_bits,
  input         io_value_out_15_8_ready,
  output        io_value_out_15_8_valid,
  output [31:0] io_value_out_15_8_bits,
  input         io_value_out_15_9_ready,
  output        io_value_out_15_9_valid,
  output [31:0] io_value_out_15_9_bits,
  input         io_value_out_15_10_ready,
  output        io_value_out_15_10_valid,
  output [31:0] io_value_out_15_10_bits,
  input         io_value_out_15_11_ready,
  output        io_value_out_15_11_valid,
  output [31:0] io_value_out_15_11_bits,
  input         io_value_out_15_12_ready,
  output        io_value_out_15_12_valid,
  output [31:0] io_value_out_15_12_bits,
  input         io_value_out_15_13_ready,
  output        io_value_out_15_13_valid,
  output [31:0] io_value_out_15_13_bits,
  input         io_value_out_15_14_ready,
  output        io_value_out_15_14_valid,
  output [31:0] io_value_out_15_14_bits,
  input         io_value_out_15_15_ready,
  output        io_value_out_15_15_valid,
  output [31:0] io_value_out_15_15_bits
);
  wire  cols_0_0_clock; // @[Stab.scala 85:60]
  wire  cols_0_0_reset; // @[Stab.scala 85:60]
  wire  cols_0_0_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_0_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_0_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_0_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_0_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_0_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_0_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_0_0_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_0_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_0_0_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_0_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_0_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_0_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_0_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_0_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_0_clock; // @[Stab.scala 85:60]
  wire  cols_1_0_reset; // @[Stab.scala 85:60]
  wire  cols_1_0_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_0_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_0_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_0_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_0_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_0_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_0_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_1_0_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_0_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_1_0_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_0_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_0_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_0_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_0_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_0_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_0_clock; // @[Stab.scala 85:60]
  wire  cols_2_0_reset; // @[Stab.scala 85:60]
  wire  cols_2_0_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_0_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_0_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_0_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_0_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_0_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_0_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_2_0_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_0_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_2_0_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_0_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_0_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_0_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_0_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_0_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_0_clock; // @[Stab.scala 85:60]
  wire  cols_3_0_reset; // @[Stab.scala 85:60]
  wire  cols_3_0_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_0_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_0_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_0_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_0_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_0_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_0_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_3_0_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_0_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_3_0_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_0_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_0_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_0_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_0_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_0_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_0_clock; // @[Stab.scala 85:60]
  wire  cols_4_0_reset; // @[Stab.scala 85:60]
  wire  cols_4_0_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_0_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_0_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_0_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_0_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_0_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_0_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_4_0_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_0_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_4_0_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_0_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_0_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_0_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_0_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_0_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_0_clock; // @[Stab.scala 85:60]
  wire  cols_5_0_reset; // @[Stab.scala 85:60]
  wire  cols_5_0_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_0_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_0_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_0_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_0_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_0_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_0_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_5_0_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_0_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_5_0_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_0_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_0_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_0_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_0_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_0_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_0_clock; // @[Stab.scala 85:60]
  wire  cols_6_0_reset; // @[Stab.scala 85:60]
  wire  cols_6_0_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_0_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_0_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_0_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_0_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_0_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_0_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_6_0_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_0_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_6_0_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_0_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_0_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_0_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_0_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_0_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_0_clock; // @[Stab.scala 85:60]
  wire  cols_7_0_reset; // @[Stab.scala 85:60]
  wire  cols_7_0_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_0_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_0_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_0_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_0_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_0_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_0_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_7_0_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_0_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_7_0_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_0_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_0_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_0_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_0_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_0_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_0_clock; // @[Stab.scala 85:60]
  wire  cols_8_0_reset; // @[Stab.scala 85:60]
  wire  cols_8_0_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_0_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_0_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_0_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_0_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_0_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_0_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_8_0_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_0_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_8_0_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_0_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_0_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_0_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_0_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_0_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_0_clock; // @[Stab.scala 85:60]
  wire  cols_9_0_reset; // @[Stab.scala 85:60]
  wire  cols_9_0_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_0_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_0_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_0_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_0_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_0_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_0_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_9_0_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_0_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_9_0_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_0_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_0_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_0_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_0_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_0_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_0_clock; // @[Stab.scala 85:60]
  wire  cols_10_0_reset; // @[Stab.scala 85:60]
  wire  cols_10_0_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_0_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_0_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_0_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_0_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_0_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_0_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_10_0_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_0_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_10_0_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_0_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_0_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_0_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_0_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_0_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_0_clock; // @[Stab.scala 85:60]
  wire  cols_11_0_reset; // @[Stab.scala 85:60]
  wire  cols_11_0_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_0_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_0_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_0_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_0_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_0_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_0_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_11_0_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_0_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_11_0_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_0_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_0_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_0_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_0_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_0_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_0_clock; // @[Stab.scala 85:60]
  wire  cols_12_0_reset; // @[Stab.scala 85:60]
  wire  cols_12_0_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_0_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_0_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_0_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_0_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_0_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_0_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_12_0_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_0_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_12_0_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_0_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_0_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_0_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_0_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_0_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_0_clock; // @[Stab.scala 85:60]
  wire  cols_13_0_reset; // @[Stab.scala 85:60]
  wire  cols_13_0_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_0_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_0_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_0_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_0_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_0_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_0_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_13_0_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_0_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_13_0_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_0_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_0_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_0_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_0_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_0_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_0_clock; // @[Stab.scala 85:60]
  wire  cols_14_0_reset; // @[Stab.scala 85:60]
  wire  cols_14_0_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_0_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_0_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_0_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_0_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_0_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_0_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_14_0_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_0_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_14_0_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_0_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_0_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_0_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_0_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_0_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_0_clock; // @[Stab.scala 85:60]
  wire  cols_15_0_reset; // @[Stab.scala 85:60]
  wire  cols_15_0_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_0_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_0_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_0_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_0_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_0_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_0_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_15_0_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_0_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_15_0_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_0_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_0_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_0_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_0_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_0_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_1_clock; // @[Stab.scala 85:60]
  wire  cols_0_1_reset; // @[Stab.scala 85:60]
  wire  cols_0_1_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_1_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_1_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_1_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_1_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_1_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_1_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_0_1_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_1_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_0_1_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_1_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_1_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_1_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_1_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_1_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_1_clock; // @[Stab.scala 85:60]
  wire  cols_1_1_reset; // @[Stab.scala 85:60]
  wire  cols_1_1_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_1_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_1_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_1_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_1_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_1_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_1_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_1_1_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_1_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_1_1_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_1_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_1_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_1_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_1_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_1_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_1_clock; // @[Stab.scala 85:60]
  wire  cols_2_1_reset; // @[Stab.scala 85:60]
  wire  cols_2_1_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_1_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_1_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_1_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_1_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_1_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_1_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_2_1_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_1_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_2_1_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_1_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_1_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_1_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_1_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_1_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_1_clock; // @[Stab.scala 85:60]
  wire  cols_3_1_reset; // @[Stab.scala 85:60]
  wire  cols_3_1_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_1_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_1_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_1_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_1_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_1_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_1_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_3_1_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_1_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_3_1_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_1_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_1_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_1_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_1_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_1_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_1_clock; // @[Stab.scala 85:60]
  wire  cols_4_1_reset; // @[Stab.scala 85:60]
  wire  cols_4_1_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_1_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_1_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_1_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_1_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_1_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_1_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_4_1_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_1_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_4_1_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_1_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_1_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_1_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_1_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_1_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_1_clock; // @[Stab.scala 85:60]
  wire  cols_5_1_reset; // @[Stab.scala 85:60]
  wire  cols_5_1_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_1_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_1_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_1_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_1_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_1_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_1_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_5_1_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_1_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_5_1_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_1_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_1_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_1_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_1_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_1_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_1_clock; // @[Stab.scala 85:60]
  wire  cols_6_1_reset; // @[Stab.scala 85:60]
  wire  cols_6_1_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_1_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_1_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_1_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_1_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_1_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_1_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_6_1_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_1_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_6_1_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_1_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_1_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_1_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_1_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_1_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_1_clock; // @[Stab.scala 85:60]
  wire  cols_7_1_reset; // @[Stab.scala 85:60]
  wire  cols_7_1_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_1_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_1_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_1_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_1_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_1_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_1_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_7_1_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_1_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_7_1_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_1_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_1_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_1_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_1_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_1_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_1_clock; // @[Stab.scala 85:60]
  wire  cols_8_1_reset; // @[Stab.scala 85:60]
  wire  cols_8_1_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_1_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_1_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_1_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_1_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_1_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_1_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_8_1_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_1_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_8_1_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_1_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_1_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_1_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_1_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_1_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_1_clock; // @[Stab.scala 85:60]
  wire  cols_9_1_reset; // @[Stab.scala 85:60]
  wire  cols_9_1_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_1_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_1_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_1_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_1_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_1_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_1_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_9_1_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_1_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_9_1_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_1_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_1_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_1_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_1_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_1_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_1_clock; // @[Stab.scala 85:60]
  wire  cols_10_1_reset; // @[Stab.scala 85:60]
  wire  cols_10_1_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_1_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_1_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_1_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_1_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_1_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_1_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_10_1_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_1_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_10_1_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_1_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_1_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_1_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_1_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_1_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_1_clock; // @[Stab.scala 85:60]
  wire  cols_11_1_reset; // @[Stab.scala 85:60]
  wire  cols_11_1_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_1_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_1_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_1_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_1_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_1_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_1_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_11_1_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_1_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_11_1_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_1_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_1_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_1_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_1_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_1_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_1_clock; // @[Stab.scala 85:60]
  wire  cols_12_1_reset; // @[Stab.scala 85:60]
  wire  cols_12_1_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_1_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_1_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_1_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_1_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_1_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_1_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_12_1_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_1_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_12_1_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_1_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_1_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_1_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_1_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_1_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_1_clock; // @[Stab.scala 85:60]
  wire  cols_13_1_reset; // @[Stab.scala 85:60]
  wire  cols_13_1_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_1_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_1_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_1_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_1_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_1_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_1_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_13_1_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_1_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_13_1_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_1_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_1_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_1_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_1_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_1_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_1_clock; // @[Stab.scala 85:60]
  wire  cols_14_1_reset; // @[Stab.scala 85:60]
  wire  cols_14_1_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_1_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_1_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_1_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_1_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_1_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_1_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_14_1_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_1_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_14_1_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_1_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_1_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_1_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_1_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_1_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_1_clock; // @[Stab.scala 85:60]
  wire  cols_15_1_reset; // @[Stab.scala 85:60]
  wire  cols_15_1_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_1_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_1_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_1_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_1_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_1_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_1_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_15_1_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_1_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_15_1_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_1_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_1_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_1_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_1_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_1_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_2_clock; // @[Stab.scala 85:60]
  wire  cols_0_2_reset; // @[Stab.scala 85:60]
  wire  cols_0_2_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_2_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_2_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_2_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_2_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_2_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_2_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_0_2_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_2_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_0_2_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_2_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_2_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_2_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_2_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_2_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_2_clock; // @[Stab.scala 85:60]
  wire  cols_1_2_reset; // @[Stab.scala 85:60]
  wire  cols_1_2_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_2_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_2_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_2_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_2_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_2_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_2_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_1_2_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_2_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_1_2_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_2_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_2_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_2_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_2_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_2_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_2_clock; // @[Stab.scala 85:60]
  wire  cols_2_2_reset; // @[Stab.scala 85:60]
  wire  cols_2_2_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_2_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_2_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_2_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_2_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_2_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_2_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_2_2_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_2_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_2_2_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_2_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_2_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_2_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_2_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_2_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_2_clock; // @[Stab.scala 85:60]
  wire  cols_3_2_reset; // @[Stab.scala 85:60]
  wire  cols_3_2_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_2_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_2_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_2_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_2_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_2_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_2_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_3_2_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_2_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_3_2_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_2_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_2_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_2_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_2_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_2_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_2_clock; // @[Stab.scala 85:60]
  wire  cols_4_2_reset; // @[Stab.scala 85:60]
  wire  cols_4_2_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_2_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_2_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_2_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_2_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_2_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_2_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_4_2_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_2_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_4_2_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_2_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_2_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_2_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_2_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_2_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_2_clock; // @[Stab.scala 85:60]
  wire  cols_5_2_reset; // @[Stab.scala 85:60]
  wire  cols_5_2_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_2_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_2_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_2_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_2_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_2_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_2_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_5_2_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_2_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_5_2_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_2_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_2_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_2_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_2_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_2_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_2_clock; // @[Stab.scala 85:60]
  wire  cols_6_2_reset; // @[Stab.scala 85:60]
  wire  cols_6_2_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_2_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_2_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_2_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_2_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_2_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_2_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_6_2_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_2_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_6_2_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_2_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_2_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_2_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_2_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_2_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_2_clock; // @[Stab.scala 85:60]
  wire  cols_7_2_reset; // @[Stab.scala 85:60]
  wire  cols_7_2_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_2_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_2_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_2_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_2_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_2_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_2_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_7_2_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_2_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_7_2_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_2_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_2_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_2_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_2_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_2_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_2_clock; // @[Stab.scala 85:60]
  wire  cols_8_2_reset; // @[Stab.scala 85:60]
  wire  cols_8_2_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_2_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_2_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_2_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_2_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_2_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_2_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_8_2_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_2_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_8_2_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_2_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_2_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_2_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_2_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_2_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_2_clock; // @[Stab.scala 85:60]
  wire  cols_9_2_reset; // @[Stab.scala 85:60]
  wire  cols_9_2_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_2_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_2_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_2_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_2_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_2_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_2_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_9_2_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_2_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_9_2_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_2_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_2_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_2_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_2_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_2_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_2_clock; // @[Stab.scala 85:60]
  wire  cols_10_2_reset; // @[Stab.scala 85:60]
  wire  cols_10_2_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_2_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_2_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_2_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_2_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_2_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_2_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_10_2_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_2_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_10_2_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_2_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_2_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_2_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_2_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_2_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_2_clock; // @[Stab.scala 85:60]
  wire  cols_11_2_reset; // @[Stab.scala 85:60]
  wire  cols_11_2_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_2_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_2_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_2_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_2_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_2_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_2_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_11_2_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_2_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_11_2_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_2_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_2_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_2_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_2_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_2_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_2_clock; // @[Stab.scala 85:60]
  wire  cols_12_2_reset; // @[Stab.scala 85:60]
  wire  cols_12_2_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_2_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_2_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_2_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_2_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_2_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_2_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_12_2_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_2_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_12_2_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_2_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_2_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_2_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_2_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_2_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_2_clock; // @[Stab.scala 85:60]
  wire  cols_13_2_reset; // @[Stab.scala 85:60]
  wire  cols_13_2_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_2_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_2_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_2_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_2_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_2_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_2_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_13_2_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_2_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_13_2_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_2_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_2_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_2_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_2_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_2_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_2_clock; // @[Stab.scala 85:60]
  wire  cols_14_2_reset; // @[Stab.scala 85:60]
  wire  cols_14_2_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_2_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_2_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_2_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_2_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_2_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_2_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_14_2_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_2_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_14_2_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_2_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_2_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_2_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_2_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_2_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_2_clock; // @[Stab.scala 85:60]
  wire  cols_15_2_reset; // @[Stab.scala 85:60]
  wire  cols_15_2_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_2_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_2_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_2_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_2_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_2_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_2_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_15_2_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_2_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_15_2_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_2_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_2_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_2_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_2_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_2_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_3_clock; // @[Stab.scala 85:60]
  wire  cols_0_3_reset; // @[Stab.scala 85:60]
  wire  cols_0_3_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_3_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_3_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_3_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_3_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_3_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_3_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_0_3_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_3_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_0_3_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_3_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_3_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_3_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_3_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_3_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_3_clock; // @[Stab.scala 85:60]
  wire  cols_1_3_reset; // @[Stab.scala 85:60]
  wire  cols_1_3_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_3_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_3_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_3_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_3_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_3_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_3_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_1_3_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_3_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_1_3_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_3_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_3_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_3_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_3_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_3_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_3_clock; // @[Stab.scala 85:60]
  wire  cols_2_3_reset; // @[Stab.scala 85:60]
  wire  cols_2_3_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_3_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_3_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_3_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_3_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_3_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_3_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_2_3_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_3_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_2_3_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_3_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_3_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_3_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_3_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_3_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_3_clock; // @[Stab.scala 85:60]
  wire  cols_3_3_reset; // @[Stab.scala 85:60]
  wire  cols_3_3_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_3_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_3_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_3_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_3_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_3_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_3_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_3_3_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_3_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_3_3_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_3_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_3_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_3_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_3_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_3_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_3_clock; // @[Stab.scala 85:60]
  wire  cols_4_3_reset; // @[Stab.scala 85:60]
  wire  cols_4_3_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_3_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_3_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_3_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_3_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_3_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_3_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_4_3_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_3_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_4_3_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_3_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_3_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_3_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_3_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_3_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_3_clock; // @[Stab.scala 85:60]
  wire  cols_5_3_reset; // @[Stab.scala 85:60]
  wire  cols_5_3_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_3_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_3_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_3_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_3_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_3_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_3_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_5_3_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_3_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_5_3_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_3_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_3_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_3_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_3_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_3_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_3_clock; // @[Stab.scala 85:60]
  wire  cols_6_3_reset; // @[Stab.scala 85:60]
  wire  cols_6_3_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_3_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_3_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_3_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_3_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_3_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_3_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_6_3_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_3_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_6_3_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_3_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_3_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_3_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_3_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_3_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_3_clock; // @[Stab.scala 85:60]
  wire  cols_7_3_reset; // @[Stab.scala 85:60]
  wire  cols_7_3_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_3_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_3_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_3_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_3_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_3_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_3_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_7_3_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_3_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_7_3_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_3_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_3_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_3_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_3_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_3_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_3_clock; // @[Stab.scala 85:60]
  wire  cols_8_3_reset; // @[Stab.scala 85:60]
  wire  cols_8_3_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_3_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_3_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_3_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_3_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_3_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_3_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_8_3_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_3_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_8_3_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_3_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_3_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_3_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_3_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_3_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_3_clock; // @[Stab.scala 85:60]
  wire  cols_9_3_reset; // @[Stab.scala 85:60]
  wire  cols_9_3_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_3_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_3_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_3_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_3_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_3_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_3_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_9_3_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_3_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_9_3_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_3_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_3_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_3_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_3_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_3_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_3_clock; // @[Stab.scala 85:60]
  wire  cols_10_3_reset; // @[Stab.scala 85:60]
  wire  cols_10_3_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_3_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_3_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_3_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_3_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_3_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_3_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_10_3_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_3_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_10_3_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_3_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_3_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_3_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_3_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_3_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_3_clock; // @[Stab.scala 85:60]
  wire  cols_11_3_reset; // @[Stab.scala 85:60]
  wire  cols_11_3_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_3_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_3_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_3_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_3_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_3_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_3_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_11_3_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_3_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_11_3_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_3_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_3_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_3_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_3_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_3_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_3_clock; // @[Stab.scala 85:60]
  wire  cols_12_3_reset; // @[Stab.scala 85:60]
  wire  cols_12_3_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_3_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_3_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_3_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_3_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_3_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_3_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_12_3_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_3_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_12_3_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_3_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_3_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_3_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_3_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_3_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_3_clock; // @[Stab.scala 85:60]
  wire  cols_13_3_reset; // @[Stab.scala 85:60]
  wire  cols_13_3_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_3_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_3_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_3_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_3_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_3_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_3_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_13_3_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_3_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_13_3_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_3_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_3_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_3_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_3_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_3_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_3_clock; // @[Stab.scala 85:60]
  wire  cols_14_3_reset; // @[Stab.scala 85:60]
  wire  cols_14_3_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_3_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_3_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_3_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_3_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_3_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_3_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_14_3_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_3_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_14_3_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_3_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_3_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_3_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_3_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_3_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_3_clock; // @[Stab.scala 85:60]
  wire  cols_15_3_reset; // @[Stab.scala 85:60]
  wire  cols_15_3_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_3_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_3_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_3_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_3_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_3_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_3_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_15_3_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_3_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_15_3_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_3_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_3_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_3_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_3_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_3_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_4_clock; // @[Stab.scala 85:60]
  wire  cols_0_4_reset; // @[Stab.scala 85:60]
  wire  cols_0_4_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_4_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_4_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_4_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_4_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_4_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_4_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_0_4_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_4_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_0_4_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_4_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_4_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_4_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_4_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_4_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_4_clock; // @[Stab.scala 85:60]
  wire  cols_1_4_reset; // @[Stab.scala 85:60]
  wire  cols_1_4_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_4_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_4_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_4_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_4_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_4_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_4_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_1_4_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_4_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_1_4_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_4_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_4_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_4_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_4_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_4_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_4_clock; // @[Stab.scala 85:60]
  wire  cols_2_4_reset; // @[Stab.scala 85:60]
  wire  cols_2_4_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_4_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_4_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_4_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_4_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_4_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_4_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_2_4_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_4_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_2_4_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_4_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_4_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_4_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_4_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_4_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_4_clock; // @[Stab.scala 85:60]
  wire  cols_3_4_reset; // @[Stab.scala 85:60]
  wire  cols_3_4_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_4_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_4_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_4_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_4_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_4_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_4_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_3_4_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_4_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_3_4_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_4_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_4_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_4_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_4_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_4_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_4_clock; // @[Stab.scala 85:60]
  wire  cols_4_4_reset; // @[Stab.scala 85:60]
  wire  cols_4_4_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_4_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_4_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_4_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_4_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_4_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_4_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_4_4_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_4_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_4_4_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_4_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_4_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_4_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_4_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_4_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_4_clock; // @[Stab.scala 85:60]
  wire  cols_5_4_reset; // @[Stab.scala 85:60]
  wire  cols_5_4_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_4_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_4_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_4_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_4_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_4_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_4_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_5_4_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_4_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_5_4_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_4_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_4_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_4_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_4_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_4_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_4_clock; // @[Stab.scala 85:60]
  wire  cols_6_4_reset; // @[Stab.scala 85:60]
  wire  cols_6_4_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_4_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_4_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_4_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_4_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_4_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_4_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_6_4_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_4_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_6_4_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_4_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_4_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_4_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_4_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_4_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_4_clock; // @[Stab.scala 85:60]
  wire  cols_7_4_reset; // @[Stab.scala 85:60]
  wire  cols_7_4_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_4_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_4_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_4_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_4_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_4_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_4_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_7_4_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_4_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_7_4_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_4_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_4_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_4_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_4_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_4_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_4_clock; // @[Stab.scala 85:60]
  wire  cols_8_4_reset; // @[Stab.scala 85:60]
  wire  cols_8_4_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_4_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_4_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_4_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_4_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_4_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_4_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_8_4_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_4_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_8_4_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_4_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_4_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_4_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_4_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_4_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_4_clock; // @[Stab.scala 85:60]
  wire  cols_9_4_reset; // @[Stab.scala 85:60]
  wire  cols_9_4_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_4_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_4_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_4_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_4_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_4_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_4_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_9_4_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_4_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_9_4_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_4_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_4_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_4_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_4_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_4_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_4_clock; // @[Stab.scala 85:60]
  wire  cols_10_4_reset; // @[Stab.scala 85:60]
  wire  cols_10_4_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_4_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_4_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_4_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_4_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_4_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_4_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_10_4_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_4_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_10_4_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_4_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_4_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_4_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_4_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_4_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_4_clock; // @[Stab.scala 85:60]
  wire  cols_11_4_reset; // @[Stab.scala 85:60]
  wire  cols_11_4_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_4_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_4_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_4_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_4_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_4_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_4_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_11_4_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_4_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_11_4_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_4_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_4_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_4_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_4_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_4_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_4_clock; // @[Stab.scala 85:60]
  wire  cols_12_4_reset; // @[Stab.scala 85:60]
  wire  cols_12_4_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_4_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_4_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_4_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_4_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_4_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_4_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_12_4_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_4_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_12_4_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_4_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_4_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_4_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_4_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_4_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_4_clock; // @[Stab.scala 85:60]
  wire  cols_13_4_reset; // @[Stab.scala 85:60]
  wire  cols_13_4_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_4_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_4_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_4_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_4_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_4_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_4_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_13_4_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_4_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_13_4_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_4_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_4_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_4_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_4_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_4_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_4_clock; // @[Stab.scala 85:60]
  wire  cols_14_4_reset; // @[Stab.scala 85:60]
  wire  cols_14_4_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_4_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_4_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_4_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_4_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_4_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_4_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_14_4_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_4_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_14_4_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_4_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_4_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_4_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_4_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_4_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_4_clock; // @[Stab.scala 85:60]
  wire  cols_15_4_reset; // @[Stab.scala 85:60]
  wire  cols_15_4_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_4_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_4_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_4_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_4_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_4_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_4_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_15_4_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_4_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_15_4_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_4_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_4_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_4_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_4_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_4_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_5_clock; // @[Stab.scala 85:60]
  wire  cols_0_5_reset; // @[Stab.scala 85:60]
  wire  cols_0_5_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_5_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_5_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_5_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_5_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_5_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_5_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_0_5_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_5_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_0_5_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_5_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_5_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_5_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_5_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_5_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_5_clock; // @[Stab.scala 85:60]
  wire  cols_1_5_reset; // @[Stab.scala 85:60]
  wire  cols_1_5_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_5_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_5_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_5_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_5_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_5_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_5_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_1_5_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_5_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_1_5_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_5_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_5_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_5_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_5_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_5_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_5_clock; // @[Stab.scala 85:60]
  wire  cols_2_5_reset; // @[Stab.scala 85:60]
  wire  cols_2_5_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_5_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_5_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_5_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_5_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_5_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_5_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_2_5_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_5_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_2_5_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_5_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_5_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_5_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_5_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_5_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_5_clock; // @[Stab.scala 85:60]
  wire  cols_3_5_reset; // @[Stab.scala 85:60]
  wire  cols_3_5_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_5_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_5_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_5_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_5_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_5_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_5_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_3_5_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_5_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_3_5_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_5_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_5_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_5_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_5_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_5_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_5_clock; // @[Stab.scala 85:60]
  wire  cols_4_5_reset; // @[Stab.scala 85:60]
  wire  cols_4_5_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_5_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_5_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_5_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_5_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_5_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_5_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_4_5_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_5_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_4_5_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_5_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_5_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_5_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_5_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_5_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_5_clock; // @[Stab.scala 85:60]
  wire  cols_5_5_reset; // @[Stab.scala 85:60]
  wire  cols_5_5_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_5_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_5_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_5_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_5_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_5_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_5_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_5_5_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_5_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_5_5_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_5_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_5_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_5_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_5_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_5_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_5_clock; // @[Stab.scala 85:60]
  wire  cols_6_5_reset; // @[Stab.scala 85:60]
  wire  cols_6_5_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_5_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_5_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_5_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_5_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_5_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_5_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_6_5_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_5_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_6_5_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_5_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_5_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_5_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_5_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_5_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_5_clock; // @[Stab.scala 85:60]
  wire  cols_7_5_reset; // @[Stab.scala 85:60]
  wire  cols_7_5_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_5_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_5_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_5_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_5_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_5_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_5_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_7_5_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_5_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_7_5_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_5_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_5_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_5_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_5_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_5_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_5_clock; // @[Stab.scala 85:60]
  wire  cols_8_5_reset; // @[Stab.scala 85:60]
  wire  cols_8_5_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_5_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_5_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_5_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_5_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_5_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_5_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_8_5_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_5_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_8_5_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_5_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_5_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_5_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_5_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_5_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_5_clock; // @[Stab.scala 85:60]
  wire  cols_9_5_reset; // @[Stab.scala 85:60]
  wire  cols_9_5_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_5_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_5_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_5_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_5_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_5_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_5_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_9_5_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_5_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_9_5_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_5_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_5_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_5_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_5_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_5_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_5_clock; // @[Stab.scala 85:60]
  wire  cols_10_5_reset; // @[Stab.scala 85:60]
  wire  cols_10_5_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_5_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_5_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_5_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_5_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_5_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_5_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_10_5_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_5_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_10_5_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_5_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_5_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_5_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_5_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_5_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_5_clock; // @[Stab.scala 85:60]
  wire  cols_11_5_reset; // @[Stab.scala 85:60]
  wire  cols_11_5_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_5_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_5_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_5_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_5_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_5_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_5_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_11_5_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_5_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_11_5_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_5_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_5_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_5_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_5_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_5_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_5_clock; // @[Stab.scala 85:60]
  wire  cols_12_5_reset; // @[Stab.scala 85:60]
  wire  cols_12_5_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_5_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_5_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_5_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_5_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_5_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_5_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_12_5_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_5_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_12_5_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_5_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_5_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_5_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_5_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_5_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_5_clock; // @[Stab.scala 85:60]
  wire  cols_13_5_reset; // @[Stab.scala 85:60]
  wire  cols_13_5_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_5_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_5_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_5_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_5_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_5_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_5_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_13_5_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_5_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_13_5_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_5_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_5_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_5_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_5_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_5_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_5_clock; // @[Stab.scala 85:60]
  wire  cols_14_5_reset; // @[Stab.scala 85:60]
  wire  cols_14_5_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_5_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_5_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_5_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_5_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_5_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_5_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_14_5_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_5_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_14_5_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_5_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_5_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_5_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_5_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_5_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_5_clock; // @[Stab.scala 85:60]
  wire  cols_15_5_reset; // @[Stab.scala 85:60]
  wire  cols_15_5_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_5_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_5_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_5_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_5_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_5_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_5_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_15_5_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_5_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_15_5_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_5_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_5_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_5_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_5_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_5_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_6_clock; // @[Stab.scala 85:60]
  wire  cols_0_6_reset; // @[Stab.scala 85:60]
  wire  cols_0_6_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_6_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_6_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_6_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_6_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_6_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_6_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_0_6_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_6_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_0_6_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_6_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_6_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_6_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_6_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_6_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_6_clock; // @[Stab.scala 85:60]
  wire  cols_1_6_reset; // @[Stab.scala 85:60]
  wire  cols_1_6_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_6_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_6_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_6_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_6_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_6_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_6_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_1_6_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_6_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_1_6_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_6_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_6_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_6_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_6_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_6_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_6_clock; // @[Stab.scala 85:60]
  wire  cols_2_6_reset; // @[Stab.scala 85:60]
  wire  cols_2_6_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_6_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_6_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_6_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_6_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_6_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_6_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_2_6_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_6_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_2_6_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_6_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_6_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_6_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_6_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_6_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_6_clock; // @[Stab.scala 85:60]
  wire  cols_3_6_reset; // @[Stab.scala 85:60]
  wire  cols_3_6_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_6_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_6_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_6_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_6_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_6_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_6_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_3_6_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_6_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_3_6_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_6_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_6_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_6_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_6_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_6_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_6_clock; // @[Stab.scala 85:60]
  wire  cols_4_6_reset; // @[Stab.scala 85:60]
  wire  cols_4_6_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_6_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_6_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_6_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_6_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_6_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_6_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_4_6_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_6_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_4_6_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_6_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_6_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_6_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_6_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_6_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_6_clock; // @[Stab.scala 85:60]
  wire  cols_5_6_reset; // @[Stab.scala 85:60]
  wire  cols_5_6_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_6_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_6_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_6_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_6_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_6_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_6_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_5_6_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_6_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_5_6_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_6_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_6_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_6_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_6_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_6_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_6_clock; // @[Stab.scala 85:60]
  wire  cols_6_6_reset; // @[Stab.scala 85:60]
  wire  cols_6_6_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_6_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_6_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_6_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_6_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_6_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_6_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_6_6_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_6_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_6_6_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_6_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_6_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_6_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_6_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_6_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_6_clock; // @[Stab.scala 85:60]
  wire  cols_7_6_reset; // @[Stab.scala 85:60]
  wire  cols_7_6_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_6_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_6_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_6_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_6_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_6_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_6_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_7_6_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_6_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_7_6_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_6_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_6_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_6_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_6_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_6_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_6_clock; // @[Stab.scala 85:60]
  wire  cols_8_6_reset; // @[Stab.scala 85:60]
  wire  cols_8_6_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_6_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_6_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_6_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_6_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_6_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_6_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_8_6_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_6_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_8_6_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_6_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_6_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_6_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_6_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_6_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_6_clock; // @[Stab.scala 85:60]
  wire  cols_9_6_reset; // @[Stab.scala 85:60]
  wire  cols_9_6_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_6_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_6_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_6_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_6_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_6_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_6_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_9_6_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_6_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_9_6_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_6_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_6_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_6_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_6_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_6_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_6_clock; // @[Stab.scala 85:60]
  wire  cols_10_6_reset; // @[Stab.scala 85:60]
  wire  cols_10_6_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_6_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_6_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_6_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_6_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_6_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_6_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_10_6_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_6_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_10_6_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_6_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_6_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_6_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_6_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_6_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_6_clock; // @[Stab.scala 85:60]
  wire  cols_11_6_reset; // @[Stab.scala 85:60]
  wire  cols_11_6_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_6_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_6_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_6_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_6_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_6_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_6_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_11_6_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_6_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_11_6_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_6_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_6_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_6_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_6_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_6_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_6_clock; // @[Stab.scala 85:60]
  wire  cols_12_6_reset; // @[Stab.scala 85:60]
  wire  cols_12_6_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_6_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_6_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_6_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_6_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_6_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_6_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_12_6_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_6_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_12_6_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_6_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_6_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_6_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_6_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_6_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_6_clock; // @[Stab.scala 85:60]
  wire  cols_13_6_reset; // @[Stab.scala 85:60]
  wire  cols_13_6_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_6_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_6_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_6_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_6_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_6_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_6_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_13_6_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_6_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_13_6_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_6_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_6_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_6_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_6_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_6_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_6_clock; // @[Stab.scala 85:60]
  wire  cols_14_6_reset; // @[Stab.scala 85:60]
  wire  cols_14_6_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_6_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_6_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_6_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_6_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_6_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_6_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_14_6_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_6_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_14_6_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_6_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_6_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_6_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_6_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_6_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_6_clock; // @[Stab.scala 85:60]
  wire  cols_15_6_reset; // @[Stab.scala 85:60]
  wire  cols_15_6_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_6_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_6_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_6_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_6_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_6_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_6_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_15_6_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_6_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_15_6_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_6_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_6_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_6_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_6_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_6_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_7_clock; // @[Stab.scala 85:60]
  wire  cols_0_7_reset; // @[Stab.scala 85:60]
  wire  cols_0_7_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_7_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_7_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_7_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_7_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_7_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_7_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_0_7_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_7_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_0_7_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_7_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_7_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_7_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_7_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_7_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_7_clock; // @[Stab.scala 85:60]
  wire  cols_1_7_reset; // @[Stab.scala 85:60]
  wire  cols_1_7_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_7_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_7_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_7_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_7_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_7_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_7_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_1_7_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_7_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_1_7_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_7_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_7_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_7_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_7_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_7_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_7_clock; // @[Stab.scala 85:60]
  wire  cols_2_7_reset; // @[Stab.scala 85:60]
  wire  cols_2_7_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_7_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_7_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_7_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_7_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_7_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_7_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_2_7_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_7_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_2_7_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_7_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_7_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_7_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_7_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_7_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_7_clock; // @[Stab.scala 85:60]
  wire  cols_3_7_reset; // @[Stab.scala 85:60]
  wire  cols_3_7_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_7_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_7_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_7_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_7_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_7_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_7_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_3_7_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_7_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_3_7_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_7_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_7_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_7_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_7_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_7_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_7_clock; // @[Stab.scala 85:60]
  wire  cols_4_7_reset; // @[Stab.scala 85:60]
  wire  cols_4_7_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_7_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_7_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_7_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_7_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_7_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_7_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_4_7_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_7_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_4_7_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_7_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_7_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_7_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_7_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_7_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_7_clock; // @[Stab.scala 85:60]
  wire  cols_5_7_reset; // @[Stab.scala 85:60]
  wire  cols_5_7_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_7_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_7_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_7_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_7_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_7_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_7_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_5_7_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_7_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_5_7_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_7_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_7_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_7_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_7_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_7_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_7_clock; // @[Stab.scala 85:60]
  wire  cols_6_7_reset; // @[Stab.scala 85:60]
  wire  cols_6_7_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_7_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_7_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_7_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_7_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_7_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_7_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_6_7_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_7_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_6_7_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_7_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_7_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_7_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_7_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_7_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_7_clock; // @[Stab.scala 85:60]
  wire  cols_7_7_reset; // @[Stab.scala 85:60]
  wire  cols_7_7_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_7_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_7_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_7_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_7_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_7_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_7_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_7_7_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_7_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_7_7_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_7_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_7_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_7_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_7_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_7_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_7_clock; // @[Stab.scala 85:60]
  wire  cols_8_7_reset; // @[Stab.scala 85:60]
  wire  cols_8_7_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_7_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_7_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_7_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_7_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_7_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_7_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_8_7_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_7_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_8_7_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_7_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_7_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_7_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_7_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_7_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_7_clock; // @[Stab.scala 85:60]
  wire  cols_9_7_reset; // @[Stab.scala 85:60]
  wire  cols_9_7_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_7_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_7_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_7_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_7_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_7_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_7_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_9_7_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_7_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_9_7_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_7_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_7_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_7_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_7_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_7_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_7_clock; // @[Stab.scala 85:60]
  wire  cols_10_7_reset; // @[Stab.scala 85:60]
  wire  cols_10_7_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_7_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_7_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_7_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_7_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_7_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_7_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_10_7_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_7_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_10_7_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_7_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_7_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_7_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_7_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_7_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_7_clock; // @[Stab.scala 85:60]
  wire  cols_11_7_reset; // @[Stab.scala 85:60]
  wire  cols_11_7_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_7_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_7_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_7_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_7_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_7_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_7_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_11_7_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_7_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_11_7_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_7_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_7_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_7_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_7_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_7_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_7_clock; // @[Stab.scala 85:60]
  wire  cols_12_7_reset; // @[Stab.scala 85:60]
  wire  cols_12_7_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_7_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_7_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_7_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_7_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_7_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_7_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_12_7_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_7_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_12_7_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_7_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_7_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_7_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_7_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_7_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_7_clock; // @[Stab.scala 85:60]
  wire  cols_13_7_reset; // @[Stab.scala 85:60]
  wire  cols_13_7_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_7_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_7_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_7_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_7_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_7_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_7_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_13_7_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_7_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_13_7_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_7_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_7_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_7_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_7_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_7_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_7_clock; // @[Stab.scala 85:60]
  wire  cols_14_7_reset; // @[Stab.scala 85:60]
  wire  cols_14_7_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_7_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_7_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_7_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_7_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_7_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_7_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_14_7_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_7_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_14_7_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_7_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_7_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_7_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_7_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_7_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_7_clock; // @[Stab.scala 85:60]
  wire  cols_15_7_reset; // @[Stab.scala 85:60]
  wire  cols_15_7_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_7_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_7_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_7_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_7_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_7_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_7_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_15_7_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_7_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_15_7_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_7_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_7_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_7_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_7_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_7_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_8_clock; // @[Stab.scala 85:60]
  wire  cols_0_8_reset; // @[Stab.scala 85:60]
  wire  cols_0_8_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_8_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_8_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_8_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_8_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_8_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_8_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_0_8_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_8_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_0_8_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_8_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_8_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_8_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_8_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_8_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_8_clock; // @[Stab.scala 85:60]
  wire  cols_1_8_reset; // @[Stab.scala 85:60]
  wire  cols_1_8_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_8_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_8_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_8_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_8_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_8_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_8_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_1_8_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_8_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_1_8_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_8_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_8_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_8_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_8_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_8_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_8_clock; // @[Stab.scala 85:60]
  wire  cols_2_8_reset; // @[Stab.scala 85:60]
  wire  cols_2_8_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_8_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_8_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_8_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_8_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_8_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_8_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_2_8_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_8_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_2_8_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_8_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_8_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_8_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_8_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_8_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_8_clock; // @[Stab.scala 85:60]
  wire  cols_3_8_reset; // @[Stab.scala 85:60]
  wire  cols_3_8_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_8_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_8_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_8_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_8_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_8_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_8_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_3_8_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_8_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_3_8_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_8_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_8_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_8_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_8_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_8_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_8_clock; // @[Stab.scala 85:60]
  wire  cols_4_8_reset; // @[Stab.scala 85:60]
  wire  cols_4_8_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_8_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_8_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_8_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_8_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_8_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_8_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_4_8_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_8_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_4_8_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_8_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_8_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_8_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_8_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_8_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_8_clock; // @[Stab.scala 85:60]
  wire  cols_5_8_reset; // @[Stab.scala 85:60]
  wire  cols_5_8_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_8_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_8_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_8_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_8_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_8_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_8_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_5_8_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_8_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_5_8_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_8_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_8_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_8_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_8_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_8_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_8_clock; // @[Stab.scala 85:60]
  wire  cols_6_8_reset; // @[Stab.scala 85:60]
  wire  cols_6_8_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_8_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_8_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_8_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_8_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_8_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_8_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_6_8_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_8_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_6_8_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_8_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_8_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_8_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_8_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_8_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_8_clock; // @[Stab.scala 85:60]
  wire  cols_7_8_reset; // @[Stab.scala 85:60]
  wire  cols_7_8_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_8_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_8_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_8_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_8_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_8_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_8_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_7_8_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_8_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_7_8_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_8_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_8_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_8_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_8_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_8_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_8_clock; // @[Stab.scala 85:60]
  wire  cols_8_8_reset; // @[Stab.scala 85:60]
  wire  cols_8_8_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_8_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_8_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_8_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_8_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_8_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_8_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_8_8_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_8_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_8_8_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_8_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_8_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_8_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_8_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_8_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_8_clock; // @[Stab.scala 85:60]
  wire  cols_9_8_reset; // @[Stab.scala 85:60]
  wire  cols_9_8_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_8_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_8_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_8_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_8_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_8_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_8_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_9_8_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_8_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_9_8_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_8_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_8_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_8_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_8_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_8_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_8_clock; // @[Stab.scala 85:60]
  wire  cols_10_8_reset; // @[Stab.scala 85:60]
  wire  cols_10_8_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_8_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_8_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_8_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_8_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_8_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_8_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_10_8_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_8_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_10_8_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_8_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_8_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_8_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_8_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_8_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_8_clock; // @[Stab.scala 85:60]
  wire  cols_11_8_reset; // @[Stab.scala 85:60]
  wire  cols_11_8_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_8_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_8_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_8_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_8_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_8_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_8_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_11_8_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_8_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_11_8_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_8_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_8_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_8_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_8_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_8_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_8_clock; // @[Stab.scala 85:60]
  wire  cols_12_8_reset; // @[Stab.scala 85:60]
  wire  cols_12_8_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_8_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_8_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_8_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_8_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_8_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_8_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_12_8_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_8_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_12_8_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_8_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_8_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_8_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_8_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_8_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_8_clock; // @[Stab.scala 85:60]
  wire  cols_13_8_reset; // @[Stab.scala 85:60]
  wire  cols_13_8_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_8_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_8_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_8_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_8_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_8_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_8_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_13_8_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_8_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_13_8_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_8_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_8_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_8_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_8_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_8_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_8_clock; // @[Stab.scala 85:60]
  wire  cols_14_8_reset; // @[Stab.scala 85:60]
  wire  cols_14_8_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_8_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_8_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_8_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_8_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_8_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_8_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_14_8_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_8_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_14_8_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_8_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_8_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_8_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_8_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_8_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_8_clock; // @[Stab.scala 85:60]
  wire  cols_15_8_reset; // @[Stab.scala 85:60]
  wire  cols_15_8_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_8_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_8_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_8_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_8_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_8_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_8_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_15_8_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_8_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_15_8_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_8_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_8_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_8_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_8_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_8_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_9_clock; // @[Stab.scala 85:60]
  wire  cols_0_9_reset; // @[Stab.scala 85:60]
  wire  cols_0_9_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_9_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_9_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_9_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_9_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_9_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_9_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_0_9_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_9_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_0_9_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_9_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_9_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_9_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_9_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_9_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_9_clock; // @[Stab.scala 85:60]
  wire  cols_1_9_reset; // @[Stab.scala 85:60]
  wire  cols_1_9_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_9_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_9_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_9_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_9_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_9_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_9_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_1_9_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_9_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_1_9_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_9_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_9_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_9_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_9_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_9_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_9_clock; // @[Stab.scala 85:60]
  wire  cols_2_9_reset; // @[Stab.scala 85:60]
  wire  cols_2_9_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_9_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_9_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_9_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_9_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_9_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_9_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_2_9_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_9_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_2_9_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_9_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_9_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_9_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_9_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_9_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_9_clock; // @[Stab.scala 85:60]
  wire  cols_3_9_reset; // @[Stab.scala 85:60]
  wire  cols_3_9_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_9_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_9_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_9_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_9_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_9_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_9_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_3_9_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_9_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_3_9_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_9_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_9_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_9_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_9_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_9_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_9_clock; // @[Stab.scala 85:60]
  wire  cols_4_9_reset; // @[Stab.scala 85:60]
  wire  cols_4_9_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_9_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_9_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_9_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_9_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_9_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_9_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_4_9_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_9_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_4_9_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_9_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_9_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_9_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_9_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_9_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_9_clock; // @[Stab.scala 85:60]
  wire  cols_5_9_reset; // @[Stab.scala 85:60]
  wire  cols_5_9_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_9_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_9_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_9_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_9_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_9_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_9_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_5_9_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_9_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_5_9_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_9_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_9_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_9_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_9_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_9_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_9_clock; // @[Stab.scala 85:60]
  wire  cols_6_9_reset; // @[Stab.scala 85:60]
  wire  cols_6_9_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_9_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_9_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_9_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_9_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_9_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_9_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_6_9_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_9_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_6_9_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_9_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_9_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_9_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_9_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_9_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_9_clock; // @[Stab.scala 85:60]
  wire  cols_7_9_reset; // @[Stab.scala 85:60]
  wire  cols_7_9_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_9_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_9_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_9_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_9_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_9_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_9_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_7_9_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_9_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_7_9_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_9_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_9_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_9_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_9_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_9_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_9_clock; // @[Stab.scala 85:60]
  wire  cols_8_9_reset; // @[Stab.scala 85:60]
  wire  cols_8_9_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_9_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_9_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_9_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_9_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_9_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_9_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_8_9_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_9_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_8_9_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_9_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_9_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_9_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_9_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_9_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_9_clock; // @[Stab.scala 85:60]
  wire  cols_9_9_reset; // @[Stab.scala 85:60]
  wire  cols_9_9_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_9_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_9_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_9_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_9_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_9_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_9_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_9_9_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_9_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_9_9_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_9_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_9_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_9_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_9_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_9_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_9_clock; // @[Stab.scala 85:60]
  wire  cols_10_9_reset; // @[Stab.scala 85:60]
  wire  cols_10_9_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_9_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_9_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_9_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_9_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_9_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_9_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_10_9_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_9_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_10_9_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_9_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_9_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_9_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_9_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_9_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_9_clock; // @[Stab.scala 85:60]
  wire  cols_11_9_reset; // @[Stab.scala 85:60]
  wire  cols_11_9_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_9_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_9_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_9_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_9_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_9_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_9_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_11_9_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_9_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_11_9_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_9_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_9_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_9_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_9_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_9_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_9_clock; // @[Stab.scala 85:60]
  wire  cols_12_9_reset; // @[Stab.scala 85:60]
  wire  cols_12_9_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_9_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_9_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_9_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_9_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_9_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_9_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_12_9_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_9_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_12_9_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_9_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_9_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_9_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_9_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_9_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_9_clock; // @[Stab.scala 85:60]
  wire  cols_13_9_reset; // @[Stab.scala 85:60]
  wire  cols_13_9_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_9_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_9_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_9_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_9_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_9_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_9_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_13_9_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_9_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_13_9_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_9_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_9_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_9_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_9_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_9_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_9_clock; // @[Stab.scala 85:60]
  wire  cols_14_9_reset; // @[Stab.scala 85:60]
  wire  cols_14_9_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_9_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_9_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_9_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_9_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_9_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_9_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_14_9_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_9_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_14_9_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_9_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_9_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_9_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_9_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_9_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_9_clock; // @[Stab.scala 85:60]
  wire  cols_15_9_reset; // @[Stab.scala 85:60]
  wire  cols_15_9_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_9_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_9_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_9_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_9_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_9_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_9_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_15_9_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_9_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_15_9_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_9_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_9_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_9_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_9_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_9_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_10_clock; // @[Stab.scala 85:60]
  wire  cols_0_10_reset; // @[Stab.scala 85:60]
  wire  cols_0_10_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_10_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_10_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_10_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_10_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_10_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_10_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_0_10_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_10_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_0_10_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_10_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_10_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_10_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_10_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_10_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_10_clock; // @[Stab.scala 85:60]
  wire  cols_1_10_reset; // @[Stab.scala 85:60]
  wire  cols_1_10_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_10_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_10_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_10_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_10_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_10_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_10_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_1_10_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_10_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_1_10_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_10_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_10_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_10_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_10_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_10_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_10_clock; // @[Stab.scala 85:60]
  wire  cols_2_10_reset; // @[Stab.scala 85:60]
  wire  cols_2_10_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_10_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_10_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_10_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_10_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_10_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_10_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_2_10_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_10_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_2_10_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_10_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_10_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_10_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_10_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_10_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_10_clock; // @[Stab.scala 85:60]
  wire  cols_3_10_reset; // @[Stab.scala 85:60]
  wire  cols_3_10_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_10_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_10_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_10_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_10_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_10_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_10_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_3_10_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_10_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_3_10_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_10_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_10_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_10_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_10_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_10_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_10_clock; // @[Stab.scala 85:60]
  wire  cols_4_10_reset; // @[Stab.scala 85:60]
  wire  cols_4_10_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_10_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_10_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_10_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_10_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_10_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_10_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_4_10_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_10_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_4_10_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_10_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_10_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_10_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_10_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_10_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_10_clock; // @[Stab.scala 85:60]
  wire  cols_5_10_reset; // @[Stab.scala 85:60]
  wire  cols_5_10_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_10_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_10_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_10_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_10_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_10_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_10_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_5_10_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_10_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_5_10_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_10_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_10_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_10_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_10_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_10_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_10_clock; // @[Stab.scala 85:60]
  wire  cols_6_10_reset; // @[Stab.scala 85:60]
  wire  cols_6_10_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_10_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_10_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_10_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_10_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_10_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_10_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_6_10_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_10_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_6_10_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_10_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_10_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_10_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_10_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_10_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_10_clock; // @[Stab.scala 85:60]
  wire  cols_7_10_reset; // @[Stab.scala 85:60]
  wire  cols_7_10_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_10_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_10_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_10_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_10_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_10_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_10_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_7_10_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_10_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_7_10_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_10_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_10_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_10_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_10_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_10_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_10_clock; // @[Stab.scala 85:60]
  wire  cols_8_10_reset; // @[Stab.scala 85:60]
  wire  cols_8_10_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_10_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_10_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_10_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_10_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_10_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_10_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_8_10_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_10_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_8_10_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_10_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_10_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_10_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_10_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_10_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_10_clock; // @[Stab.scala 85:60]
  wire  cols_9_10_reset; // @[Stab.scala 85:60]
  wire  cols_9_10_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_10_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_10_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_10_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_10_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_10_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_10_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_9_10_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_10_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_9_10_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_10_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_10_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_10_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_10_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_10_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_10_clock; // @[Stab.scala 85:60]
  wire  cols_10_10_reset; // @[Stab.scala 85:60]
  wire  cols_10_10_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_10_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_10_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_10_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_10_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_10_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_10_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_10_10_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_10_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_10_10_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_10_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_10_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_10_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_10_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_10_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_10_clock; // @[Stab.scala 85:60]
  wire  cols_11_10_reset; // @[Stab.scala 85:60]
  wire  cols_11_10_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_10_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_10_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_10_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_10_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_10_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_10_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_11_10_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_10_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_11_10_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_10_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_10_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_10_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_10_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_10_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_10_clock; // @[Stab.scala 85:60]
  wire  cols_12_10_reset; // @[Stab.scala 85:60]
  wire  cols_12_10_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_10_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_10_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_10_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_10_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_10_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_10_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_12_10_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_10_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_12_10_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_10_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_10_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_10_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_10_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_10_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_10_clock; // @[Stab.scala 85:60]
  wire  cols_13_10_reset; // @[Stab.scala 85:60]
  wire  cols_13_10_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_10_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_10_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_10_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_10_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_10_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_10_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_13_10_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_10_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_13_10_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_10_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_10_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_10_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_10_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_10_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_10_clock; // @[Stab.scala 85:60]
  wire  cols_14_10_reset; // @[Stab.scala 85:60]
  wire  cols_14_10_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_10_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_10_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_10_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_10_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_10_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_10_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_14_10_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_10_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_14_10_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_10_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_10_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_10_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_10_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_10_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_10_clock; // @[Stab.scala 85:60]
  wire  cols_15_10_reset; // @[Stab.scala 85:60]
  wire  cols_15_10_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_10_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_10_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_10_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_10_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_10_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_10_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_15_10_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_10_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_15_10_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_10_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_10_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_10_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_10_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_10_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_11_clock; // @[Stab.scala 85:60]
  wire  cols_0_11_reset; // @[Stab.scala 85:60]
  wire  cols_0_11_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_11_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_11_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_11_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_11_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_11_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_11_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_0_11_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_11_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_0_11_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_11_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_11_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_11_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_11_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_11_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_11_clock; // @[Stab.scala 85:60]
  wire  cols_1_11_reset; // @[Stab.scala 85:60]
  wire  cols_1_11_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_11_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_11_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_11_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_11_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_11_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_11_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_1_11_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_11_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_1_11_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_11_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_11_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_11_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_11_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_11_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_11_clock; // @[Stab.scala 85:60]
  wire  cols_2_11_reset; // @[Stab.scala 85:60]
  wire  cols_2_11_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_11_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_11_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_11_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_11_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_11_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_11_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_2_11_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_11_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_2_11_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_11_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_11_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_11_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_11_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_11_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_11_clock; // @[Stab.scala 85:60]
  wire  cols_3_11_reset; // @[Stab.scala 85:60]
  wire  cols_3_11_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_11_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_11_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_11_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_11_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_11_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_11_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_3_11_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_11_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_3_11_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_11_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_11_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_11_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_11_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_11_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_11_clock; // @[Stab.scala 85:60]
  wire  cols_4_11_reset; // @[Stab.scala 85:60]
  wire  cols_4_11_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_11_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_11_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_11_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_11_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_11_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_11_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_4_11_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_11_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_4_11_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_11_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_11_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_11_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_11_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_11_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_11_clock; // @[Stab.scala 85:60]
  wire  cols_5_11_reset; // @[Stab.scala 85:60]
  wire  cols_5_11_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_11_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_11_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_11_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_11_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_11_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_11_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_5_11_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_11_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_5_11_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_11_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_11_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_11_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_11_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_11_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_11_clock; // @[Stab.scala 85:60]
  wire  cols_6_11_reset; // @[Stab.scala 85:60]
  wire  cols_6_11_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_11_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_11_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_11_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_11_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_11_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_11_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_6_11_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_11_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_6_11_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_11_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_11_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_11_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_11_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_11_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_11_clock; // @[Stab.scala 85:60]
  wire  cols_7_11_reset; // @[Stab.scala 85:60]
  wire  cols_7_11_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_11_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_11_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_11_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_11_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_11_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_11_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_7_11_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_11_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_7_11_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_11_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_11_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_11_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_11_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_11_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_11_clock; // @[Stab.scala 85:60]
  wire  cols_8_11_reset; // @[Stab.scala 85:60]
  wire  cols_8_11_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_11_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_11_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_11_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_11_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_11_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_11_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_8_11_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_11_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_8_11_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_11_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_11_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_11_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_11_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_11_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_11_clock; // @[Stab.scala 85:60]
  wire  cols_9_11_reset; // @[Stab.scala 85:60]
  wire  cols_9_11_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_11_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_11_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_11_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_11_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_11_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_11_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_9_11_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_11_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_9_11_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_11_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_11_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_11_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_11_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_11_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_11_clock; // @[Stab.scala 85:60]
  wire  cols_10_11_reset; // @[Stab.scala 85:60]
  wire  cols_10_11_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_11_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_11_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_11_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_11_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_11_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_11_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_10_11_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_11_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_10_11_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_11_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_11_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_11_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_11_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_11_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_11_clock; // @[Stab.scala 85:60]
  wire  cols_11_11_reset; // @[Stab.scala 85:60]
  wire  cols_11_11_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_11_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_11_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_11_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_11_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_11_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_11_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_11_11_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_11_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_11_11_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_11_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_11_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_11_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_11_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_11_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_11_clock; // @[Stab.scala 85:60]
  wire  cols_12_11_reset; // @[Stab.scala 85:60]
  wire  cols_12_11_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_11_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_11_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_11_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_11_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_11_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_11_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_12_11_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_11_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_12_11_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_11_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_11_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_11_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_11_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_11_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_11_clock; // @[Stab.scala 85:60]
  wire  cols_13_11_reset; // @[Stab.scala 85:60]
  wire  cols_13_11_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_11_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_11_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_11_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_11_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_11_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_11_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_13_11_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_11_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_13_11_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_11_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_11_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_11_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_11_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_11_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_11_clock; // @[Stab.scala 85:60]
  wire  cols_14_11_reset; // @[Stab.scala 85:60]
  wire  cols_14_11_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_11_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_11_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_11_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_11_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_11_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_11_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_14_11_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_11_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_14_11_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_11_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_11_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_11_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_11_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_11_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_11_clock; // @[Stab.scala 85:60]
  wire  cols_15_11_reset; // @[Stab.scala 85:60]
  wire  cols_15_11_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_11_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_11_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_11_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_11_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_11_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_11_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_15_11_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_11_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_15_11_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_11_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_11_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_11_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_11_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_11_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_12_clock; // @[Stab.scala 85:60]
  wire  cols_0_12_reset; // @[Stab.scala 85:60]
  wire  cols_0_12_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_12_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_12_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_12_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_12_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_12_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_12_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_0_12_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_12_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_0_12_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_12_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_12_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_12_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_12_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_12_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_12_clock; // @[Stab.scala 85:60]
  wire  cols_1_12_reset; // @[Stab.scala 85:60]
  wire  cols_1_12_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_12_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_12_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_12_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_12_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_12_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_12_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_1_12_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_12_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_1_12_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_12_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_12_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_12_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_12_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_12_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_12_clock; // @[Stab.scala 85:60]
  wire  cols_2_12_reset; // @[Stab.scala 85:60]
  wire  cols_2_12_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_12_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_12_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_12_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_12_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_12_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_12_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_2_12_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_12_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_2_12_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_12_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_12_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_12_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_12_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_12_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_12_clock; // @[Stab.scala 85:60]
  wire  cols_3_12_reset; // @[Stab.scala 85:60]
  wire  cols_3_12_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_12_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_12_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_12_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_12_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_12_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_12_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_3_12_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_12_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_3_12_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_12_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_12_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_12_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_12_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_12_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_12_clock; // @[Stab.scala 85:60]
  wire  cols_4_12_reset; // @[Stab.scala 85:60]
  wire  cols_4_12_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_12_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_12_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_12_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_12_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_12_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_12_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_4_12_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_12_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_4_12_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_12_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_12_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_12_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_12_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_12_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_12_clock; // @[Stab.scala 85:60]
  wire  cols_5_12_reset; // @[Stab.scala 85:60]
  wire  cols_5_12_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_12_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_12_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_12_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_12_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_12_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_12_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_5_12_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_12_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_5_12_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_12_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_12_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_12_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_12_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_12_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_12_clock; // @[Stab.scala 85:60]
  wire  cols_6_12_reset; // @[Stab.scala 85:60]
  wire  cols_6_12_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_12_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_12_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_12_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_12_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_12_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_12_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_6_12_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_12_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_6_12_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_12_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_12_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_12_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_12_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_12_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_12_clock; // @[Stab.scala 85:60]
  wire  cols_7_12_reset; // @[Stab.scala 85:60]
  wire  cols_7_12_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_12_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_12_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_12_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_12_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_12_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_12_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_7_12_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_12_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_7_12_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_12_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_12_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_12_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_12_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_12_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_12_clock; // @[Stab.scala 85:60]
  wire  cols_8_12_reset; // @[Stab.scala 85:60]
  wire  cols_8_12_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_12_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_12_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_12_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_12_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_12_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_12_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_8_12_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_12_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_8_12_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_12_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_12_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_12_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_12_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_12_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_12_clock; // @[Stab.scala 85:60]
  wire  cols_9_12_reset; // @[Stab.scala 85:60]
  wire  cols_9_12_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_12_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_12_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_12_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_12_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_12_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_12_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_9_12_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_12_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_9_12_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_12_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_12_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_12_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_12_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_12_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_12_clock; // @[Stab.scala 85:60]
  wire  cols_10_12_reset; // @[Stab.scala 85:60]
  wire  cols_10_12_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_12_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_12_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_12_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_12_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_12_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_12_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_10_12_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_12_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_10_12_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_12_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_12_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_12_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_12_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_12_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_12_clock; // @[Stab.scala 85:60]
  wire  cols_11_12_reset; // @[Stab.scala 85:60]
  wire  cols_11_12_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_12_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_12_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_12_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_12_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_12_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_12_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_11_12_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_12_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_11_12_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_12_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_12_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_12_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_12_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_12_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_12_clock; // @[Stab.scala 85:60]
  wire  cols_12_12_reset; // @[Stab.scala 85:60]
  wire  cols_12_12_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_12_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_12_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_12_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_12_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_12_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_12_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_12_12_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_12_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_12_12_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_12_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_12_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_12_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_12_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_12_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_12_clock; // @[Stab.scala 85:60]
  wire  cols_13_12_reset; // @[Stab.scala 85:60]
  wire  cols_13_12_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_12_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_12_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_12_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_12_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_12_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_12_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_13_12_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_12_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_13_12_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_12_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_12_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_12_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_12_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_12_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_12_clock; // @[Stab.scala 85:60]
  wire  cols_14_12_reset; // @[Stab.scala 85:60]
  wire  cols_14_12_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_12_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_12_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_12_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_12_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_12_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_12_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_14_12_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_12_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_14_12_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_12_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_12_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_12_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_12_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_12_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_12_clock; // @[Stab.scala 85:60]
  wire  cols_15_12_reset; // @[Stab.scala 85:60]
  wire  cols_15_12_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_12_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_12_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_12_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_12_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_12_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_12_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_15_12_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_12_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_15_12_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_12_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_12_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_12_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_12_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_12_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_13_clock; // @[Stab.scala 85:60]
  wire  cols_0_13_reset; // @[Stab.scala 85:60]
  wire  cols_0_13_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_13_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_13_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_13_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_13_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_13_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_13_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_0_13_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_13_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_0_13_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_13_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_13_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_13_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_13_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_13_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_13_clock; // @[Stab.scala 85:60]
  wire  cols_1_13_reset; // @[Stab.scala 85:60]
  wire  cols_1_13_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_13_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_13_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_13_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_13_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_13_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_13_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_1_13_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_13_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_1_13_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_13_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_13_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_13_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_13_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_13_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_13_clock; // @[Stab.scala 85:60]
  wire  cols_2_13_reset; // @[Stab.scala 85:60]
  wire  cols_2_13_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_13_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_13_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_13_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_13_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_13_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_13_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_2_13_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_13_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_2_13_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_13_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_13_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_13_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_13_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_13_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_13_clock; // @[Stab.scala 85:60]
  wire  cols_3_13_reset; // @[Stab.scala 85:60]
  wire  cols_3_13_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_13_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_13_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_13_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_13_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_13_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_13_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_3_13_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_13_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_3_13_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_13_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_13_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_13_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_13_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_13_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_13_clock; // @[Stab.scala 85:60]
  wire  cols_4_13_reset; // @[Stab.scala 85:60]
  wire  cols_4_13_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_13_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_13_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_13_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_13_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_13_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_13_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_4_13_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_13_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_4_13_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_13_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_13_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_13_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_13_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_13_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_13_clock; // @[Stab.scala 85:60]
  wire  cols_5_13_reset; // @[Stab.scala 85:60]
  wire  cols_5_13_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_13_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_13_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_13_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_13_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_13_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_13_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_5_13_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_13_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_5_13_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_13_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_13_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_13_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_13_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_13_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_13_clock; // @[Stab.scala 85:60]
  wire  cols_6_13_reset; // @[Stab.scala 85:60]
  wire  cols_6_13_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_13_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_13_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_13_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_13_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_13_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_13_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_6_13_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_13_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_6_13_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_13_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_13_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_13_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_13_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_13_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_13_clock; // @[Stab.scala 85:60]
  wire  cols_7_13_reset; // @[Stab.scala 85:60]
  wire  cols_7_13_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_13_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_13_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_13_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_13_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_13_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_13_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_7_13_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_13_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_7_13_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_13_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_13_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_13_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_13_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_13_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_13_clock; // @[Stab.scala 85:60]
  wire  cols_8_13_reset; // @[Stab.scala 85:60]
  wire  cols_8_13_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_13_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_13_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_13_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_13_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_13_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_13_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_8_13_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_13_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_8_13_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_13_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_13_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_13_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_13_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_13_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_13_clock; // @[Stab.scala 85:60]
  wire  cols_9_13_reset; // @[Stab.scala 85:60]
  wire  cols_9_13_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_13_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_13_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_13_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_13_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_13_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_13_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_9_13_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_13_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_9_13_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_13_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_13_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_13_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_13_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_13_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_13_clock; // @[Stab.scala 85:60]
  wire  cols_10_13_reset; // @[Stab.scala 85:60]
  wire  cols_10_13_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_13_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_13_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_13_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_13_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_13_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_13_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_10_13_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_13_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_10_13_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_13_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_13_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_13_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_13_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_13_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_13_clock; // @[Stab.scala 85:60]
  wire  cols_11_13_reset; // @[Stab.scala 85:60]
  wire  cols_11_13_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_13_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_13_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_13_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_13_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_13_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_13_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_11_13_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_13_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_11_13_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_13_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_13_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_13_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_13_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_13_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_13_clock; // @[Stab.scala 85:60]
  wire  cols_12_13_reset; // @[Stab.scala 85:60]
  wire  cols_12_13_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_13_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_13_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_13_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_13_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_13_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_13_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_12_13_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_13_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_12_13_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_13_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_13_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_13_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_13_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_13_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_13_clock; // @[Stab.scala 85:60]
  wire  cols_13_13_reset; // @[Stab.scala 85:60]
  wire  cols_13_13_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_13_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_13_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_13_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_13_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_13_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_13_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_13_13_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_13_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_13_13_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_13_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_13_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_13_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_13_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_13_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_13_clock; // @[Stab.scala 85:60]
  wire  cols_14_13_reset; // @[Stab.scala 85:60]
  wire  cols_14_13_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_13_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_13_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_13_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_13_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_13_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_13_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_14_13_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_13_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_14_13_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_13_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_13_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_13_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_13_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_13_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_13_clock; // @[Stab.scala 85:60]
  wire  cols_15_13_reset; // @[Stab.scala 85:60]
  wire  cols_15_13_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_13_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_13_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_13_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_13_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_13_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_13_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_15_13_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_13_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_15_13_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_13_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_13_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_13_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_13_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_13_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_14_clock; // @[Stab.scala 85:60]
  wire  cols_0_14_reset; // @[Stab.scala 85:60]
  wire  cols_0_14_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_14_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_14_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_14_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_14_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_14_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_14_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_0_14_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_14_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_0_14_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_14_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_14_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_14_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_14_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_14_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_14_clock; // @[Stab.scala 85:60]
  wire  cols_1_14_reset; // @[Stab.scala 85:60]
  wire  cols_1_14_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_14_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_14_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_14_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_14_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_14_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_14_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_1_14_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_14_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_1_14_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_14_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_14_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_14_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_14_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_14_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_14_clock; // @[Stab.scala 85:60]
  wire  cols_2_14_reset; // @[Stab.scala 85:60]
  wire  cols_2_14_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_14_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_14_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_14_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_14_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_14_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_14_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_2_14_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_14_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_2_14_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_14_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_14_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_14_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_14_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_14_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_14_clock; // @[Stab.scala 85:60]
  wire  cols_3_14_reset; // @[Stab.scala 85:60]
  wire  cols_3_14_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_14_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_14_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_14_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_14_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_14_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_14_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_3_14_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_14_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_3_14_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_14_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_14_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_14_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_14_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_14_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_14_clock; // @[Stab.scala 85:60]
  wire  cols_4_14_reset; // @[Stab.scala 85:60]
  wire  cols_4_14_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_14_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_14_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_14_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_14_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_14_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_14_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_4_14_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_14_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_4_14_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_14_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_14_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_14_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_14_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_14_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_14_clock; // @[Stab.scala 85:60]
  wire  cols_5_14_reset; // @[Stab.scala 85:60]
  wire  cols_5_14_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_14_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_14_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_14_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_14_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_14_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_14_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_5_14_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_14_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_5_14_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_14_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_14_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_14_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_14_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_14_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_14_clock; // @[Stab.scala 85:60]
  wire  cols_6_14_reset; // @[Stab.scala 85:60]
  wire  cols_6_14_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_14_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_14_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_14_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_14_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_14_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_14_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_6_14_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_14_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_6_14_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_14_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_14_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_14_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_14_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_14_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_14_clock; // @[Stab.scala 85:60]
  wire  cols_7_14_reset; // @[Stab.scala 85:60]
  wire  cols_7_14_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_14_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_14_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_14_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_14_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_14_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_14_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_7_14_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_14_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_7_14_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_14_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_14_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_14_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_14_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_14_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_14_clock; // @[Stab.scala 85:60]
  wire  cols_8_14_reset; // @[Stab.scala 85:60]
  wire  cols_8_14_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_14_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_14_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_14_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_14_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_14_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_14_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_8_14_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_14_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_8_14_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_14_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_14_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_14_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_14_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_14_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_14_clock; // @[Stab.scala 85:60]
  wire  cols_9_14_reset; // @[Stab.scala 85:60]
  wire  cols_9_14_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_14_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_14_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_14_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_14_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_14_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_14_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_9_14_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_14_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_9_14_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_14_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_14_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_14_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_14_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_14_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_14_clock; // @[Stab.scala 85:60]
  wire  cols_10_14_reset; // @[Stab.scala 85:60]
  wire  cols_10_14_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_14_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_14_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_14_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_14_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_14_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_14_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_10_14_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_14_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_10_14_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_14_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_14_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_14_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_14_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_14_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_14_clock; // @[Stab.scala 85:60]
  wire  cols_11_14_reset; // @[Stab.scala 85:60]
  wire  cols_11_14_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_14_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_14_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_14_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_14_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_14_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_14_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_11_14_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_14_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_11_14_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_14_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_14_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_14_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_14_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_14_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_14_clock; // @[Stab.scala 85:60]
  wire  cols_12_14_reset; // @[Stab.scala 85:60]
  wire  cols_12_14_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_14_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_14_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_14_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_14_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_14_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_14_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_12_14_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_14_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_12_14_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_14_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_14_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_14_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_14_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_14_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_14_clock; // @[Stab.scala 85:60]
  wire  cols_13_14_reset; // @[Stab.scala 85:60]
  wire  cols_13_14_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_14_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_14_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_14_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_14_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_14_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_14_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_13_14_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_14_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_13_14_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_14_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_14_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_14_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_14_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_14_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_14_clock; // @[Stab.scala 85:60]
  wire  cols_14_14_reset; // @[Stab.scala 85:60]
  wire  cols_14_14_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_14_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_14_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_14_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_14_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_14_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_14_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_14_14_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_14_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_14_14_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_14_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_14_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_14_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_14_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_14_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_14_clock; // @[Stab.scala 85:60]
  wire  cols_15_14_reset; // @[Stab.scala 85:60]
  wire  cols_15_14_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_14_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_14_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_14_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_14_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_14_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_14_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_15_14_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_14_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_15_14_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_14_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_14_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_14_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_14_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_14_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_15_clock; // @[Stab.scala 85:60]
  wire  cols_0_15_reset; // @[Stab.scala 85:60]
  wire  cols_0_15_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_15_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_15_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_15_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_0_15_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_15_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_0_15_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_0_15_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_15_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_0_15_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_15_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_15_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_0_15_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_0_15_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_0_15_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_15_clock; // @[Stab.scala 85:60]
  wire  cols_1_15_reset; // @[Stab.scala 85:60]
  wire  cols_1_15_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_15_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_15_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_15_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_1_15_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_15_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_1_15_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_1_15_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_15_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_1_15_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_15_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_15_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_1_15_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_1_15_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_1_15_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_15_clock; // @[Stab.scala 85:60]
  wire  cols_2_15_reset; // @[Stab.scala 85:60]
  wire  cols_2_15_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_15_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_15_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_15_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_2_15_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_15_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_2_15_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_2_15_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_15_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_2_15_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_15_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_15_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_2_15_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_2_15_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_2_15_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_15_clock; // @[Stab.scala 85:60]
  wire  cols_3_15_reset; // @[Stab.scala 85:60]
  wire  cols_3_15_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_15_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_15_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_15_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_3_15_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_15_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_3_15_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_3_15_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_15_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_3_15_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_15_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_15_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_3_15_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_3_15_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_3_15_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_15_clock; // @[Stab.scala 85:60]
  wire  cols_4_15_reset; // @[Stab.scala 85:60]
  wire  cols_4_15_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_15_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_15_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_15_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_4_15_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_15_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_4_15_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_4_15_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_15_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_4_15_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_15_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_15_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_4_15_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_4_15_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_4_15_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_15_clock; // @[Stab.scala 85:60]
  wire  cols_5_15_reset; // @[Stab.scala 85:60]
  wire  cols_5_15_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_15_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_15_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_15_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_5_15_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_15_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_5_15_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_5_15_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_15_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_5_15_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_15_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_15_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_5_15_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_5_15_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_5_15_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_15_clock; // @[Stab.scala 85:60]
  wire  cols_6_15_reset; // @[Stab.scala 85:60]
  wire  cols_6_15_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_15_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_15_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_15_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_6_15_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_15_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_6_15_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_6_15_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_15_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_6_15_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_15_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_15_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_6_15_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_6_15_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_6_15_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_15_clock; // @[Stab.scala 85:60]
  wire  cols_7_15_reset; // @[Stab.scala 85:60]
  wire  cols_7_15_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_15_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_15_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_15_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_7_15_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_15_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_7_15_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_7_15_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_15_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_7_15_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_15_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_15_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_7_15_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_7_15_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_7_15_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_15_clock; // @[Stab.scala 85:60]
  wire  cols_8_15_reset; // @[Stab.scala 85:60]
  wire  cols_8_15_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_15_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_15_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_15_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_8_15_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_15_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_8_15_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_8_15_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_15_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_8_15_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_15_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_15_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_8_15_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_8_15_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_8_15_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_15_clock; // @[Stab.scala 85:60]
  wire  cols_9_15_reset; // @[Stab.scala 85:60]
  wire  cols_9_15_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_15_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_15_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_15_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_9_15_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_15_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_9_15_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_9_15_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_15_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_9_15_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_15_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_15_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_9_15_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_9_15_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_9_15_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_15_clock; // @[Stab.scala 85:60]
  wire  cols_10_15_reset; // @[Stab.scala 85:60]
  wire  cols_10_15_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_15_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_15_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_15_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_10_15_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_15_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_10_15_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_10_15_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_15_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_10_15_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_15_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_15_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_10_15_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_10_15_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_10_15_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_15_clock; // @[Stab.scala 85:60]
  wire  cols_11_15_reset; // @[Stab.scala 85:60]
  wire  cols_11_15_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_15_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_15_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_15_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_11_15_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_15_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_11_15_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_11_15_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_15_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_11_15_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_15_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_15_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_11_15_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_11_15_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_11_15_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_15_clock; // @[Stab.scala 85:60]
  wire  cols_12_15_reset; // @[Stab.scala 85:60]
  wire  cols_12_15_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_15_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_15_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_15_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_12_15_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_15_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_12_15_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_12_15_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_15_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_12_15_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_15_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_15_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_12_15_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_12_15_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_12_15_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_15_clock; // @[Stab.scala 85:60]
  wire  cols_13_15_reset; // @[Stab.scala 85:60]
  wire  cols_13_15_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_15_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_15_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_15_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_13_15_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_15_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_13_15_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_13_15_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_15_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_13_15_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_15_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_15_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_13_15_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_13_15_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_13_15_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_15_clock; // @[Stab.scala 85:60]
  wire  cols_14_15_reset; // @[Stab.scala 85:60]
  wire  cols_14_15_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_15_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_15_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_15_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_14_15_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_15_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_14_15_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_14_15_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_15_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_14_15_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_15_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_15_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_14_15_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_14_15_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_14_15_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_15_clock; // @[Stab.scala 85:60]
  wire  cols_15_15_reset; // @[Stab.scala 85:60]
  wire  cols_15_15_io_left_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_15_io_left_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_15_io_left_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_15_io_top_in_ready; // @[Stab.scala 85:60]
  wire  cols_15_15_io_top_in_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_15_io_top_in_bits; // @[Stab.scala 85:60]
  wire  cols_15_15_io_sum_ready; // @[Stab.scala 85:60]
  wire  cols_15_15_io_sum_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_15_io_sum_bits; // @[Stab.scala 85:60]
  wire  cols_15_15_io_right_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_15_io_right_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_15_io_right_out_bits; // @[Stab.scala 85:60]
  wire  cols_15_15_io_bottom_out_ready; // @[Stab.scala 85:60]
  wire  cols_15_15_io_bottom_out_valid; // @[Stab.scala 85:60]
  wire [31:0] cols_15_15_io_bottom_out_bits; // @[Stab.scala 85:60]
  wire  q_clock; // @[Decoupled.scala 361:21]
  wire  q_reset; // @[Decoupled.scala 361:21]
  wire  q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_1_clock; // @[Decoupled.scala 361:21]
  wire  q_1_reset; // @[Decoupled.scala 361:21]
  wire  q_1_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_1_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_1_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_1_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_1_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_1_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_2_clock; // @[Decoupled.scala 361:21]
  wire  q_2_reset; // @[Decoupled.scala 361:21]
  wire  q_2_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_2_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_2_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_2_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_2_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_2_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_3_clock; // @[Decoupled.scala 361:21]
  wire  q_3_reset; // @[Decoupled.scala 361:21]
  wire  q_3_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_3_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_3_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_3_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_3_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_3_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_4_clock; // @[Decoupled.scala 361:21]
  wire  q_4_reset; // @[Decoupled.scala 361:21]
  wire  q_4_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_4_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_4_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_4_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_4_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_4_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_5_clock; // @[Decoupled.scala 361:21]
  wire  q_5_reset; // @[Decoupled.scala 361:21]
  wire  q_5_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_5_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_5_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_5_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_5_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_5_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_6_clock; // @[Decoupled.scala 361:21]
  wire  q_6_reset; // @[Decoupled.scala 361:21]
  wire  q_6_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_6_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_6_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_6_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_6_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_6_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_7_clock; // @[Decoupled.scala 361:21]
  wire  q_7_reset; // @[Decoupled.scala 361:21]
  wire  q_7_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_7_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_7_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_7_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_7_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_7_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_8_clock; // @[Decoupled.scala 361:21]
  wire  q_8_reset; // @[Decoupled.scala 361:21]
  wire  q_8_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_8_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_8_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_8_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_8_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_8_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_9_clock; // @[Decoupled.scala 361:21]
  wire  q_9_reset; // @[Decoupled.scala 361:21]
  wire  q_9_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_9_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_9_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_9_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_9_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_9_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_10_clock; // @[Decoupled.scala 361:21]
  wire  q_10_reset; // @[Decoupled.scala 361:21]
  wire  q_10_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_10_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_10_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_10_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_10_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_10_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_11_clock; // @[Decoupled.scala 361:21]
  wire  q_11_reset; // @[Decoupled.scala 361:21]
  wire  q_11_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_11_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_11_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_11_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_11_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_11_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_12_clock; // @[Decoupled.scala 361:21]
  wire  q_12_reset; // @[Decoupled.scala 361:21]
  wire  q_12_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_12_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_12_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_12_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_12_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_12_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_13_clock; // @[Decoupled.scala 361:21]
  wire  q_13_reset; // @[Decoupled.scala 361:21]
  wire  q_13_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_13_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_13_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_13_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_13_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_13_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_14_clock; // @[Decoupled.scala 361:21]
  wire  q_14_reset; // @[Decoupled.scala 361:21]
  wire  q_14_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_14_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_14_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_14_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_14_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_14_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_15_clock; // @[Decoupled.scala 361:21]
  wire  q_15_reset; // @[Decoupled.scala 361:21]
  wire  q_15_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_15_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_15_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_15_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_15_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_15_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_16_clock; // @[Decoupled.scala 361:21]
  wire  q_16_reset; // @[Decoupled.scala 361:21]
  wire  q_16_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_16_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_16_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_16_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_16_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_16_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_17_clock; // @[Decoupled.scala 361:21]
  wire  q_17_reset; // @[Decoupled.scala 361:21]
  wire  q_17_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_17_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_17_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_17_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_17_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_17_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_18_clock; // @[Decoupled.scala 361:21]
  wire  q_18_reset; // @[Decoupled.scala 361:21]
  wire  q_18_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_18_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_18_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_18_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_18_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_18_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_19_clock; // @[Decoupled.scala 361:21]
  wire  q_19_reset; // @[Decoupled.scala 361:21]
  wire  q_19_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_19_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_19_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_19_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_19_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_19_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_20_clock; // @[Decoupled.scala 361:21]
  wire  q_20_reset; // @[Decoupled.scala 361:21]
  wire  q_20_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_20_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_20_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_20_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_20_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_20_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_21_clock; // @[Decoupled.scala 361:21]
  wire  q_21_reset; // @[Decoupled.scala 361:21]
  wire  q_21_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_21_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_21_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_21_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_21_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_21_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_22_clock; // @[Decoupled.scala 361:21]
  wire  q_22_reset; // @[Decoupled.scala 361:21]
  wire  q_22_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_22_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_22_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_22_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_22_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_22_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_23_clock; // @[Decoupled.scala 361:21]
  wire  q_23_reset; // @[Decoupled.scala 361:21]
  wire  q_23_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_23_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_23_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_23_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_23_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_23_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_24_clock; // @[Decoupled.scala 361:21]
  wire  q_24_reset; // @[Decoupled.scala 361:21]
  wire  q_24_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_24_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_24_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_24_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_24_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_24_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_25_clock; // @[Decoupled.scala 361:21]
  wire  q_25_reset; // @[Decoupled.scala 361:21]
  wire  q_25_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_25_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_25_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_25_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_25_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_25_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_26_clock; // @[Decoupled.scala 361:21]
  wire  q_26_reset; // @[Decoupled.scala 361:21]
  wire  q_26_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_26_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_26_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_26_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_26_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_26_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_27_clock; // @[Decoupled.scala 361:21]
  wire  q_27_reset; // @[Decoupled.scala 361:21]
  wire  q_27_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_27_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_27_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_27_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_27_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_27_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_28_clock; // @[Decoupled.scala 361:21]
  wire  q_28_reset; // @[Decoupled.scala 361:21]
  wire  q_28_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_28_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_28_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_28_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_28_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_28_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_29_clock; // @[Decoupled.scala 361:21]
  wire  q_29_reset; // @[Decoupled.scala 361:21]
  wire  q_29_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_29_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_29_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_29_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_29_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_29_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_30_clock; // @[Decoupled.scala 361:21]
  wire  q_30_reset; // @[Decoupled.scala 361:21]
  wire  q_30_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_30_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_30_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_30_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_30_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_30_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_31_clock; // @[Decoupled.scala 361:21]
  wire  q_31_reset; // @[Decoupled.scala 361:21]
  wire  q_31_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_31_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_31_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_31_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_31_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_31_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_32_clock; // @[Decoupled.scala 361:21]
  wire  q_32_reset; // @[Decoupled.scala 361:21]
  wire  q_32_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_32_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_32_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_32_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_32_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_32_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_33_clock; // @[Decoupled.scala 361:21]
  wire  q_33_reset; // @[Decoupled.scala 361:21]
  wire  q_33_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_33_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_33_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_33_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_33_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_33_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_34_clock; // @[Decoupled.scala 361:21]
  wire  q_34_reset; // @[Decoupled.scala 361:21]
  wire  q_34_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_34_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_34_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_34_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_34_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_34_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_35_clock; // @[Decoupled.scala 361:21]
  wire  q_35_reset; // @[Decoupled.scala 361:21]
  wire  q_35_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_35_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_35_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_35_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_35_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_35_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_36_clock; // @[Decoupled.scala 361:21]
  wire  q_36_reset; // @[Decoupled.scala 361:21]
  wire  q_36_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_36_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_36_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_36_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_36_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_36_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_37_clock; // @[Decoupled.scala 361:21]
  wire  q_37_reset; // @[Decoupled.scala 361:21]
  wire  q_37_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_37_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_37_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_37_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_37_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_37_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_38_clock; // @[Decoupled.scala 361:21]
  wire  q_38_reset; // @[Decoupled.scala 361:21]
  wire  q_38_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_38_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_38_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_38_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_38_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_38_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_39_clock; // @[Decoupled.scala 361:21]
  wire  q_39_reset; // @[Decoupled.scala 361:21]
  wire  q_39_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_39_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_39_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_39_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_39_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_39_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_40_clock; // @[Decoupled.scala 361:21]
  wire  q_40_reset; // @[Decoupled.scala 361:21]
  wire  q_40_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_40_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_40_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_40_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_40_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_40_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_41_clock; // @[Decoupled.scala 361:21]
  wire  q_41_reset; // @[Decoupled.scala 361:21]
  wire  q_41_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_41_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_41_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_41_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_41_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_41_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_42_clock; // @[Decoupled.scala 361:21]
  wire  q_42_reset; // @[Decoupled.scala 361:21]
  wire  q_42_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_42_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_42_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_42_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_42_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_42_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_43_clock; // @[Decoupled.scala 361:21]
  wire  q_43_reset; // @[Decoupled.scala 361:21]
  wire  q_43_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_43_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_43_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_43_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_43_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_43_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_44_clock; // @[Decoupled.scala 361:21]
  wire  q_44_reset; // @[Decoupled.scala 361:21]
  wire  q_44_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_44_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_44_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_44_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_44_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_44_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_45_clock; // @[Decoupled.scala 361:21]
  wire  q_45_reset; // @[Decoupled.scala 361:21]
  wire  q_45_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_45_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_45_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_45_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_45_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_45_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_46_clock; // @[Decoupled.scala 361:21]
  wire  q_46_reset; // @[Decoupled.scala 361:21]
  wire  q_46_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_46_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_46_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_46_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_46_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_46_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_47_clock; // @[Decoupled.scala 361:21]
  wire  q_47_reset; // @[Decoupled.scala 361:21]
  wire  q_47_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_47_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_47_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_47_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_47_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_47_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_48_clock; // @[Decoupled.scala 361:21]
  wire  q_48_reset; // @[Decoupled.scala 361:21]
  wire  q_48_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_48_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_48_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_48_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_48_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_48_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_49_clock; // @[Decoupled.scala 361:21]
  wire  q_49_reset; // @[Decoupled.scala 361:21]
  wire  q_49_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_49_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_49_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_49_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_49_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_49_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_50_clock; // @[Decoupled.scala 361:21]
  wire  q_50_reset; // @[Decoupled.scala 361:21]
  wire  q_50_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_50_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_50_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_50_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_50_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_50_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_51_clock; // @[Decoupled.scala 361:21]
  wire  q_51_reset; // @[Decoupled.scala 361:21]
  wire  q_51_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_51_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_51_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_51_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_51_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_51_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_52_clock; // @[Decoupled.scala 361:21]
  wire  q_52_reset; // @[Decoupled.scala 361:21]
  wire  q_52_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_52_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_52_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_52_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_52_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_52_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_53_clock; // @[Decoupled.scala 361:21]
  wire  q_53_reset; // @[Decoupled.scala 361:21]
  wire  q_53_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_53_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_53_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_53_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_53_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_53_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_54_clock; // @[Decoupled.scala 361:21]
  wire  q_54_reset; // @[Decoupled.scala 361:21]
  wire  q_54_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_54_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_54_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_54_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_54_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_54_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_55_clock; // @[Decoupled.scala 361:21]
  wire  q_55_reset; // @[Decoupled.scala 361:21]
  wire  q_55_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_55_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_55_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_55_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_55_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_55_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_56_clock; // @[Decoupled.scala 361:21]
  wire  q_56_reset; // @[Decoupled.scala 361:21]
  wire  q_56_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_56_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_56_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_56_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_56_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_56_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_57_clock; // @[Decoupled.scala 361:21]
  wire  q_57_reset; // @[Decoupled.scala 361:21]
  wire  q_57_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_57_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_57_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_57_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_57_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_57_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_58_clock; // @[Decoupled.scala 361:21]
  wire  q_58_reset; // @[Decoupled.scala 361:21]
  wire  q_58_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_58_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_58_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_58_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_58_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_58_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_59_clock; // @[Decoupled.scala 361:21]
  wire  q_59_reset; // @[Decoupled.scala 361:21]
  wire  q_59_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_59_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_59_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_59_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_59_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_59_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_60_clock; // @[Decoupled.scala 361:21]
  wire  q_60_reset; // @[Decoupled.scala 361:21]
  wire  q_60_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_60_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_60_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_60_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_60_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_60_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_61_clock; // @[Decoupled.scala 361:21]
  wire  q_61_reset; // @[Decoupled.scala 361:21]
  wire  q_61_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_61_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_61_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_61_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_61_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_61_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_62_clock; // @[Decoupled.scala 361:21]
  wire  q_62_reset; // @[Decoupled.scala 361:21]
  wire  q_62_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_62_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_62_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_62_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_62_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_62_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_63_clock; // @[Decoupled.scala 361:21]
  wire  q_63_reset; // @[Decoupled.scala 361:21]
  wire  q_63_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_63_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_63_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_63_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_63_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_63_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_64_clock; // @[Decoupled.scala 361:21]
  wire  q_64_reset; // @[Decoupled.scala 361:21]
  wire  q_64_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_64_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_64_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_64_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_64_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_64_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_65_clock; // @[Decoupled.scala 361:21]
  wire  q_65_reset; // @[Decoupled.scala 361:21]
  wire  q_65_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_65_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_65_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_65_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_65_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_65_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_66_clock; // @[Decoupled.scala 361:21]
  wire  q_66_reset; // @[Decoupled.scala 361:21]
  wire  q_66_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_66_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_66_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_66_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_66_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_66_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_67_clock; // @[Decoupled.scala 361:21]
  wire  q_67_reset; // @[Decoupled.scala 361:21]
  wire  q_67_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_67_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_67_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_67_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_67_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_67_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_68_clock; // @[Decoupled.scala 361:21]
  wire  q_68_reset; // @[Decoupled.scala 361:21]
  wire  q_68_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_68_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_68_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_68_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_68_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_68_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_69_clock; // @[Decoupled.scala 361:21]
  wire  q_69_reset; // @[Decoupled.scala 361:21]
  wire  q_69_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_69_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_69_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_69_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_69_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_69_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_70_clock; // @[Decoupled.scala 361:21]
  wire  q_70_reset; // @[Decoupled.scala 361:21]
  wire  q_70_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_70_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_70_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_70_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_70_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_70_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_71_clock; // @[Decoupled.scala 361:21]
  wire  q_71_reset; // @[Decoupled.scala 361:21]
  wire  q_71_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_71_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_71_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_71_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_71_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_71_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_72_clock; // @[Decoupled.scala 361:21]
  wire  q_72_reset; // @[Decoupled.scala 361:21]
  wire  q_72_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_72_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_72_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_72_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_72_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_72_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_73_clock; // @[Decoupled.scala 361:21]
  wire  q_73_reset; // @[Decoupled.scala 361:21]
  wire  q_73_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_73_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_73_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_73_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_73_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_73_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_74_clock; // @[Decoupled.scala 361:21]
  wire  q_74_reset; // @[Decoupled.scala 361:21]
  wire  q_74_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_74_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_74_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_74_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_74_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_74_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_75_clock; // @[Decoupled.scala 361:21]
  wire  q_75_reset; // @[Decoupled.scala 361:21]
  wire  q_75_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_75_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_75_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_75_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_75_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_75_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_76_clock; // @[Decoupled.scala 361:21]
  wire  q_76_reset; // @[Decoupled.scala 361:21]
  wire  q_76_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_76_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_76_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_76_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_76_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_76_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_77_clock; // @[Decoupled.scala 361:21]
  wire  q_77_reset; // @[Decoupled.scala 361:21]
  wire  q_77_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_77_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_77_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_77_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_77_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_77_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_78_clock; // @[Decoupled.scala 361:21]
  wire  q_78_reset; // @[Decoupled.scala 361:21]
  wire  q_78_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_78_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_78_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_78_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_78_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_78_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_79_clock; // @[Decoupled.scala 361:21]
  wire  q_79_reset; // @[Decoupled.scala 361:21]
  wire  q_79_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_79_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_79_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_79_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_79_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_79_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_80_clock; // @[Decoupled.scala 361:21]
  wire  q_80_reset; // @[Decoupled.scala 361:21]
  wire  q_80_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_80_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_80_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_80_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_80_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_80_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_81_clock; // @[Decoupled.scala 361:21]
  wire  q_81_reset; // @[Decoupled.scala 361:21]
  wire  q_81_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_81_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_81_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_81_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_81_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_81_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_82_clock; // @[Decoupled.scala 361:21]
  wire  q_82_reset; // @[Decoupled.scala 361:21]
  wire  q_82_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_82_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_82_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_82_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_82_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_82_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_83_clock; // @[Decoupled.scala 361:21]
  wire  q_83_reset; // @[Decoupled.scala 361:21]
  wire  q_83_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_83_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_83_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_83_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_83_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_83_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_84_clock; // @[Decoupled.scala 361:21]
  wire  q_84_reset; // @[Decoupled.scala 361:21]
  wire  q_84_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_84_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_84_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_84_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_84_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_84_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_85_clock; // @[Decoupled.scala 361:21]
  wire  q_85_reset; // @[Decoupled.scala 361:21]
  wire  q_85_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_85_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_85_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_85_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_85_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_85_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_86_clock; // @[Decoupled.scala 361:21]
  wire  q_86_reset; // @[Decoupled.scala 361:21]
  wire  q_86_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_86_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_86_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_86_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_86_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_86_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_87_clock; // @[Decoupled.scala 361:21]
  wire  q_87_reset; // @[Decoupled.scala 361:21]
  wire  q_87_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_87_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_87_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_87_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_87_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_87_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_88_clock; // @[Decoupled.scala 361:21]
  wire  q_88_reset; // @[Decoupled.scala 361:21]
  wire  q_88_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_88_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_88_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_88_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_88_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_88_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_89_clock; // @[Decoupled.scala 361:21]
  wire  q_89_reset; // @[Decoupled.scala 361:21]
  wire  q_89_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_89_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_89_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_89_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_89_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_89_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_90_clock; // @[Decoupled.scala 361:21]
  wire  q_90_reset; // @[Decoupled.scala 361:21]
  wire  q_90_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_90_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_90_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_90_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_90_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_90_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_91_clock; // @[Decoupled.scala 361:21]
  wire  q_91_reset; // @[Decoupled.scala 361:21]
  wire  q_91_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_91_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_91_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_91_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_91_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_91_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_92_clock; // @[Decoupled.scala 361:21]
  wire  q_92_reset; // @[Decoupled.scala 361:21]
  wire  q_92_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_92_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_92_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_92_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_92_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_92_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_93_clock; // @[Decoupled.scala 361:21]
  wire  q_93_reset; // @[Decoupled.scala 361:21]
  wire  q_93_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_93_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_93_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_93_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_93_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_93_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_94_clock; // @[Decoupled.scala 361:21]
  wire  q_94_reset; // @[Decoupled.scala 361:21]
  wire  q_94_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_94_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_94_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_94_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_94_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_94_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_95_clock; // @[Decoupled.scala 361:21]
  wire  q_95_reset; // @[Decoupled.scala 361:21]
  wire  q_95_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_95_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_95_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_95_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_95_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_95_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_96_clock; // @[Decoupled.scala 361:21]
  wire  q_96_reset; // @[Decoupled.scala 361:21]
  wire  q_96_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_96_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_96_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_96_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_96_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_96_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_97_clock; // @[Decoupled.scala 361:21]
  wire  q_97_reset; // @[Decoupled.scala 361:21]
  wire  q_97_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_97_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_97_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_97_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_97_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_97_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_98_clock; // @[Decoupled.scala 361:21]
  wire  q_98_reset; // @[Decoupled.scala 361:21]
  wire  q_98_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_98_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_98_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_98_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_98_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_98_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_99_clock; // @[Decoupled.scala 361:21]
  wire  q_99_reset; // @[Decoupled.scala 361:21]
  wire  q_99_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_99_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_99_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_99_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_99_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_99_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_100_clock; // @[Decoupled.scala 361:21]
  wire  q_100_reset; // @[Decoupled.scala 361:21]
  wire  q_100_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_100_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_100_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_100_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_100_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_100_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_101_clock; // @[Decoupled.scala 361:21]
  wire  q_101_reset; // @[Decoupled.scala 361:21]
  wire  q_101_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_101_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_101_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_101_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_101_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_101_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_102_clock; // @[Decoupled.scala 361:21]
  wire  q_102_reset; // @[Decoupled.scala 361:21]
  wire  q_102_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_102_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_102_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_102_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_102_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_102_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_103_clock; // @[Decoupled.scala 361:21]
  wire  q_103_reset; // @[Decoupled.scala 361:21]
  wire  q_103_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_103_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_103_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_103_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_103_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_103_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_104_clock; // @[Decoupled.scala 361:21]
  wire  q_104_reset; // @[Decoupled.scala 361:21]
  wire  q_104_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_104_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_104_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_104_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_104_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_104_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_105_clock; // @[Decoupled.scala 361:21]
  wire  q_105_reset; // @[Decoupled.scala 361:21]
  wire  q_105_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_105_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_105_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_105_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_105_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_105_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_106_clock; // @[Decoupled.scala 361:21]
  wire  q_106_reset; // @[Decoupled.scala 361:21]
  wire  q_106_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_106_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_106_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_106_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_106_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_106_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_107_clock; // @[Decoupled.scala 361:21]
  wire  q_107_reset; // @[Decoupled.scala 361:21]
  wire  q_107_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_107_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_107_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_107_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_107_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_107_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_108_clock; // @[Decoupled.scala 361:21]
  wire  q_108_reset; // @[Decoupled.scala 361:21]
  wire  q_108_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_108_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_108_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_108_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_108_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_108_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_109_clock; // @[Decoupled.scala 361:21]
  wire  q_109_reset; // @[Decoupled.scala 361:21]
  wire  q_109_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_109_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_109_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_109_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_109_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_109_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_110_clock; // @[Decoupled.scala 361:21]
  wire  q_110_reset; // @[Decoupled.scala 361:21]
  wire  q_110_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_110_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_110_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_110_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_110_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_110_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_111_clock; // @[Decoupled.scala 361:21]
  wire  q_111_reset; // @[Decoupled.scala 361:21]
  wire  q_111_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_111_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_111_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_111_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_111_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_111_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_112_clock; // @[Decoupled.scala 361:21]
  wire  q_112_reset; // @[Decoupled.scala 361:21]
  wire  q_112_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_112_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_112_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_112_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_112_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_112_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_113_clock; // @[Decoupled.scala 361:21]
  wire  q_113_reset; // @[Decoupled.scala 361:21]
  wire  q_113_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_113_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_113_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_113_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_113_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_113_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_114_clock; // @[Decoupled.scala 361:21]
  wire  q_114_reset; // @[Decoupled.scala 361:21]
  wire  q_114_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_114_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_114_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_114_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_114_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_114_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_115_clock; // @[Decoupled.scala 361:21]
  wire  q_115_reset; // @[Decoupled.scala 361:21]
  wire  q_115_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_115_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_115_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_115_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_115_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_115_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_116_clock; // @[Decoupled.scala 361:21]
  wire  q_116_reset; // @[Decoupled.scala 361:21]
  wire  q_116_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_116_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_116_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_116_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_116_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_116_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_117_clock; // @[Decoupled.scala 361:21]
  wire  q_117_reset; // @[Decoupled.scala 361:21]
  wire  q_117_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_117_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_117_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_117_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_117_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_117_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_118_clock; // @[Decoupled.scala 361:21]
  wire  q_118_reset; // @[Decoupled.scala 361:21]
  wire  q_118_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_118_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_118_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_118_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_118_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_118_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_119_clock; // @[Decoupled.scala 361:21]
  wire  q_119_reset; // @[Decoupled.scala 361:21]
  wire  q_119_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_119_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_119_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_119_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_119_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_119_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_120_clock; // @[Decoupled.scala 361:21]
  wire  q_120_reset; // @[Decoupled.scala 361:21]
  wire  q_120_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_120_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_120_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_120_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_120_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_120_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_121_clock; // @[Decoupled.scala 361:21]
  wire  q_121_reset; // @[Decoupled.scala 361:21]
  wire  q_121_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_121_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_121_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_121_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_121_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_121_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_122_clock; // @[Decoupled.scala 361:21]
  wire  q_122_reset; // @[Decoupled.scala 361:21]
  wire  q_122_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_122_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_122_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_122_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_122_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_122_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_123_clock; // @[Decoupled.scala 361:21]
  wire  q_123_reset; // @[Decoupled.scala 361:21]
  wire  q_123_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_123_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_123_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_123_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_123_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_123_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_124_clock; // @[Decoupled.scala 361:21]
  wire  q_124_reset; // @[Decoupled.scala 361:21]
  wire  q_124_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_124_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_124_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_124_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_124_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_124_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_125_clock; // @[Decoupled.scala 361:21]
  wire  q_125_reset; // @[Decoupled.scala 361:21]
  wire  q_125_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_125_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_125_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_125_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_125_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_125_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_126_clock; // @[Decoupled.scala 361:21]
  wire  q_126_reset; // @[Decoupled.scala 361:21]
  wire  q_126_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_126_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_126_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_126_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_126_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_126_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_127_clock; // @[Decoupled.scala 361:21]
  wire  q_127_reset; // @[Decoupled.scala 361:21]
  wire  q_127_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_127_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_127_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_127_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_127_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_127_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_128_clock; // @[Decoupled.scala 361:21]
  wire  q_128_reset; // @[Decoupled.scala 361:21]
  wire  q_128_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_128_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_128_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_128_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_128_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_128_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_129_clock; // @[Decoupled.scala 361:21]
  wire  q_129_reset; // @[Decoupled.scala 361:21]
  wire  q_129_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_129_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_129_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_129_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_129_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_129_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_130_clock; // @[Decoupled.scala 361:21]
  wire  q_130_reset; // @[Decoupled.scala 361:21]
  wire  q_130_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_130_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_130_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_130_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_130_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_130_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_131_clock; // @[Decoupled.scala 361:21]
  wire  q_131_reset; // @[Decoupled.scala 361:21]
  wire  q_131_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_131_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_131_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_131_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_131_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_131_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_132_clock; // @[Decoupled.scala 361:21]
  wire  q_132_reset; // @[Decoupled.scala 361:21]
  wire  q_132_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_132_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_132_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_132_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_132_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_132_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_133_clock; // @[Decoupled.scala 361:21]
  wire  q_133_reset; // @[Decoupled.scala 361:21]
  wire  q_133_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_133_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_133_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_133_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_133_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_133_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_134_clock; // @[Decoupled.scala 361:21]
  wire  q_134_reset; // @[Decoupled.scala 361:21]
  wire  q_134_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_134_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_134_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_134_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_134_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_134_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_135_clock; // @[Decoupled.scala 361:21]
  wire  q_135_reset; // @[Decoupled.scala 361:21]
  wire  q_135_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_135_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_135_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_135_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_135_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_135_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_136_clock; // @[Decoupled.scala 361:21]
  wire  q_136_reset; // @[Decoupled.scala 361:21]
  wire  q_136_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_136_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_136_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_136_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_136_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_136_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_137_clock; // @[Decoupled.scala 361:21]
  wire  q_137_reset; // @[Decoupled.scala 361:21]
  wire  q_137_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_137_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_137_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_137_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_137_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_137_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_138_clock; // @[Decoupled.scala 361:21]
  wire  q_138_reset; // @[Decoupled.scala 361:21]
  wire  q_138_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_138_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_138_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_138_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_138_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_138_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_139_clock; // @[Decoupled.scala 361:21]
  wire  q_139_reset; // @[Decoupled.scala 361:21]
  wire  q_139_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_139_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_139_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_139_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_139_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_139_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_140_clock; // @[Decoupled.scala 361:21]
  wire  q_140_reset; // @[Decoupled.scala 361:21]
  wire  q_140_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_140_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_140_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_140_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_140_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_140_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_141_clock; // @[Decoupled.scala 361:21]
  wire  q_141_reset; // @[Decoupled.scala 361:21]
  wire  q_141_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_141_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_141_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_141_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_141_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_141_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_142_clock; // @[Decoupled.scala 361:21]
  wire  q_142_reset; // @[Decoupled.scala 361:21]
  wire  q_142_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_142_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_142_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_142_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_142_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_142_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_143_clock; // @[Decoupled.scala 361:21]
  wire  q_143_reset; // @[Decoupled.scala 361:21]
  wire  q_143_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_143_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_143_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_143_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_143_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_143_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_144_clock; // @[Decoupled.scala 361:21]
  wire  q_144_reset; // @[Decoupled.scala 361:21]
  wire  q_144_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_144_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_144_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_144_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_144_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_144_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_145_clock; // @[Decoupled.scala 361:21]
  wire  q_145_reset; // @[Decoupled.scala 361:21]
  wire  q_145_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_145_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_145_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_145_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_145_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_145_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_146_clock; // @[Decoupled.scala 361:21]
  wire  q_146_reset; // @[Decoupled.scala 361:21]
  wire  q_146_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_146_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_146_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_146_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_146_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_146_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_147_clock; // @[Decoupled.scala 361:21]
  wire  q_147_reset; // @[Decoupled.scala 361:21]
  wire  q_147_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_147_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_147_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_147_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_147_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_147_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_148_clock; // @[Decoupled.scala 361:21]
  wire  q_148_reset; // @[Decoupled.scala 361:21]
  wire  q_148_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_148_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_148_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_148_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_148_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_148_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_149_clock; // @[Decoupled.scala 361:21]
  wire  q_149_reset; // @[Decoupled.scala 361:21]
  wire  q_149_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_149_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_149_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_149_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_149_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_149_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_150_clock; // @[Decoupled.scala 361:21]
  wire  q_150_reset; // @[Decoupled.scala 361:21]
  wire  q_150_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_150_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_150_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_150_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_150_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_150_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_151_clock; // @[Decoupled.scala 361:21]
  wire  q_151_reset; // @[Decoupled.scala 361:21]
  wire  q_151_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_151_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_151_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_151_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_151_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_151_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_152_clock; // @[Decoupled.scala 361:21]
  wire  q_152_reset; // @[Decoupled.scala 361:21]
  wire  q_152_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_152_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_152_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_152_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_152_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_152_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_153_clock; // @[Decoupled.scala 361:21]
  wire  q_153_reset; // @[Decoupled.scala 361:21]
  wire  q_153_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_153_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_153_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_153_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_153_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_153_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_154_clock; // @[Decoupled.scala 361:21]
  wire  q_154_reset; // @[Decoupled.scala 361:21]
  wire  q_154_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_154_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_154_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_154_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_154_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_154_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_155_clock; // @[Decoupled.scala 361:21]
  wire  q_155_reset; // @[Decoupled.scala 361:21]
  wire  q_155_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_155_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_155_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_155_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_155_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_155_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_156_clock; // @[Decoupled.scala 361:21]
  wire  q_156_reset; // @[Decoupled.scala 361:21]
  wire  q_156_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_156_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_156_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_156_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_156_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_156_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_157_clock; // @[Decoupled.scala 361:21]
  wire  q_157_reset; // @[Decoupled.scala 361:21]
  wire  q_157_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_157_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_157_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_157_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_157_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_157_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_158_clock; // @[Decoupled.scala 361:21]
  wire  q_158_reset; // @[Decoupled.scala 361:21]
  wire  q_158_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_158_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_158_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_158_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_158_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_158_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_159_clock; // @[Decoupled.scala 361:21]
  wire  q_159_reset; // @[Decoupled.scala 361:21]
  wire  q_159_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_159_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_159_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_159_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_159_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_159_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_160_clock; // @[Decoupled.scala 361:21]
  wire  q_160_reset; // @[Decoupled.scala 361:21]
  wire  q_160_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_160_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_160_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_160_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_160_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_160_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_161_clock; // @[Decoupled.scala 361:21]
  wire  q_161_reset; // @[Decoupled.scala 361:21]
  wire  q_161_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_161_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_161_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_161_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_161_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_161_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_162_clock; // @[Decoupled.scala 361:21]
  wire  q_162_reset; // @[Decoupled.scala 361:21]
  wire  q_162_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_162_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_162_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_162_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_162_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_162_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_163_clock; // @[Decoupled.scala 361:21]
  wire  q_163_reset; // @[Decoupled.scala 361:21]
  wire  q_163_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_163_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_163_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_163_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_163_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_163_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_164_clock; // @[Decoupled.scala 361:21]
  wire  q_164_reset; // @[Decoupled.scala 361:21]
  wire  q_164_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_164_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_164_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_164_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_164_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_164_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_165_clock; // @[Decoupled.scala 361:21]
  wire  q_165_reset; // @[Decoupled.scala 361:21]
  wire  q_165_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_165_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_165_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_165_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_165_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_165_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_166_clock; // @[Decoupled.scala 361:21]
  wire  q_166_reset; // @[Decoupled.scala 361:21]
  wire  q_166_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_166_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_166_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_166_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_166_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_166_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_167_clock; // @[Decoupled.scala 361:21]
  wire  q_167_reset; // @[Decoupled.scala 361:21]
  wire  q_167_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_167_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_167_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_167_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_167_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_167_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_168_clock; // @[Decoupled.scala 361:21]
  wire  q_168_reset; // @[Decoupled.scala 361:21]
  wire  q_168_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_168_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_168_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_168_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_168_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_168_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_169_clock; // @[Decoupled.scala 361:21]
  wire  q_169_reset; // @[Decoupled.scala 361:21]
  wire  q_169_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_169_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_169_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_169_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_169_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_169_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_170_clock; // @[Decoupled.scala 361:21]
  wire  q_170_reset; // @[Decoupled.scala 361:21]
  wire  q_170_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_170_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_170_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_170_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_170_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_170_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_171_clock; // @[Decoupled.scala 361:21]
  wire  q_171_reset; // @[Decoupled.scala 361:21]
  wire  q_171_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_171_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_171_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_171_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_171_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_171_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_172_clock; // @[Decoupled.scala 361:21]
  wire  q_172_reset; // @[Decoupled.scala 361:21]
  wire  q_172_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_172_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_172_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_172_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_172_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_172_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_173_clock; // @[Decoupled.scala 361:21]
  wire  q_173_reset; // @[Decoupled.scala 361:21]
  wire  q_173_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_173_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_173_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_173_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_173_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_173_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_174_clock; // @[Decoupled.scala 361:21]
  wire  q_174_reset; // @[Decoupled.scala 361:21]
  wire  q_174_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_174_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_174_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_174_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_174_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_174_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_175_clock; // @[Decoupled.scala 361:21]
  wire  q_175_reset; // @[Decoupled.scala 361:21]
  wire  q_175_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_175_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_175_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_175_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_175_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_175_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_176_clock; // @[Decoupled.scala 361:21]
  wire  q_176_reset; // @[Decoupled.scala 361:21]
  wire  q_176_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_176_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_176_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_176_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_176_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_176_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_177_clock; // @[Decoupled.scala 361:21]
  wire  q_177_reset; // @[Decoupled.scala 361:21]
  wire  q_177_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_177_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_177_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_177_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_177_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_177_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_178_clock; // @[Decoupled.scala 361:21]
  wire  q_178_reset; // @[Decoupled.scala 361:21]
  wire  q_178_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_178_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_178_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_178_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_178_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_178_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_179_clock; // @[Decoupled.scala 361:21]
  wire  q_179_reset; // @[Decoupled.scala 361:21]
  wire  q_179_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_179_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_179_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_179_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_179_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_179_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_180_clock; // @[Decoupled.scala 361:21]
  wire  q_180_reset; // @[Decoupled.scala 361:21]
  wire  q_180_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_180_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_180_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_180_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_180_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_180_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_181_clock; // @[Decoupled.scala 361:21]
  wire  q_181_reset; // @[Decoupled.scala 361:21]
  wire  q_181_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_181_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_181_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_181_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_181_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_181_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_182_clock; // @[Decoupled.scala 361:21]
  wire  q_182_reset; // @[Decoupled.scala 361:21]
  wire  q_182_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_182_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_182_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_182_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_182_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_182_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_183_clock; // @[Decoupled.scala 361:21]
  wire  q_183_reset; // @[Decoupled.scala 361:21]
  wire  q_183_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_183_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_183_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_183_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_183_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_183_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_184_clock; // @[Decoupled.scala 361:21]
  wire  q_184_reset; // @[Decoupled.scala 361:21]
  wire  q_184_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_184_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_184_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_184_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_184_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_184_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_185_clock; // @[Decoupled.scala 361:21]
  wire  q_185_reset; // @[Decoupled.scala 361:21]
  wire  q_185_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_185_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_185_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_185_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_185_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_185_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_186_clock; // @[Decoupled.scala 361:21]
  wire  q_186_reset; // @[Decoupled.scala 361:21]
  wire  q_186_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_186_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_186_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_186_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_186_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_186_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_187_clock; // @[Decoupled.scala 361:21]
  wire  q_187_reset; // @[Decoupled.scala 361:21]
  wire  q_187_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_187_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_187_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_187_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_187_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_187_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_188_clock; // @[Decoupled.scala 361:21]
  wire  q_188_reset; // @[Decoupled.scala 361:21]
  wire  q_188_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_188_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_188_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_188_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_188_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_188_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_189_clock; // @[Decoupled.scala 361:21]
  wire  q_189_reset; // @[Decoupled.scala 361:21]
  wire  q_189_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_189_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_189_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_189_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_189_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_189_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_190_clock; // @[Decoupled.scala 361:21]
  wire  q_190_reset; // @[Decoupled.scala 361:21]
  wire  q_190_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_190_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_190_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_190_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_190_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_190_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_191_clock; // @[Decoupled.scala 361:21]
  wire  q_191_reset; // @[Decoupled.scala 361:21]
  wire  q_191_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_191_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_191_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_191_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_191_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_191_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_192_clock; // @[Decoupled.scala 361:21]
  wire  q_192_reset; // @[Decoupled.scala 361:21]
  wire  q_192_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_192_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_192_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_192_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_192_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_192_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_193_clock; // @[Decoupled.scala 361:21]
  wire  q_193_reset; // @[Decoupled.scala 361:21]
  wire  q_193_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_193_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_193_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_193_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_193_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_193_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_194_clock; // @[Decoupled.scala 361:21]
  wire  q_194_reset; // @[Decoupled.scala 361:21]
  wire  q_194_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_194_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_194_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_194_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_194_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_194_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_195_clock; // @[Decoupled.scala 361:21]
  wire  q_195_reset; // @[Decoupled.scala 361:21]
  wire  q_195_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_195_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_195_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_195_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_195_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_195_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_196_clock; // @[Decoupled.scala 361:21]
  wire  q_196_reset; // @[Decoupled.scala 361:21]
  wire  q_196_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_196_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_196_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_196_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_196_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_196_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_197_clock; // @[Decoupled.scala 361:21]
  wire  q_197_reset; // @[Decoupled.scala 361:21]
  wire  q_197_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_197_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_197_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_197_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_197_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_197_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_198_clock; // @[Decoupled.scala 361:21]
  wire  q_198_reset; // @[Decoupled.scala 361:21]
  wire  q_198_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_198_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_198_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_198_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_198_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_198_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_199_clock; // @[Decoupled.scala 361:21]
  wire  q_199_reset; // @[Decoupled.scala 361:21]
  wire  q_199_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_199_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_199_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_199_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_199_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_199_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_200_clock; // @[Decoupled.scala 361:21]
  wire  q_200_reset; // @[Decoupled.scala 361:21]
  wire  q_200_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_200_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_200_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_200_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_200_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_200_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_201_clock; // @[Decoupled.scala 361:21]
  wire  q_201_reset; // @[Decoupled.scala 361:21]
  wire  q_201_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_201_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_201_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_201_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_201_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_201_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_202_clock; // @[Decoupled.scala 361:21]
  wire  q_202_reset; // @[Decoupled.scala 361:21]
  wire  q_202_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_202_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_202_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_202_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_202_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_202_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_203_clock; // @[Decoupled.scala 361:21]
  wire  q_203_reset; // @[Decoupled.scala 361:21]
  wire  q_203_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_203_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_203_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_203_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_203_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_203_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_204_clock; // @[Decoupled.scala 361:21]
  wire  q_204_reset; // @[Decoupled.scala 361:21]
  wire  q_204_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_204_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_204_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_204_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_204_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_204_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_205_clock; // @[Decoupled.scala 361:21]
  wire  q_205_reset; // @[Decoupled.scala 361:21]
  wire  q_205_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_205_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_205_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_205_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_205_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_205_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_206_clock; // @[Decoupled.scala 361:21]
  wire  q_206_reset; // @[Decoupled.scala 361:21]
  wire  q_206_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_206_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_206_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_206_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_206_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_206_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_207_clock; // @[Decoupled.scala 361:21]
  wire  q_207_reset; // @[Decoupled.scala 361:21]
  wire  q_207_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_207_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_207_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_207_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_207_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_207_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_208_clock; // @[Decoupled.scala 361:21]
  wire  q_208_reset; // @[Decoupled.scala 361:21]
  wire  q_208_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_208_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_208_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_208_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_208_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_208_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_209_clock; // @[Decoupled.scala 361:21]
  wire  q_209_reset; // @[Decoupled.scala 361:21]
  wire  q_209_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_209_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_209_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_209_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_209_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_209_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_210_clock; // @[Decoupled.scala 361:21]
  wire  q_210_reset; // @[Decoupled.scala 361:21]
  wire  q_210_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_210_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_210_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_210_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_210_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_210_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_211_clock; // @[Decoupled.scala 361:21]
  wire  q_211_reset; // @[Decoupled.scala 361:21]
  wire  q_211_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_211_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_211_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_211_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_211_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_211_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_212_clock; // @[Decoupled.scala 361:21]
  wire  q_212_reset; // @[Decoupled.scala 361:21]
  wire  q_212_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_212_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_212_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_212_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_212_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_212_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_213_clock; // @[Decoupled.scala 361:21]
  wire  q_213_reset; // @[Decoupled.scala 361:21]
  wire  q_213_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_213_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_213_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_213_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_213_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_213_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_214_clock; // @[Decoupled.scala 361:21]
  wire  q_214_reset; // @[Decoupled.scala 361:21]
  wire  q_214_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_214_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_214_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_214_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_214_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_214_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_215_clock; // @[Decoupled.scala 361:21]
  wire  q_215_reset; // @[Decoupled.scala 361:21]
  wire  q_215_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_215_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_215_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_215_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_215_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_215_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_216_clock; // @[Decoupled.scala 361:21]
  wire  q_216_reset; // @[Decoupled.scala 361:21]
  wire  q_216_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_216_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_216_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_216_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_216_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_216_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_217_clock; // @[Decoupled.scala 361:21]
  wire  q_217_reset; // @[Decoupled.scala 361:21]
  wire  q_217_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_217_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_217_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_217_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_217_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_217_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_218_clock; // @[Decoupled.scala 361:21]
  wire  q_218_reset; // @[Decoupled.scala 361:21]
  wire  q_218_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_218_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_218_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_218_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_218_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_218_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_219_clock; // @[Decoupled.scala 361:21]
  wire  q_219_reset; // @[Decoupled.scala 361:21]
  wire  q_219_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_219_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_219_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_219_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_219_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_219_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_220_clock; // @[Decoupled.scala 361:21]
  wire  q_220_reset; // @[Decoupled.scala 361:21]
  wire  q_220_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_220_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_220_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_220_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_220_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_220_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_221_clock; // @[Decoupled.scala 361:21]
  wire  q_221_reset; // @[Decoupled.scala 361:21]
  wire  q_221_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_221_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_221_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_221_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_221_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_221_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_222_clock; // @[Decoupled.scala 361:21]
  wire  q_222_reset; // @[Decoupled.scala 361:21]
  wire  q_222_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_222_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_222_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_222_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_222_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_222_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_223_clock; // @[Decoupled.scala 361:21]
  wire  q_223_reset; // @[Decoupled.scala 361:21]
  wire  q_223_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_223_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_223_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_223_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_223_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_223_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_224_clock; // @[Decoupled.scala 361:21]
  wire  q_224_reset; // @[Decoupled.scala 361:21]
  wire  q_224_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_224_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_224_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_224_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_224_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_224_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_225_clock; // @[Decoupled.scala 361:21]
  wire  q_225_reset; // @[Decoupled.scala 361:21]
  wire  q_225_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_225_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_225_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_225_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_225_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_225_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_226_clock; // @[Decoupled.scala 361:21]
  wire  q_226_reset; // @[Decoupled.scala 361:21]
  wire  q_226_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_226_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_226_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_226_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_226_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_226_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_227_clock; // @[Decoupled.scala 361:21]
  wire  q_227_reset; // @[Decoupled.scala 361:21]
  wire  q_227_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_227_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_227_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_227_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_227_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_227_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_228_clock; // @[Decoupled.scala 361:21]
  wire  q_228_reset; // @[Decoupled.scala 361:21]
  wire  q_228_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_228_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_228_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_228_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_228_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_228_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_229_clock; // @[Decoupled.scala 361:21]
  wire  q_229_reset; // @[Decoupled.scala 361:21]
  wire  q_229_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_229_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_229_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_229_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_229_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_229_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_230_clock; // @[Decoupled.scala 361:21]
  wire  q_230_reset; // @[Decoupled.scala 361:21]
  wire  q_230_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_230_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_230_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_230_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_230_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_230_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_231_clock; // @[Decoupled.scala 361:21]
  wire  q_231_reset; // @[Decoupled.scala 361:21]
  wire  q_231_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_231_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_231_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_231_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_231_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_231_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_232_clock; // @[Decoupled.scala 361:21]
  wire  q_232_reset; // @[Decoupled.scala 361:21]
  wire  q_232_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_232_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_232_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_232_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_232_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_232_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_233_clock; // @[Decoupled.scala 361:21]
  wire  q_233_reset; // @[Decoupled.scala 361:21]
  wire  q_233_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_233_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_233_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_233_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_233_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_233_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_234_clock; // @[Decoupled.scala 361:21]
  wire  q_234_reset; // @[Decoupled.scala 361:21]
  wire  q_234_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_234_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_234_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_234_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_234_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_234_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_235_clock; // @[Decoupled.scala 361:21]
  wire  q_235_reset; // @[Decoupled.scala 361:21]
  wire  q_235_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_235_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_235_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_235_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_235_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_235_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_236_clock; // @[Decoupled.scala 361:21]
  wire  q_236_reset; // @[Decoupled.scala 361:21]
  wire  q_236_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_236_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_236_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_236_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_236_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_236_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_237_clock; // @[Decoupled.scala 361:21]
  wire  q_237_reset; // @[Decoupled.scala 361:21]
  wire  q_237_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_237_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_237_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_237_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_237_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_237_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_238_clock; // @[Decoupled.scala 361:21]
  wire  q_238_reset; // @[Decoupled.scala 361:21]
  wire  q_238_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_238_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_238_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_238_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_238_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_238_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_239_clock; // @[Decoupled.scala 361:21]
  wire  q_239_reset; // @[Decoupled.scala 361:21]
  wire  q_239_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_239_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_239_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_239_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_239_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_239_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_240_clock; // @[Decoupled.scala 361:21]
  wire  q_240_reset; // @[Decoupled.scala 361:21]
  wire  q_240_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_240_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_240_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_240_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_240_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_240_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_241_clock; // @[Decoupled.scala 361:21]
  wire  q_241_reset; // @[Decoupled.scala 361:21]
  wire  q_241_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_241_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_241_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_241_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_241_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_241_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_242_clock; // @[Decoupled.scala 361:21]
  wire  q_242_reset; // @[Decoupled.scala 361:21]
  wire  q_242_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_242_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_242_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_242_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_242_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_242_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_243_clock; // @[Decoupled.scala 361:21]
  wire  q_243_reset; // @[Decoupled.scala 361:21]
  wire  q_243_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_243_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_243_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_243_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_243_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_243_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_244_clock; // @[Decoupled.scala 361:21]
  wire  q_244_reset; // @[Decoupled.scala 361:21]
  wire  q_244_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_244_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_244_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_244_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_244_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_244_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_245_clock; // @[Decoupled.scala 361:21]
  wire  q_245_reset; // @[Decoupled.scala 361:21]
  wire  q_245_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_245_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_245_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_245_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_245_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_245_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_246_clock; // @[Decoupled.scala 361:21]
  wire  q_246_reset; // @[Decoupled.scala 361:21]
  wire  q_246_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_246_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_246_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_246_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_246_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_246_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_247_clock; // @[Decoupled.scala 361:21]
  wire  q_247_reset; // @[Decoupled.scala 361:21]
  wire  q_247_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_247_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_247_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_247_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_247_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_247_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_248_clock; // @[Decoupled.scala 361:21]
  wire  q_248_reset; // @[Decoupled.scala 361:21]
  wire  q_248_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_248_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_248_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_248_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_248_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_248_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_249_clock; // @[Decoupled.scala 361:21]
  wire  q_249_reset; // @[Decoupled.scala 361:21]
  wire  q_249_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_249_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_249_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_249_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_249_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_249_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_250_clock; // @[Decoupled.scala 361:21]
  wire  q_250_reset; // @[Decoupled.scala 361:21]
  wire  q_250_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_250_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_250_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_250_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_250_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_250_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_251_clock; // @[Decoupled.scala 361:21]
  wire  q_251_reset; // @[Decoupled.scala 361:21]
  wire  q_251_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_251_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_251_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_251_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_251_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_251_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_252_clock; // @[Decoupled.scala 361:21]
  wire  q_252_reset; // @[Decoupled.scala 361:21]
  wire  q_252_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_252_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_252_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_252_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_252_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_252_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_253_clock; // @[Decoupled.scala 361:21]
  wire  q_253_reset; // @[Decoupled.scala 361:21]
  wire  q_253_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_253_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_253_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_253_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_253_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_253_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_254_clock; // @[Decoupled.scala 361:21]
  wire  q_254_reset; // @[Decoupled.scala 361:21]
  wire  q_254_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_254_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_254_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_254_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_254_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_254_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_255_clock; // @[Decoupled.scala 361:21]
  wire  q_255_reset; // @[Decoupled.scala 361:21]
  wire  q_255_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_255_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_255_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_255_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_255_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_255_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_256_clock; // @[Decoupled.scala 361:21]
  wire  q_256_reset; // @[Decoupled.scala 361:21]
  wire  q_256_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_256_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_256_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_256_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_256_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_256_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_257_clock; // @[Decoupled.scala 361:21]
  wire  q_257_reset; // @[Decoupled.scala 361:21]
  wire  q_257_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_257_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_257_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_257_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_257_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_257_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_258_clock; // @[Decoupled.scala 361:21]
  wire  q_258_reset; // @[Decoupled.scala 361:21]
  wire  q_258_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_258_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_258_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_258_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_258_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_258_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_259_clock; // @[Decoupled.scala 361:21]
  wire  q_259_reset; // @[Decoupled.scala 361:21]
  wire  q_259_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_259_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_259_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_259_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_259_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_259_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_260_clock; // @[Decoupled.scala 361:21]
  wire  q_260_reset; // @[Decoupled.scala 361:21]
  wire  q_260_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_260_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_260_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_260_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_260_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_260_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_261_clock; // @[Decoupled.scala 361:21]
  wire  q_261_reset; // @[Decoupled.scala 361:21]
  wire  q_261_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_261_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_261_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_261_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_261_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_261_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_262_clock; // @[Decoupled.scala 361:21]
  wire  q_262_reset; // @[Decoupled.scala 361:21]
  wire  q_262_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_262_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_262_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_262_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_262_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_262_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_263_clock; // @[Decoupled.scala 361:21]
  wire  q_263_reset; // @[Decoupled.scala 361:21]
  wire  q_263_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_263_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_263_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_263_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_263_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_263_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_264_clock; // @[Decoupled.scala 361:21]
  wire  q_264_reset; // @[Decoupled.scala 361:21]
  wire  q_264_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_264_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_264_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_264_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_264_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_264_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_265_clock; // @[Decoupled.scala 361:21]
  wire  q_265_reset; // @[Decoupled.scala 361:21]
  wire  q_265_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_265_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_265_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_265_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_265_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_265_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_266_clock; // @[Decoupled.scala 361:21]
  wire  q_266_reset; // @[Decoupled.scala 361:21]
  wire  q_266_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_266_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_266_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_266_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_266_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_266_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_267_clock; // @[Decoupled.scala 361:21]
  wire  q_267_reset; // @[Decoupled.scala 361:21]
  wire  q_267_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_267_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_267_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_267_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_267_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_267_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_268_clock; // @[Decoupled.scala 361:21]
  wire  q_268_reset; // @[Decoupled.scala 361:21]
  wire  q_268_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_268_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_268_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_268_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_268_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_268_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_269_clock; // @[Decoupled.scala 361:21]
  wire  q_269_reset; // @[Decoupled.scala 361:21]
  wire  q_269_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_269_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_269_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_269_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_269_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_269_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_270_clock; // @[Decoupled.scala 361:21]
  wire  q_270_reset; // @[Decoupled.scala 361:21]
  wire  q_270_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_270_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_270_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_270_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_270_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_270_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_271_clock; // @[Decoupled.scala 361:21]
  wire  q_271_reset; // @[Decoupled.scala 361:21]
  wire  q_271_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_271_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_271_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_271_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_271_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_271_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_272_clock; // @[Decoupled.scala 361:21]
  wire  q_272_reset; // @[Decoupled.scala 361:21]
  wire  q_272_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_272_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_272_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_272_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_272_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_272_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_273_clock; // @[Decoupled.scala 361:21]
  wire  q_273_reset; // @[Decoupled.scala 361:21]
  wire  q_273_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_273_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_273_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_273_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_273_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_273_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_274_clock; // @[Decoupled.scala 361:21]
  wire  q_274_reset; // @[Decoupled.scala 361:21]
  wire  q_274_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_274_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_274_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_274_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_274_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_274_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_275_clock; // @[Decoupled.scala 361:21]
  wire  q_275_reset; // @[Decoupled.scala 361:21]
  wire  q_275_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_275_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_275_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_275_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_275_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_275_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_276_clock; // @[Decoupled.scala 361:21]
  wire  q_276_reset; // @[Decoupled.scala 361:21]
  wire  q_276_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_276_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_276_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_276_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_276_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_276_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_277_clock; // @[Decoupled.scala 361:21]
  wire  q_277_reset; // @[Decoupled.scala 361:21]
  wire  q_277_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_277_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_277_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_277_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_277_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_277_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_278_clock; // @[Decoupled.scala 361:21]
  wire  q_278_reset; // @[Decoupled.scala 361:21]
  wire  q_278_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_278_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_278_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_278_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_278_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_278_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_279_clock; // @[Decoupled.scala 361:21]
  wire  q_279_reset; // @[Decoupled.scala 361:21]
  wire  q_279_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_279_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_279_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_279_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_279_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_279_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_280_clock; // @[Decoupled.scala 361:21]
  wire  q_280_reset; // @[Decoupled.scala 361:21]
  wire  q_280_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_280_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_280_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_280_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_280_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_280_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_281_clock; // @[Decoupled.scala 361:21]
  wire  q_281_reset; // @[Decoupled.scala 361:21]
  wire  q_281_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_281_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_281_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_281_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_281_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_281_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_282_clock; // @[Decoupled.scala 361:21]
  wire  q_282_reset; // @[Decoupled.scala 361:21]
  wire  q_282_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_282_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_282_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_282_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_282_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_282_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_283_clock; // @[Decoupled.scala 361:21]
  wire  q_283_reset; // @[Decoupled.scala 361:21]
  wire  q_283_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_283_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_283_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_283_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_283_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_283_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_284_clock; // @[Decoupled.scala 361:21]
  wire  q_284_reset; // @[Decoupled.scala 361:21]
  wire  q_284_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_284_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_284_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_284_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_284_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_284_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_285_clock; // @[Decoupled.scala 361:21]
  wire  q_285_reset; // @[Decoupled.scala 361:21]
  wire  q_285_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_285_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_285_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_285_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_285_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_285_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_286_clock; // @[Decoupled.scala 361:21]
  wire  q_286_reset; // @[Decoupled.scala 361:21]
  wire  q_286_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_286_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_286_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_286_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_286_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_286_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_287_clock; // @[Decoupled.scala 361:21]
  wire  q_287_reset; // @[Decoupled.scala 361:21]
  wire  q_287_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_287_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_287_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_287_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_287_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_287_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_288_clock; // @[Decoupled.scala 361:21]
  wire  q_288_reset; // @[Decoupled.scala 361:21]
  wire  q_288_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_288_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_288_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_288_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_288_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_288_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_289_clock; // @[Decoupled.scala 361:21]
  wire  q_289_reset; // @[Decoupled.scala 361:21]
  wire  q_289_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_289_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_289_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_289_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_289_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_289_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_290_clock; // @[Decoupled.scala 361:21]
  wire  q_290_reset; // @[Decoupled.scala 361:21]
  wire  q_290_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_290_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_290_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_290_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_290_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_290_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_291_clock; // @[Decoupled.scala 361:21]
  wire  q_291_reset; // @[Decoupled.scala 361:21]
  wire  q_291_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_291_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_291_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_291_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_291_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_291_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_292_clock; // @[Decoupled.scala 361:21]
  wire  q_292_reset; // @[Decoupled.scala 361:21]
  wire  q_292_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_292_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_292_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_292_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_292_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_292_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_293_clock; // @[Decoupled.scala 361:21]
  wire  q_293_reset; // @[Decoupled.scala 361:21]
  wire  q_293_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_293_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_293_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_293_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_293_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_293_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_294_clock; // @[Decoupled.scala 361:21]
  wire  q_294_reset; // @[Decoupled.scala 361:21]
  wire  q_294_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_294_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_294_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_294_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_294_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_294_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_295_clock; // @[Decoupled.scala 361:21]
  wire  q_295_reset; // @[Decoupled.scala 361:21]
  wire  q_295_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_295_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_295_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_295_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_295_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_295_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_296_clock; // @[Decoupled.scala 361:21]
  wire  q_296_reset; // @[Decoupled.scala 361:21]
  wire  q_296_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_296_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_296_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_296_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_296_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_296_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_297_clock; // @[Decoupled.scala 361:21]
  wire  q_297_reset; // @[Decoupled.scala 361:21]
  wire  q_297_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_297_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_297_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_297_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_297_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_297_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_298_clock; // @[Decoupled.scala 361:21]
  wire  q_298_reset; // @[Decoupled.scala 361:21]
  wire  q_298_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_298_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_298_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_298_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_298_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_298_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_299_clock; // @[Decoupled.scala 361:21]
  wire  q_299_reset; // @[Decoupled.scala 361:21]
  wire  q_299_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_299_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_299_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_299_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_299_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_299_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_300_clock; // @[Decoupled.scala 361:21]
  wire  q_300_reset; // @[Decoupled.scala 361:21]
  wire  q_300_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_300_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_300_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_300_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_300_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_300_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_301_clock; // @[Decoupled.scala 361:21]
  wire  q_301_reset; // @[Decoupled.scala 361:21]
  wire  q_301_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_301_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_301_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_301_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_301_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_301_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_302_clock; // @[Decoupled.scala 361:21]
  wire  q_302_reset; // @[Decoupled.scala 361:21]
  wire  q_302_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_302_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_302_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_302_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_302_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_302_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_303_clock; // @[Decoupled.scala 361:21]
  wire  q_303_reset; // @[Decoupled.scala 361:21]
  wire  q_303_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_303_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_303_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_303_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_303_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_303_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_304_clock; // @[Decoupled.scala 361:21]
  wire  q_304_reset; // @[Decoupled.scala 361:21]
  wire  q_304_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_304_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_304_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_304_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_304_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_304_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_305_clock; // @[Decoupled.scala 361:21]
  wire  q_305_reset; // @[Decoupled.scala 361:21]
  wire  q_305_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_305_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_305_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_305_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_305_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_305_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_306_clock; // @[Decoupled.scala 361:21]
  wire  q_306_reset; // @[Decoupled.scala 361:21]
  wire  q_306_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_306_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_306_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_306_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_306_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_306_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_307_clock; // @[Decoupled.scala 361:21]
  wire  q_307_reset; // @[Decoupled.scala 361:21]
  wire  q_307_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_307_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_307_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_307_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_307_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_307_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_308_clock; // @[Decoupled.scala 361:21]
  wire  q_308_reset; // @[Decoupled.scala 361:21]
  wire  q_308_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_308_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_308_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_308_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_308_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_308_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_309_clock; // @[Decoupled.scala 361:21]
  wire  q_309_reset; // @[Decoupled.scala 361:21]
  wire  q_309_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_309_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_309_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_309_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_309_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_309_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_310_clock; // @[Decoupled.scala 361:21]
  wire  q_310_reset; // @[Decoupled.scala 361:21]
  wire  q_310_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_310_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_310_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_310_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_310_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_310_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_311_clock; // @[Decoupled.scala 361:21]
  wire  q_311_reset; // @[Decoupled.scala 361:21]
  wire  q_311_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_311_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_311_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_311_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_311_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_311_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_312_clock; // @[Decoupled.scala 361:21]
  wire  q_312_reset; // @[Decoupled.scala 361:21]
  wire  q_312_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_312_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_312_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_312_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_312_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_312_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_313_clock; // @[Decoupled.scala 361:21]
  wire  q_313_reset; // @[Decoupled.scala 361:21]
  wire  q_313_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_313_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_313_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_313_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_313_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_313_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_314_clock; // @[Decoupled.scala 361:21]
  wire  q_314_reset; // @[Decoupled.scala 361:21]
  wire  q_314_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_314_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_314_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_314_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_314_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_314_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_315_clock; // @[Decoupled.scala 361:21]
  wire  q_315_reset; // @[Decoupled.scala 361:21]
  wire  q_315_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_315_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_315_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_315_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_315_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_315_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_316_clock; // @[Decoupled.scala 361:21]
  wire  q_316_reset; // @[Decoupled.scala 361:21]
  wire  q_316_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_316_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_316_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_316_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_316_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_316_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_317_clock; // @[Decoupled.scala 361:21]
  wire  q_317_reset; // @[Decoupled.scala 361:21]
  wire  q_317_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_317_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_317_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_317_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_317_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_317_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_318_clock; // @[Decoupled.scala 361:21]
  wire  q_318_reset; // @[Decoupled.scala 361:21]
  wire  q_318_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_318_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_318_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_318_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_318_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_318_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_319_clock; // @[Decoupled.scala 361:21]
  wire  q_319_reset; // @[Decoupled.scala 361:21]
  wire  q_319_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_319_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_319_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_319_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_319_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_319_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_320_clock; // @[Decoupled.scala 361:21]
  wire  q_320_reset; // @[Decoupled.scala 361:21]
  wire  q_320_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_320_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_320_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_320_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_320_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_320_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_321_clock; // @[Decoupled.scala 361:21]
  wire  q_321_reset; // @[Decoupled.scala 361:21]
  wire  q_321_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_321_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_321_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_321_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_321_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_321_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_322_clock; // @[Decoupled.scala 361:21]
  wire  q_322_reset; // @[Decoupled.scala 361:21]
  wire  q_322_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_322_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_322_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_322_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_322_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_322_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_323_clock; // @[Decoupled.scala 361:21]
  wire  q_323_reset; // @[Decoupled.scala 361:21]
  wire  q_323_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_323_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_323_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_323_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_323_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_323_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_324_clock; // @[Decoupled.scala 361:21]
  wire  q_324_reset; // @[Decoupled.scala 361:21]
  wire  q_324_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_324_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_324_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_324_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_324_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_324_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_325_clock; // @[Decoupled.scala 361:21]
  wire  q_325_reset; // @[Decoupled.scala 361:21]
  wire  q_325_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_325_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_325_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_325_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_325_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_325_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_326_clock; // @[Decoupled.scala 361:21]
  wire  q_326_reset; // @[Decoupled.scala 361:21]
  wire  q_326_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_326_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_326_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_326_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_326_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_326_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_327_clock; // @[Decoupled.scala 361:21]
  wire  q_327_reset; // @[Decoupled.scala 361:21]
  wire  q_327_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_327_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_327_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_327_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_327_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_327_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_328_clock; // @[Decoupled.scala 361:21]
  wire  q_328_reset; // @[Decoupled.scala 361:21]
  wire  q_328_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_328_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_328_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_328_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_328_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_328_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_329_clock; // @[Decoupled.scala 361:21]
  wire  q_329_reset; // @[Decoupled.scala 361:21]
  wire  q_329_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_329_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_329_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_329_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_329_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_329_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_330_clock; // @[Decoupled.scala 361:21]
  wire  q_330_reset; // @[Decoupled.scala 361:21]
  wire  q_330_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_330_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_330_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_330_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_330_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_330_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_331_clock; // @[Decoupled.scala 361:21]
  wire  q_331_reset; // @[Decoupled.scala 361:21]
  wire  q_331_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_331_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_331_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_331_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_331_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_331_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_332_clock; // @[Decoupled.scala 361:21]
  wire  q_332_reset; // @[Decoupled.scala 361:21]
  wire  q_332_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_332_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_332_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_332_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_332_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_332_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_333_clock; // @[Decoupled.scala 361:21]
  wire  q_333_reset; // @[Decoupled.scala 361:21]
  wire  q_333_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_333_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_333_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_333_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_333_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_333_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_334_clock; // @[Decoupled.scala 361:21]
  wire  q_334_reset; // @[Decoupled.scala 361:21]
  wire  q_334_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_334_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_334_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_334_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_334_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_334_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_335_clock; // @[Decoupled.scala 361:21]
  wire  q_335_reset; // @[Decoupled.scala 361:21]
  wire  q_335_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_335_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_335_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_335_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_335_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_335_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_336_clock; // @[Decoupled.scala 361:21]
  wire  q_336_reset; // @[Decoupled.scala 361:21]
  wire  q_336_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_336_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_336_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_336_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_336_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_336_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_337_clock; // @[Decoupled.scala 361:21]
  wire  q_337_reset; // @[Decoupled.scala 361:21]
  wire  q_337_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_337_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_337_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_337_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_337_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_337_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_338_clock; // @[Decoupled.scala 361:21]
  wire  q_338_reset; // @[Decoupled.scala 361:21]
  wire  q_338_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_338_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_338_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_338_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_338_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_338_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_339_clock; // @[Decoupled.scala 361:21]
  wire  q_339_reset; // @[Decoupled.scala 361:21]
  wire  q_339_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_339_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_339_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_339_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_339_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_339_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_340_clock; // @[Decoupled.scala 361:21]
  wire  q_340_reset; // @[Decoupled.scala 361:21]
  wire  q_340_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_340_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_340_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_340_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_340_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_340_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_341_clock; // @[Decoupled.scala 361:21]
  wire  q_341_reset; // @[Decoupled.scala 361:21]
  wire  q_341_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_341_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_341_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_341_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_341_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_341_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_342_clock; // @[Decoupled.scala 361:21]
  wire  q_342_reset; // @[Decoupled.scala 361:21]
  wire  q_342_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_342_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_342_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_342_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_342_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_342_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_343_clock; // @[Decoupled.scala 361:21]
  wire  q_343_reset; // @[Decoupled.scala 361:21]
  wire  q_343_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_343_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_343_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_343_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_343_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_343_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_344_clock; // @[Decoupled.scala 361:21]
  wire  q_344_reset; // @[Decoupled.scala 361:21]
  wire  q_344_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_344_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_344_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_344_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_344_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_344_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_345_clock; // @[Decoupled.scala 361:21]
  wire  q_345_reset; // @[Decoupled.scala 361:21]
  wire  q_345_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_345_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_345_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_345_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_345_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_345_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_346_clock; // @[Decoupled.scala 361:21]
  wire  q_346_reset; // @[Decoupled.scala 361:21]
  wire  q_346_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_346_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_346_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_346_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_346_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_346_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_347_clock; // @[Decoupled.scala 361:21]
  wire  q_347_reset; // @[Decoupled.scala 361:21]
  wire  q_347_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_347_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_347_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_347_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_347_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_347_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_348_clock; // @[Decoupled.scala 361:21]
  wire  q_348_reset; // @[Decoupled.scala 361:21]
  wire  q_348_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_348_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_348_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_348_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_348_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_348_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_349_clock; // @[Decoupled.scala 361:21]
  wire  q_349_reset; // @[Decoupled.scala 361:21]
  wire  q_349_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_349_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_349_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_349_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_349_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_349_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_350_clock; // @[Decoupled.scala 361:21]
  wire  q_350_reset; // @[Decoupled.scala 361:21]
  wire  q_350_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_350_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_350_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_350_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_350_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_350_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_351_clock; // @[Decoupled.scala 361:21]
  wire  q_351_reset; // @[Decoupled.scala 361:21]
  wire  q_351_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_351_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_351_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_351_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_351_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_351_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_352_clock; // @[Decoupled.scala 361:21]
  wire  q_352_reset; // @[Decoupled.scala 361:21]
  wire  q_352_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_352_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_352_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_352_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_352_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_352_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_353_clock; // @[Decoupled.scala 361:21]
  wire  q_353_reset; // @[Decoupled.scala 361:21]
  wire  q_353_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_353_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_353_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_353_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_353_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_353_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_354_clock; // @[Decoupled.scala 361:21]
  wire  q_354_reset; // @[Decoupled.scala 361:21]
  wire  q_354_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_354_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_354_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_354_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_354_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_354_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_355_clock; // @[Decoupled.scala 361:21]
  wire  q_355_reset; // @[Decoupled.scala 361:21]
  wire  q_355_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_355_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_355_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_355_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_355_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_355_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_356_clock; // @[Decoupled.scala 361:21]
  wire  q_356_reset; // @[Decoupled.scala 361:21]
  wire  q_356_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_356_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_356_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_356_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_356_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_356_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_357_clock; // @[Decoupled.scala 361:21]
  wire  q_357_reset; // @[Decoupled.scala 361:21]
  wire  q_357_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_357_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_357_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_357_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_357_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_357_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_358_clock; // @[Decoupled.scala 361:21]
  wire  q_358_reset; // @[Decoupled.scala 361:21]
  wire  q_358_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_358_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_358_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_358_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_358_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_358_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_359_clock; // @[Decoupled.scala 361:21]
  wire  q_359_reset; // @[Decoupled.scala 361:21]
  wire  q_359_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_359_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_359_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_359_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_359_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_359_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_360_clock; // @[Decoupled.scala 361:21]
  wire  q_360_reset; // @[Decoupled.scala 361:21]
  wire  q_360_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_360_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_360_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_360_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_360_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_360_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_361_clock; // @[Decoupled.scala 361:21]
  wire  q_361_reset; // @[Decoupled.scala 361:21]
  wire  q_361_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_361_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_361_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_361_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_361_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_361_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_362_clock; // @[Decoupled.scala 361:21]
  wire  q_362_reset; // @[Decoupled.scala 361:21]
  wire  q_362_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_362_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_362_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_362_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_362_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_362_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_363_clock; // @[Decoupled.scala 361:21]
  wire  q_363_reset; // @[Decoupled.scala 361:21]
  wire  q_363_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_363_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_363_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_363_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_363_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_363_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_364_clock; // @[Decoupled.scala 361:21]
  wire  q_364_reset; // @[Decoupled.scala 361:21]
  wire  q_364_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_364_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_364_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_364_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_364_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_364_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_365_clock; // @[Decoupled.scala 361:21]
  wire  q_365_reset; // @[Decoupled.scala 361:21]
  wire  q_365_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_365_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_365_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_365_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_365_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_365_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_366_clock; // @[Decoupled.scala 361:21]
  wire  q_366_reset; // @[Decoupled.scala 361:21]
  wire  q_366_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_366_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_366_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_366_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_366_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_366_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_367_clock; // @[Decoupled.scala 361:21]
  wire  q_367_reset; // @[Decoupled.scala 361:21]
  wire  q_367_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_367_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_367_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_367_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_367_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_367_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_368_clock; // @[Decoupled.scala 361:21]
  wire  q_368_reset; // @[Decoupled.scala 361:21]
  wire  q_368_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_368_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_368_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_368_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_368_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_368_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_369_clock; // @[Decoupled.scala 361:21]
  wire  q_369_reset; // @[Decoupled.scala 361:21]
  wire  q_369_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_369_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_369_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_369_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_369_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_369_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_370_clock; // @[Decoupled.scala 361:21]
  wire  q_370_reset; // @[Decoupled.scala 361:21]
  wire  q_370_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_370_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_370_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_370_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_370_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_370_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_371_clock; // @[Decoupled.scala 361:21]
  wire  q_371_reset; // @[Decoupled.scala 361:21]
  wire  q_371_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_371_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_371_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_371_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_371_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_371_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_372_clock; // @[Decoupled.scala 361:21]
  wire  q_372_reset; // @[Decoupled.scala 361:21]
  wire  q_372_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_372_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_372_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_372_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_372_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_372_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_373_clock; // @[Decoupled.scala 361:21]
  wire  q_373_reset; // @[Decoupled.scala 361:21]
  wire  q_373_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_373_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_373_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_373_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_373_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_373_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_374_clock; // @[Decoupled.scala 361:21]
  wire  q_374_reset; // @[Decoupled.scala 361:21]
  wire  q_374_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_374_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_374_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_374_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_374_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_374_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_375_clock; // @[Decoupled.scala 361:21]
  wire  q_375_reset; // @[Decoupled.scala 361:21]
  wire  q_375_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_375_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_375_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_375_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_375_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_375_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_376_clock; // @[Decoupled.scala 361:21]
  wire  q_376_reset; // @[Decoupled.scala 361:21]
  wire  q_376_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_376_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_376_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_376_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_376_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_376_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_377_clock; // @[Decoupled.scala 361:21]
  wire  q_377_reset; // @[Decoupled.scala 361:21]
  wire  q_377_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_377_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_377_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_377_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_377_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_377_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_378_clock; // @[Decoupled.scala 361:21]
  wire  q_378_reset; // @[Decoupled.scala 361:21]
  wire  q_378_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_378_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_378_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_378_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_378_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_378_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_379_clock; // @[Decoupled.scala 361:21]
  wire  q_379_reset; // @[Decoupled.scala 361:21]
  wire  q_379_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_379_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_379_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_379_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_379_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_379_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_380_clock; // @[Decoupled.scala 361:21]
  wire  q_380_reset; // @[Decoupled.scala 361:21]
  wire  q_380_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_380_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_380_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_380_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_380_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_380_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_381_clock; // @[Decoupled.scala 361:21]
  wire  q_381_reset; // @[Decoupled.scala 361:21]
  wire  q_381_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_381_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_381_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_381_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_381_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_381_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_382_clock; // @[Decoupled.scala 361:21]
  wire  q_382_reset; // @[Decoupled.scala 361:21]
  wire  q_382_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_382_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_382_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_382_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_382_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_382_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_383_clock; // @[Decoupled.scala 361:21]
  wire  q_383_reset; // @[Decoupled.scala 361:21]
  wire  q_383_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_383_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_383_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_383_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_383_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_383_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_384_clock; // @[Decoupled.scala 361:21]
  wire  q_384_reset; // @[Decoupled.scala 361:21]
  wire  q_384_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_384_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_384_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_384_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_384_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_384_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_385_clock; // @[Decoupled.scala 361:21]
  wire  q_385_reset; // @[Decoupled.scala 361:21]
  wire  q_385_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_385_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_385_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_385_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_385_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_385_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_386_clock; // @[Decoupled.scala 361:21]
  wire  q_386_reset; // @[Decoupled.scala 361:21]
  wire  q_386_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_386_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_386_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_386_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_386_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_386_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_387_clock; // @[Decoupled.scala 361:21]
  wire  q_387_reset; // @[Decoupled.scala 361:21]
  wire  q_387_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_387_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_387_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_387_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_387_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_387_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_388_clock; // @[Decoupled.scala 361:21]
  wire  q_388_reset; // @[Decoupled.scala 361:21]
  wire  q_388_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_388_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_388_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_388_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_388_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_388_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_389_clock; // @[Decoupled.scala 361:21]
  wire  q_389_reset; // @[Decoupled.scala 361:21]
  wire  q_389_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_389_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_389_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_389_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_389_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_389_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_390_clock; // @[Decoupled.scala 361:21]
  wire  q_390_reset; // @[Decoupled.scala 361:21]
  wire  q_390_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_390_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_390_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_390_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_390_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_390_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_391_clock; // @[Decoupled.scala 361:21]
  wire  q_391_reset; // @[Decoupled.scala 361:21]
  wire  q_391_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_391_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_391_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_391_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_391_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_391_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_392_clock; // @[Decoupled.scala 361:21]
  wire  q_392_reset; // @[Decoupled.scala 361:21]
  wire  q_392_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_392_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_392_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_392_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_392_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_392_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_393_clock; // @[Decoupled.scala 361:21]
  wire  q_393_reset; // @[Decoupled.scala 361:21]
  wire  q_393_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_393_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_393_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_393_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_393_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_393_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_394_clock; // @[Decoupled.scala 361:21]
  wire  q_394_reset; // @[Decoupled.scala 361:21]
  wire  q_394_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_394_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_394_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_394_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_394_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_394_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_395_clock; // @[Decoupled.scala 361:21]
  wire  q_395_reset; // @[Decoupled.scala 361:21]
  wire  q_395_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_395_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_395_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_395_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_395_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_395_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_396_clock; // @[Decoupled.scala 361:21]
  wire  q_396_reset; // @[Decoupled.scala 361:21]
  wire  q_396_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_396_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_396_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_396_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_396_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_396_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_397_clock; // @[Decoupled.scala 361:21]
  wire  q_397_reset; // @[Decoupled.scala 361:21]
  wire  q_397_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_397_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_397_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_397_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_397_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_397_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_398_clock; // @[Decoupled.scala 361:21]
  wire  q_398_reset; // @[Decoupled.scala 361:21]
  wire  q_398_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_398_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_398_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_398_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_398_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_398_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_399_clock; // @[Decoupled.scala 361:21]
  wire  q_399_reset; // @[Decoupled.scala 361:21]
  wire  q_399_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_399_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_399_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_399_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_399_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_399_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_400_clock; // @[Decoupled.scala 361:21]
  wire  q_400_reset; // @[Decoupled.scala 361:21]
  wire  q_400_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_400_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_400_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_400_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_400_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_400_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_401_clock; // @[Decoupled.scala 361:21]
  wire  q_401_reset; // @[Decoupled.scala 361:21]
  wire  q_401_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_401_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_401_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_401_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_401_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_401_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_402_clock; // @[Decoupled.scala 361:21]
  wire  q_402_reset; // @[Decoupled.scala 361:21]
  wire  q_402_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_402_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_402_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_402_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_402_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_402_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_403_clock; // @[Decoupled.scala 361:21]
  wire  q_403_reset; // @[Decoupled.scala 361:21]
  wire  q_403_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_403_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_403_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_403_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_403_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_403_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_404_clock; // @[Decoupled.scala 361:21]
  wire  q_404_reset; // @[Decoupled.scala 361:21]
  wire  q_404_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_404_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_404_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_404_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_404_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_404_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_405_clock; // @[Decoupled.scala 361:21]
  wire  q_405_reset; // @[Decoupled.scala 361:21]
  wire  q_405_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_405_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_405_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_405_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_405_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_405_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_406_clock; // @[Decoupled.scala 361:21]
  wire  q_406_reset; // @[Decoupled.scala 361:21]
  wire  q_406_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_406_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_406_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_406_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_406_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_406_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_407_clock; // @[Decoupled.scala 361:21]
  wire  q_407_reset; // @[Decoupled.scala 361:21]
  wire  q_407_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_407_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_407_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_407_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_407_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_407_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_408_clock; // @[Decoupled.scala 361:21]
  wire  q_408_reset; // @[Decoupled.scala 361:21]
  wire  q_408_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_408_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_408_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_408_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_408_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_408_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_409_clock; // @[Decoupled.scala 361:21]
  wire  q_409_reset; // @[Decoupled.scala 361:21]
  wire  q_409_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_409_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_409_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_409_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_409_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_409_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_410_clock; // @[Decoupled.scala 361:21]
  wire  q_410_reset; // @[Decoupled.scala 361:21]
  wire  q_410_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_410_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_410_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_410_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_410_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_410_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_411_clock; // @[Decoupled.scala 361:21]
  wire  q_411_reset; // @[Decoupled.scala 361:21]
  wire  q_411_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_411_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_411_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_411_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_411_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_411_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_412_clock; // @[Decoupled.scala 361:21]
  wire  q_412_reset; // @[Decoupled.scala 361:21]
  wire  q_412_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_412_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_412_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_412_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_412_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_412_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_413_clock; // @[Decoupled.scala 361:21]
  wire  q_413_reset; // @[Decoupled.scala 361:21]
  wire  q_413_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_413_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_413_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_413_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_413_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_413_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_414_clock; // @[Decoupled.scala 361:21]
  wire  q_414_reset; // @[Decoupled.scala 361:21]
  wire  q_414_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_414_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_414_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_414_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_414_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_414_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_415_clock; // @[Decoupled.scala 361:21]
  wire  q_415_reset; // @[Decoupled.scala 361:21]
  wire  q_415_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_415_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_415_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_415_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_415_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_415_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_416_clock; // @[Decoupled.scala 361:21]
  wire  q_416_reset; // @[Decoupled.scala 361:21]
  wire  q_416_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_416_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_416_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_416_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_416_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_416_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_417_clock; // @[Decoupled.scala 361:21]
  wire  q_417_reset; // @[Decoupled.scala 361:21]
  wire  q_417_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_417_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_417_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_417_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_417_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_417_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_418_clock; // @[Decoupled.scala 361:21]
  wire  q_418_reset; // @[Decoupled.scala 361:21]
  wire  q_418_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_418_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_418_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_418_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_418_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_418_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_419_clock; // @[Decoupled.scala 361:21]
  wire  q_419_reset; // @[Decoupled.scala 361:21]
  wire  q_419_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_419_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_419_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_419_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_419_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_419_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_420_clock; // @[Decoupled.scala 361:21]
  wire  q_420_reset; // @[Decoupled.scala 361:21]
  wire  q_420_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_420_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_420_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_420_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_420_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_420_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_421_clock; // @[Decoupled.scala 361:21]
  wire  q_421_reset; // @[Decoupled.scala 361:21]
  wire  q_421_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_421_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_421_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_421_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_421_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_421_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_422_clock; // @[Decoupled.scala 361:21]
  wire  q_422_reset; // @[Decoupled.scala 361:21]
  wire  q_422_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_422_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_422_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_422_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_422_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_422_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_423_clock; // @[Decoupled.scala 361:21]
  wire  q_423_reset; // @[Decoupled.scala 361:21]
  wire  q_423_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_423_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_423_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_423_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_423_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_423_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_424_clock; // @[Decoupled.scala 361:21]
  wire  q_424_reset; // @[Decoupled.scala 361:21]
  wire  q_424_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_424_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_424_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_424_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_424_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_424_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_425_clock; // @[Decoupled.scala 361:21]
  wire  q_425_reset; // @[Decoupled.scala 361:21]
  wire  q_425_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_425_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_425_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_425_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_425_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_425_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_426_clock; // @[Decoupled.scala 361:21]
  wire  q_426_reset; // @[Decoupled.scala 361:21]
  wire  q_426_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_426_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_426_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_426_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_426_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_426_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_427_clock; // @[Decoupled.scala 361:21]
  wire  q_427_reset; // @[Decoupled.scala 361:21]
  wire  q_427_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_427_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_427_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_427_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_427_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_427_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_428_clock; // @[Decoupled.scala 361:21]
  wire  q_428_reset; // @[Decoupled.scala 361:21]
  wire  q_428_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_428_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_428_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_428_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_428_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_428_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_429_clock; // @[Decoupled.scala 361:21]
  wire  q_429_reset; // @[Decoupled.scala 361:21]
  wire  q_429_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_429_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_429_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_429_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_429_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_429_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_430_clock; // @[Decoupled.scala 361:21]
  wire  q_430_reset; // @[Decoupled.scala 361:21]
  wire  q_430_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_430_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_430_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_430_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_430_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_430_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_431_clock; // @[Decoupled.scala 361:21]
  wire  q_431_reset; // @[Decoupled.scala 361:21]
  wire  q_431_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_431_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_431_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_431_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_431_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_431_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_432_clock; // @[Decoupled.scala 361:21]
  wire  q_432_reset; // @[Decoupled.scala 361:21]
  wire  q_432_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_432_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_432_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_432_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_432_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_432_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_433_clock; // @[Decoupled.scala 361:21]
  wire  q_433_reset; // @[Decoupled.scala 361:21]
  wire  q_433_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_433_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_433_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_433_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_433_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_433_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_434_clock; // @[Decoupled.scala 361:21]
  wire  q_434_reset; // @[Decoupled.scala 361:21]
  wire  q_434_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_434_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_434_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_434_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_434_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_434_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_435_clock; // @[Decoupled.scala 361:21]
  wire  q_435_reset; // @[Decoupled.scala 361:21]
  wire  q_435_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_435_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_435_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_435_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_435_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_435_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_436_clock; // @[Decoupled.scala 361:21]
  wire  q_436_reset; // @[Decoupled.scala 361:21]
  wire  q_436_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_436_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_436_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_436_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_436_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_436_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_437_clock; // @[Decoupled.scala 361:21]
  wire  q_437_reset; // @[Decoupled.scala 361:21]
  wire  q_437_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_437_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_437_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_437_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_437_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_437_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_438_clock; // @[Decoupled.scala 361:21]
  wire  q_438_reset; // @[Decoupled.scala 361:21]
  wire  q_438_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_438_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_438_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_438_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_438_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_438_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_439_clock; // @[Decoupled.scala 361:21]
  wire  q_439_reset; // @[Decoupled.scala 361:21]
  wire  q_439_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_439_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_439_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_439_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_439_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_439_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_440_clock; // @[Decoupled.scala 361:21]
  wire  q_440_reset; // @[Decoupled.scala 361:21]
  wire  q_440_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_440_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_440_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_440_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_440_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_440_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_441_clock; // @[Decoupled.scala 361:21]
  wire  q_441_reset; // @[Decoupled.scala 361:21]
  wire  q_441_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_441_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_441_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_441_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_441_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_441_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_442_clock; // @[Decoupled.scala 361:21]
  wire  q_442_reset; // @[Decoupled.scala 361:21]
  wire  q_442_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_442_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_442_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_442_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_442_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_442_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_443_clock; // @[Decoupled.scala 361:21]
  wire  q_443_reset; // @[Decoupled.scala 361:21]
  wire  q_443_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_443_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_443_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_443_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_443_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_443_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_444_clock; // @[Decoupled.scala 361:21]
  wire  q_444_reset; // @[Decoupled.scala 361:21]
  wire  q_444_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_444_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_444_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_444_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_444_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_444_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_445_clock; // @[Decoupled.scala 361:21]
  wire  q_445_reset; // @[Decoupled.scala 361:21]
  wire  q_445_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_445_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_445_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_445_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_445_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_445_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_446_clock; // @[Decoupled.scala 361:21]
  wire  q_446_reset; // @[Decoupled.scala 361:21]
  wire  q_446_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_446_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_446_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_446_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_446_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_446_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_447_clock; // @[Decoupled.scala 361:21]
  wire  q_447_reset; // @[Decoupled.scala 361:21]
  wire  q_447_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_447_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_447_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_447_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_447_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_447_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_448_clock; // @[Decoupled.scala 361:21]
  wire  q_448_reset; // @[Decoupled.scala 361:21]
  wire  q_448_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_448_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_448_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_448_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_448_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_448_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_449_clock; // @[Decoupled.scala 361:21]
  wire  q_449_reset; // @[Decoupled.scala 361:21]
  wire  q_449_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_449_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_449_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_449_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_449_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_449_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_450_clock; // @[Decoupled.scala 361:21]
  wire  q_450_reset; // @[Decoupled.scala 361:21]
  wire  q_450_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_450_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_450_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_450_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_450_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_450_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_451_clock; // @[Decoupled.scala 361:21]
  wire  q_451_reset; // @[Decoupled.scala 361:21]
  wire  q_451_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_451_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_451_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_451_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_451_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_451_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_452_clock; // @[Decoupled.scala 361:21]
  wire  q_452_reset; // @[Decoupled.scala 361:21]
  wire  q_452_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_452_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_452_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_452_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_452_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_452_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_453_clock; // @[Decoupled.scala 361:21]
  wire  q_453_reset; // @[Decoupled.scala 361:21]
  wire  q_453_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_453_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_453_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_453_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_453_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_453_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_454_clock; // @[Decoupled.scala 361:21]
  wire  q_454_reset; // @[Decoupled.scala 361:21]
  wire  q_454_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_454_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_454_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_454_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_454_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_454_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_455_clock; // @[Decoupled.scala 361:21]
  wire  q_455_reset; // @[Decoupled.scala 361:21]
  wire  q_455_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_455_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_455_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_455_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_455_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_455_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_456_clock; // @[Decoupled.scala 361:21]
  wire  q_456_reset; // @[Decoupled.scala 361:21]
  wire  q_456_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_456_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_456_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_456_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_456_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_456_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_457_clock; // @[Decoupled.scala 361:21]
  wire  q_457_reset; // @[Decoupled.scala 361:21]
  wire  q_457_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_457_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_457_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_457_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_457_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_457_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_458_clock; // @[Decoupled.scala 361:21]
  wire  q_458_reset; // @[Decoupled.scala 361:21]
  wire  q_458_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_458_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_458_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_458_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_458_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_458_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_459_clock; // @[Decoupled.scala 361:21]
  wire  q_459_reset; // @[Decoupled.scala 361:21]
  wire  q_459_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_459_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_459_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_459_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_459_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_459_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_460_clock; // @[Decoupled.scala 361:21]
  wire  q_460_reset; // @[Decoupled.scala 361:21]
  wire  q_460_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_460_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_460_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_460_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_460_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_460_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_461_clock; // @[Decoupled.scala 361:21]
  wire  q_461_reset; // @[Decoupled.scala 361:21]
  wire  q_461_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_461_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_461_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_461_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_461_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_461_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_462_clock; // @[Decoupled.scala 361:21]
  wire  q_462_reset; // @[Decoupled.scala 361:21]
  wire  q_462_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_462_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_462_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_462_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_462_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_462_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_463_clock; // @[Decoupled.scala 361:21]
  wire  q_463_reset; // @[Decoupled.scala 361:21]
  wire  q_463_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_463_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_463_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_463_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_463_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_463_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_464_clock; // @[Decoupled.scala 361:21]
  wire  q_464_reset; // @[Decoupled.scala 361:21]
  wire  q_464_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_464_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_464_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_464_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_464_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_464_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_465_clock; // @[Decoupled.scala 361:21]
  wire  q_465_reset; // @[Decoupled.scala 361:21]
  wire  q_465_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_465_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_465_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_465_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_465_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_465_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_466_clock; // @[Decoupled.scala 361:21]
  wire  q_466_reset; // @[Decoupled.scala 361:21]
  wire  q_466_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_466_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_466_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_466_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_466_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_466_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_467_clock; // @[Decoupled.scala 361:21]
  wire  q_467_reset; // @[Decoupled.scala 361:21]
  wire  q_467_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_467_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_467_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_467_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_467_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_467_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_468_clock; // @[Decoupled.scala 361:21]
  wire  q_468_reset; // @[Decoupled.scala 361:21]
  wire  q_468_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_468_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_468_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_468_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_468_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_468_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_469_clock; // @[Decoupled.scala 361:21]
  wire  q_469_reset; // @[Decoupled.scala 361:21]
  wire  q_469_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_469_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_469_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_469_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_469_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_469_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_470_clock; // @[Decoupled.scala 361:21]
  wire  q_470_reset; // @[Decoupled.scala 361:21]
  wire  q_470_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_470_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_470_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_470_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_470_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_470_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_471_clock; // @[Decoupled.scala 361:21]
  wire  q_471_reset; // @[Decoupled.scala 361:21]
  wire  q_471_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_471_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_471_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_471_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_471_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_471_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_472_clock; // @[Decoupled.scala 361:21]
  wire  q_472_reset; // @[Decoupled.scala 361:21]
  wire  q_472_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_472_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_472_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_472_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_472_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_472_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_473_clock; // @[Decoupled.scala 361:21]
  wire  q_473_reset; // @[Decoupled.scala 361:21]
  wire  q_473_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_473_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_473_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_473_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_473_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_473_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_474_clock; // @[Decoupled.scala 361:21]
  wire  q_474_reset; // @[Decoupled.scala 361:21]
  wire  q_474_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_474_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_474_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_474_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_474_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_474_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_475_clock; // @[Decoupled.scala 361:21]
  wire  q_475_reset; // @[Decoupled.scala 361:21]
  wire  q_475_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_475_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_475_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_475_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_475_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_475_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_476_clock; // @[Decoupled.scala 361:21]
  wire  q_476_reset; // @[Decoupled.scala 361:21]
  wire  q_476_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_476_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_476_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_476_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_476_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_476_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_477_clock; // @[Decoupled.scala 361:21]
  wire  q_477_reset; // @[Decoupled.scala 361:21]
  wire  q_477_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_477_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_477_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_477_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_477_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_477_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_478_clock; // @[Decoupled.scala 361:21]
  wire  q_478_reset; // @[Decoupled.scala 361:21]
  wire  q_478_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_478_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_478_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_478_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_478_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_478_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_479_clock; // @[Decoupled.scala 361:21]
  wire  q_479_reset; // @[Decoupled.scala 361:21]
  wire  q_479_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_479_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_479_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_479_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_479_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_479_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_480_clock; // @[Decoupled.scala 361:21]
  wire  q_480_reset; // @[Decoupled.scala 361:21]
  wire  q_480_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_480_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_480_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_480_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_480_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_480_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_481_clock; // @[Decoupled.scala 361:21]
  wire  q_481_reset; // @[Decoupled.scala 361:21]
  wire  q_481_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_481_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_481_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_481_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_481_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_481_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_482_clock; // @[Decoupled.scala 361:21]
  wire  q_482_reset; // @[Decoupled.scala 361:21]
  wire  q_482_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_482_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_482_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_482_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_482_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_482_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_483_clock; // @[Decoupled.scala 361:21]
  wire  q_483_reset; // @[Decoupled.scala 361:21]
  wire  q_483_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_483_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_483_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_483_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_483_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_483_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_484_clock; // @[Decoupled.scala 361:21]
  wire  q_484_reset; // @[Decoupled.scala 361:21]
  wire  q_484_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_484_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_484_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_484_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_484_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_484_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_485_clock; // @[Decoupled.scala 361:21]
  wire  q_485_reset; // @[Decoupled.scala 361:21]
  wire  q_485_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_485_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_485_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_485_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_485_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_485_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_486_clock; // @[Decoupled.scala 361:21]
  wire  q_486_reset; // @[Decoupled.scala 361:21]
  wire  q_486_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_486_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_486_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_486_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_486_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_486_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_487_clock; // @[Decoupled.scala 361:21]
  wire  q_487_reset; // @[Decoupled.scala 361:21]
  wire  q_487_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_487_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_487_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_487_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_487_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_487_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_488_clock; // @[Decoupled.scala 361:21]
  wire  q_488_reset; // @[Decoupled.scala 361:21]
  wire  q_488_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_488_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_488_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_488_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_488_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_488_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_489_clock; // @[Decoupled.scala 361:21]
  wire  q_489_reset; // @[Decoupled.scala 361:21]
  wire  q_489_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_489_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_489_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_489_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_489_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_489_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_490_clock; // @[Decoupled.scala 361:21]
  wire  q_490_reset; // @[Decoupled.scala 361:21]
  wire  q_490_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_490_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_490_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_490_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_490_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_490_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_491_clock; // @[Decoupled.scala 361:21]
  wire  q_491_reset; // @[Decoupled.scala 361:21]
  wire  q_491_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_491_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_491_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_491_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_491_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_491_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_492_clock; // @[Decoupled.scala 361:21]
  wire  q_492_reset; // @[Decoupled.scala 361:21]
  wire  q_492_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_492_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_492_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_492_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_492_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_492_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_493_clock; // @[Decoupled.scala 361:21]
  wire  q_493_reset; // @[Decoupled.scala 361:21]
  wire  q_493_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_493_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_493_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_493_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_493_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_493_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_494_clock; // @[Decoupled.scala 361:21]
  wire  q_494_reset; // @[Decoupled.scala 361:21]
  wire  q_494_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_494_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_494_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_494_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_494_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_494_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_495_clock; // @[Decoupled.scala 361:21]
  wire  q_495_reset; // @[Decoupled.scala 361:21]
  wire  q_495_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_495_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_495_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_495_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_495_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_495_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_496_clock; // @[Decoupled.scala 361:21]
  wire  q_496_reset; // @[Decoupled.scala 361:21]
  wire  q_496_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_496_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_496_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_496_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_496_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_496_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_497_clock; // @[Decoupled.scala 361:21]
  wire  q_497_reset; // @[Decoupled.scala 361:21]
  wire  q_497_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_497_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_497_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_497_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_497_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_497_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_498_clock; // @[Decoupled.scala 361:21]
  wire  q_498_reset; // @[Decoupled.scala 361:21]
  wire  q_498_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_498_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_498_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_498_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_498_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_498_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_499_clock; // @[Decoupled.scala 361:21]
  wire  q_499_reset; // @[Decoupled.scala 361:21]
  wire  q_499_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_499_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_499_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_499_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_499_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_499_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_500_clock; // @[Decoupled.scala 361:21]
  wire  q_500_reset; // @[Decoupled.scala 361:21]
  wire  q_500_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_500_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_500_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_500_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_500_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_500_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_501_clock; // @[Decoupled.scala 361:21]
  wire  q_501_reset; // @[Decoupled.scala 361:21]
  wire  q_501_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_501_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_501_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_501_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_501_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_501_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_502_clock; // @[Decoupled.scala 361:21]
  wire  q_502_reset; // @[Decoupled.scala 361:21]
  wire  q_502_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_502_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_502_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_502_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_502_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_502_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_503_clock; // @[Decoupled.scala 361:21]
  wire  q_503_reset; // @[Decoupled.scala 361:21]
  wire  q_503_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_503_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_503_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_503_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_503_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_503_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_504_clock; // @[Decoupled.scala 361:21]
  wire  q_504_reset; // @[Decoupled.scala 361:21]
  wire  q_504_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_504_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_504_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_504_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_504_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_504_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_505_clock; // @[Decoupled.scala 361:21]
  wire  q_505_reset; // @[Decoupled.scala 361:21]
  wire  q_505_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_505_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_505_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_505_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_505_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_505_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_506_clock; // @[Decoupled.scala 361:21]
  wire  q_506_reset; // @[Decoupled.scala 361:21]
  wire  q_506_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_506_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_506_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_506_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_506_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_506_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_507_clock; // @[Decoupled.scala 361:21]
  wire  q_507_reset; // @[Decoupled.scala 361:21]
  wire  q_507_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_507_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_507_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_507_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_507_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_507_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_508_clock; // @[Decoupled.scala 361:21]
  wire  q_508_reset; // @[Decoupled.scala 361:21]
  wire  q_508_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_508_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_508_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_508_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_508_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_508_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_509_clock; // @[Decoupled.scala 361:21]
  wire  q_509_reset; // @[Decoupled.scala 361:21]
  wire  q_509_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_509_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_509_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_509_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_509_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_509_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_510_clock; // @[Decoupled.scala 361:21]
  wire  q_510_reset; // @[Decoupled.scala 361:21]
  wire  q_510_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_510_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_510_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_510_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_510_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_510_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_511_clock; // @[Decoupled.scala 361:21]
  wire  q_511_reset; // @[Decoupled.scala 361:21]
  wire  q_511_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_511_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_511_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_511_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_511_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_511_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_512_clock; // @[Decoupled.scala 361:21]
  wire  q_512_reset; // @[Decoupled.scala 361:21]
  wire  q_512_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_512_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_512_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_512_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_512_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_512_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_513_clock; // @[Decoupled.scala 361:21]
  wire  q_513_reset; // @[Decoupled.scala 361:21]
  wire  q_513_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_513_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_513_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_513_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_513_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_513_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_514_clock; // @[Decoupled.scala 361:21]
  wire  q_514_reset; // @[Decoupled.scala 361:21]
  wire  q_514_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_514_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_514_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_514_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_514_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_514_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_515_clock; // @[Decoupled.scala 361:21]
  wire  q_515_reset; // @[Decoupled.scala 361:21]
  wire  q_515_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_515_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_515_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_515_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_515_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_515_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_516_clock; // @[Decoupled.scala 361:21]
  wire  q_516_reset; // @[Decoupled.scala 361:21]
  wire  q_516_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_516_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_516_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_516_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_516_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_516_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_517_clock; // @[Decoupled.scala 361:21]
  wire  q_517_reset; // @[Decoupled.scala 361:21]
  wire  q_517_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_517_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_517_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_517_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_517_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_517_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_518_clock; // @[Decoupled.scala 361:21]
  wire  q_518_reset; // @[Decoupled.scala 361:21]
  wire  q_518_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_518_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_518_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_518_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_518_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_518_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_519_clock; // @[Decoupled.scala 361:21]
  wire  q_519_reset; // @[Decoupled.scala 361:21]
  wire  q_519_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_519_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_519_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_519_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_519_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_519_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_520_clock; // @[Decoupled.scala 361:21]
  wire  q_520_reset; // @[Decoupled.scala 361:21]
  wire  q_520_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_520_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_520_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_520_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_520_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_520_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_521_clock; // @[Decoupled.scala 361:21]
  wire  q_521_reset; // @[Decoupled.scala 361:21]
  wire  q_521_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_521_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_521_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_521_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_521_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_521_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_522_clock; // @[Decoupled.scala 361:21]
  wire  q_522_reset; // @[Decoupled.scala 361:21]
  wire  q_522_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_522_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_522_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_522_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_522_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_522_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_523_clock; // @[Decoupled.scala 361:21]
  wire  q_523_reset; // @[Decoupled.scala 361:21]
  wire  q_523_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_523_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_523_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_523_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_523_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_523_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_524_clock; // @[Decoupled.scala 361:21]
  wire  q_524_reset; // @[Decoupled.scala 361:21]
  wire  q_524_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_524_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_524_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_524_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_524_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_524_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_525_clock; // @[Decoupled.scala 361:21]
  wire  q_525_reset; // @[Decoupled.scala 361:21]
  wire  q_525_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_525_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_525_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_525_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_525_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_525_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_526_clock; // @[Decoupled.scala 361:21]
  wire  q_526_reset; // @[Decoupled.scala 361:21]
  wire  q_526_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_526_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_526_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_526_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_526_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_526_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_527_clock; // @[Decoupled.scala 361:21]
  wire  q_527_reset; // @[Decoupled.scala 361:21]
  wire  q_527_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_527_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_527_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_527_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_527_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_527_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_528_clock; // @[Decoupled.scala 361:21]
  wire  q_528_reset; // @[Decoupled.scala 361:21]
  wire  q_528_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_528_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_528_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_528_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_528_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_528_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_529_clock; // @[Decoupled.scala 361:21]
  wire  q_529_reset; // @[Decoupled.scala 361:21]
  wire  q_529_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_529_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_529_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_529_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_529_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_529_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_530_clock; // @[Decoupled.scala 361:21]
  wire  q_530_reset; // @[Decoupled.scala 361:21]
  wire  q_530_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_530_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_530_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_530_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_530_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_530_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_531_clock; // @[Decoupled.scala 361:21]
  wire  q_531_reset; // @[Decoupled.scala 361:21]
  wire  q_531_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_531_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_531_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_531_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_531_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_531_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_532_clock; // @[Decoupled.scala 361:21]
  wire  q_532_reset; // @[Decoupled.scala 361:21]
  wire  q_532_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_532_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_532_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_532_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_532_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_532_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_533_clock; // @[Decoupled.scala 361:21]
  wire  q_533_reset; // @[Decoupled.scala 361:21]
  wire  q_533_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_533_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_533_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_533_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_533_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_533_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_534_clock; // @[Decoupled.scala 361:21]
  wire  q_534_reset; // @[Decoupled.scala 361:21]
  wire  q_534_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_534_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_534_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_534_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_534_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_534_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_535_clock; // @[Decoupled.scala 361:21]
  wire  q_535_reset; // @[Decoupled.scala 361:21]
  wire  q_535_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_535_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_535_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_535_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_535_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_535_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_536_clock; // @[Decoupled.scala 361:21]
  wire  q_536_reset; // @[Decoupled.scala 361:21]
  wire  q_536_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_536_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_536_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_536_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_536_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_536_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_537_clock; // @[Decoupled.scala 361:21]
  wire  q_537_reset; // @[Decoupled.scala 361:21]
  wire  q_537_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_537_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_537_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_537_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_537_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_537_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_538_clock; // @[Decoupled.scala 361:21]
  wire  q_538_reset; // @[Decoupled.scala 361:21]
  wire  q_538_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_538_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_538_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_538_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_538_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_538_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_539_clock; // @[Decoupled.scala 361:21]
  wire  q_539_reset; // @[Decoupled.scala 361:21]
  wire  q_539_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_539_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_539_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_539_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_539_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_539_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_540_clock; // @[Decoupled.scala 361:21]
  wire  q_540_reset; // @[Decoupled.scala 361:21]
  wire  q_540_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_540_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_540_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_540_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_540_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_540_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_541_clock; // @[Decoupled.scala 361:21]
  wire  q_541_reset; // @[Decoupled.scala 361:21]
  wire  q_541_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_541_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_541_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_541_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_541_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_541_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_542_clock; // @[Decoupled.scala 361:21]
  wire  q_542_reset; // @[Decoupled.scala 361:21]
  wire  q_542_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_542_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_542_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_542_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_542_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_542_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_543_clock; // @[Decoupled.scala 361:21]
  wire  q_543_reset; // @[Decoupled.scala 361:21]
  wire  q_543_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_543_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_543_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_543_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_543_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_543_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_544_clock; // @[Decoupled.scala 361:21]
  wire  q_544_reset; // @[Decoupled.scala 361:21]
  wire  q_544_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_544_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_544_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_544_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_544_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_544_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_545_clock; // @[Decoupled.scala 361:21]
  wire  q_545_reset; // @[Decoupled.scala 361:21]
  wire  q_545_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_545_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_545_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_545_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_545_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_545_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_546_clock; // @[Decoupled.scala 361:21]
  wire  q_546_reset; // @[Decoupled.scala 361:21]
  wire  q_546_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_546_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_546_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_546_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_546_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_546_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_547_clock; // @[Decoupled.scala 361:21]
  wire  q_547_reset; // @[Decoupled.scala 361:21]
  wire  q_547_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_547_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_547_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_547_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_547_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_547_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_548_clock; // @[Decoupled.scala 361:21]
  wire  q_548_reset; // @[Decoupled.scala 361:21]
  wire  q_548_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_548_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_548_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_548_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_548_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_548_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_549_clock; // @[Decoupled.scala 361:21]
  wire  q_549_reset; // @[Decoupled.scala 361:21]
  wire  q_549_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_549_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_549_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_549_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_549_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_549_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_550_clock; // @[Decoupled.scala 361:21]
  wire  q_550_reset; // @[Decoupled.scala 361:21]
  wire  q_550_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_550_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_550_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_550_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_550_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_550_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_551_clock; // @[Decoupled.scala 361:21]
  wire  q_551_reset; // @[Decoupled.scala 361:21]
  wire  q_551_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_551_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_551_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_551_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_551_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_551_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_552_clock; // @[Decoupled.scala 361:21]
  wire  q_552_reset; // @[Decoupled.scala 361:21]
  wire  q_552_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_552_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_552_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_552_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_552_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_552_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_553_clock; // @[Decoupled.scala 361:21]
  wire  q_553_reset; // @[Decoupled.scala 361:21]
  wire  q_553_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_553_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_553_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_553_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_553_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_553_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_554_clock; // @[Decoupled.scala 361:21]
  wire  q_554_reset; // @[Decoupled.scala 361:21]
  wire  q_554_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_554_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_554_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_554_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_554_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_554_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_555_clock; // @[Decoupled.scala 361:21]
  wire  q_555_reset; // @[Decoupled.scala 361:21]
  wire  q_555_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_555_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_555_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_555_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_555_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_555_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_556_clock; // @[Decoupled.scala 361:21]
  wire  q_556_reset; // @[Decoupled.scala 361:21]
  wire  q_556_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_556_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_556_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_556_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_556_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_556_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_557_clock; // @[Decoupled.scala 361:21]
  wire  q_557_reset; // @[Decoupled.scala 361:21]
  wire  q_557_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_557_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_557_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_557_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_557_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_557_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_558_clock; // @[Decoupled.scala 361:21]
  wire  q_558_reset; // @[Decoupled.scala 361:21]
  wire  q_558_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_558_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_558_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_558_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_558_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_558_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_559_clock; // @[Decoupled.scala 361:21]
  wire  q_559_reset; // @[Decoupled.scala 361:21]
  wire  q_559_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_559_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_559_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_559_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_559_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_559_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_560_clock; // @[Decoupled.scala 361:21]
  wire  q_560_reset; // @[Decoupled.scala 361:21]
  wire  q_560_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_560_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_560_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_560_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_560_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_560_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_561_clock; // @[Decoupled.scala 361:21]
  wire  q_561_reset; // @[Decoupled.scala 361:21]
  wire  q_561_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_561_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_561_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_561_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_561_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_561_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_562_clock; // @[Decoupled.scala 361:21]
  wire  q_562_reset; // @[Decoupled.scala 361:21]
  wire  q_562_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_562_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_562_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_562_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_562_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_562_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_563_clock; // @[Decoupled.scala 361:21]
  wire  q_563_reset; // @[Decoupled.scala 361:21]
  wire  q_563_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_563_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_563_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_563_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_563_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_563_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_564_clock; // @[Decoupled.scala 361:21]
  wire  q_564_reset; // @[Decoupled.scala 361:21]
  wire  q_564_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_564_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_564_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_564_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_564_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_564_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_565_clock; // @[Decoupled.scala 361:21]
  wire  q_565_reset; // @[Decoupled.scala 361:21]
  wire  q_565_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_565_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_565_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_565_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_565_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_565_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_566_clock; // @[Decoupled.scala 361:21]
  wire  q_566_reset; // @[Decoupled.scala 361:21]
  wire  q_566_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_566_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_566_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_566_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_566_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_566_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_567_clock; // @[Decoupled.scala 361:21]
  wire  q_567_reset; // @[Decoupled.scala 361:21]
  wire  q_567_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_567_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_567_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_567_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_567_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_567_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_568_clock; // @[Decoupled.scala 361:21]
  wire  q_568_reset; // @[Decoupled.scala 361:21]
  wire  q_568_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_568_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_568_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_568_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_568_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_568_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_569_clock; // @[Decoupled.scala 361:21]
  wire  q_569_reset; // @[Decoupled.scala 361:21]
  wire  q_569_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_569_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_569_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_569_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_569_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_569_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_570_clock; // @[Decoupled.scala 361:21]
  wire  q_570_reset; // @[Decoupled.scala 361:21]
  wire  q_570_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_570_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_570_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_570_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_570_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_570_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_571_clock; // @[Decoupled.scala 361:21]
  wire  q_571_reset; // @[Decoupled.scala 361:21]
  wire  q_571_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_571_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_571_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_571_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_571_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_571_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_572_clock; // @[Decoupled.scala 361:21]
  wire  q_572_reset; // @[Decoupled.scala 361:21]
  wire  q_572_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_572_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_572_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_572_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_572_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_572_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_573_clock; // @[Decoupled.scala 361:21]
  wire  q_573_reset; // @[Decoupled.scala 361:21]
  wire  q_573_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_573_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_573_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_573_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_573_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_573_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_574_clock; // @[Decoupled.scala 361:21]
  wire  q_574_reset; // @[Decoupled.scala 361:21]
  wire  q_574_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_574_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_574_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_574_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_574_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_574_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_575_clock; // @[Decoupled.scala 361:21]
  wire  q_575_reset; // @[Decoupled.scala 361:21]
  wire  q_575_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_575_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_575_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_575_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_575_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_575_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_576_clock; // @[Decoupled.scala 361:21]
  wire  q_576_reset; // @[Decoupled.scala 361:21]
  wire  q_576_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_576_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_576_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_576_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_576_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_576_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_577_clock; // @[Decoupled.scala 361:21]
  wire  q_577_reset; // @[Decoupled.scala 361:21]
  wire  q_577_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_577_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_577_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_577_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_577_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_577_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_578_clock; // @[Decoupled.scala 361:21]
  wire  q_578_reset; // @[Decoupled.scala 361:21]
  wire  q_578_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_578_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_578_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_578_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_578_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_578_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_579_clock; // @[Decoupled.scala 361:21]
  wire  q_579_reset; // @[Decoupled.scala 361:21]
  wire  q_579_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_579_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_579_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_579_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_579_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_579_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_580_clock; // @[Decoupled.scala 361:21]
  wire  q_580_reset; // @[Decoupled.scala 361:21]
  wire  q_580_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_580_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_580_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_580_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_580_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_580_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_581_clock; // @[Decoupled.scala 361:21]
  wire  q_581_reset; // @[Decoupled.scala 361:21]
  wire  q_581_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_581_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_581_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_581_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_581_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_581_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_582_clock; // @[Decoupled.scala 361:21]
  wire  q_582_reset; // @[Decoupled.scala 361:21]
  wire  q_582_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_582_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_582_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_582_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_582_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_582_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_583_clock; // @[Decoupled.scala 361:21]
  wire  q_583_reset; // @[Decoupled.scala 361:21]
  wire  q_583_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_583_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_583_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_583_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_583_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_583_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_584_clock; // @[Decoupled.scala 361:21]
  wire  q_584_reset; // @[Decoupled.scala 361:21]
  wire  q_584_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_584_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_584_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_584_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_584_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_584_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_585_clock; // @[Decoupled.scala 361:21]
  wire  q_585_reset; // @[Decoupled.scala 361:21]
  wire  q_585_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_585_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_585_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_585_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_585_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_585_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_586_clock; // @[Decoupled.scala 361:21]
  wire  q_586_reset; // @[Decoupled.scala 361:21]
  wire  q_586_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_586_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_586_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_586_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_586_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_586_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_587_clock; // @[Decoupled.scala 361:21]
  wire  q_587_reset; // @[Decoupled.scala 361:21]
  wire  q_587_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_587_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_587_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_587_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_587_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_587_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_588_clock; // @[Decoupled.scala 361:21]
  wire  q_588_reset; // @[Decoupled.scala 361:21]
  wire  q_588_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_588_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_588_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_588_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_588_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_588_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_589_clock; // @[Decoupled.scala 361:21]
  wire  q_589_reset; // @[Decoupled.scala 361:21]
  wire  q_589_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_589_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_589_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_589_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_589_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_589_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_590_clock; // @[Decoupled.scala 361:21]
  wire  q_590_reset; // @[Decoupled.scala 361:21]
  wire  q_590_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_590_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_590_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_590_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_590_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_590_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_591_clock; // @[Decoupled.scala 361:21]
  wire  q_591_reset; // @[Decoupled.scala 361:21]
  wire  q_591_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_591_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_591_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_591_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_591_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_591_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_592_clock; // @[Decoupled.scala 361:21]
  wire  q_592_reset; // @[Decoupled.scala 361:21]
  wire  q_592_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_592_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_592_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_592_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_592_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_592_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_593_clock; // @[Decoupled.scala 361:21]
  wire  q_593_reset; // @[Decoupled.scala 361:21]
  wire  q_593_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_593_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_593_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_593_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_593_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_593_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_594_clock; // @[Decoupled.scala 361:21]
  wire  q_594_reset; // @[Decoupled.scala 361:21]
  wire  q_594_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_594_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_594_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_594_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_594_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_594_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_595_clock; // @[Decoupled.scala 361:21]
  wire  q_595_reset; // @[Decoupled.scala 361:21]
  wire  q_595_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_595_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_595_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_595_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_595_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_595_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_596_clock; // @[Decoupled.scala 361:21]
  wire  q_596_reset; // @[Decoupled.scala 361:21]
  wire  q_596_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_596_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_596_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_596_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_596_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_596_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_597_clock; // @[Decoupled.scala 361:21]
  wire  q_597_reset; // @[Decoupled.scala 361:21]
  wire  q_597_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_597_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_597_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_597_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_597_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_597_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_598_clock; // @[Decoupled.scala 361:21]
  wire  q_598_reset; // @[Decoupled.scala 361:21]
  wire  q_598_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_598_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_598_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_598_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_598_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_598_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_599_clock; // @[Decoupled.scala 361:21]
  wire  q_599_reset; // @[Decoupled.scala 361:21]
  wire  q_599_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_599_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_599_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_599_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_599_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_599_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_600_clock; // @[Decoupled.scala 361:21]
  wire  q_600_reset; // @[Decoupled.scala 361:21]
  wire  q_600_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_600_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_600_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_600_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_600_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_600_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_601_clock; // @[Decoupled.scala 361:21]
  wire  q_601_reset; // @[Decoupled.scala 361:21]
  wire  q_601_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_601_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_601_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_601_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_601_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_601_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_602_clock; // @[Decoupled.scala 361:21]
  wire  q_602_reset; // @[Decoupled.scala 361:21]
  wire  q_602_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_602_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_602_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_602_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_602_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_602_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_603_clock; // @[Decoupled.scala 361:21]
  wire  q_603_reset; // @[Decoupled.scala 361:21]
  wire  q_603_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_603_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_603_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_603_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_603_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_603_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_604_clock; // @[Decoupled.scala 361:21]
  wire  q_604_reset; // @[Decoupled.scala 361:21]
  wire  q_604_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_604_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_604_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_604_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_604_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_604_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_605_clock; // @[Decoupled.scala 361:21]
  wire  q_605_reset; // @[Decoupled.scala 361:21]
  wire  q_605_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_605_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_605_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_605_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_605_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_605_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_606_clock; // @[Decoupled.scala 361:21]
  wire  q_606_reset; // @[Decoupled.scala 361:21]
  wire  q_606_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_606_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_606_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_606_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_606_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_606_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_607_clock; // @[Decoupled.scala 361:21]
  wire  q_607_reset; // @[Decoupled.scala 361:21]
  wire  q_607_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_607_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_607_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_607_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_607_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_607_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_608_clock; // @[Decoupled.scala 361:21]
  wire  q_608_reset; // @[Decoupled.scala 361:21]
  wire  q_608_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_608_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_608_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_608_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_608_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_608_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_609_clock; // @[Decoupled.scala 361:21]
  wire  q_609_reset; // @[Decoupled.scala 361:21]
  wire  q_609_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_609_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_609_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_609_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_609_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_609_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_610_clock; // @[Decoupled.scala 361:21]
  wire  q_610_reset; // @[Decoupled.scala 361:21]
  wire  q_610_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_610_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_610_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_610_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_610_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_610_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_611_clock; // @[Decoupled.scala 361:21]
  wire  q_611_reset; // @[Decoupled.scala 361:21]
  wire  q_611_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_611_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_611_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_611_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_611_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_611_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_612_clock; // @[Decoupled.scala 361:21]
  wire  q_612_reset; // @[Decoupled.scala 361:21]
  wire  q_612_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_612_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_612_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_612_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_612_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_612_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_613_clock; // @[Decoupled.scala 361:21]
  wire  q_613_reset; // @[Decoupled.scala 361:21]
  wire  q_613_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_613_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_613_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_613_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_613_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_613_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_614_clock; // @[Decoupled.scala 361:21]
  wire  q_614_reset; // @[Decoupled.scala 361:21]
  wire  q_614_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_614_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_614_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_614_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_614_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_614_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_615_clock; // @[Decoupled.scala 361:21]
  wire  q_615_reset; // @[Decoupled.scala 361:21]
  wire  q_615_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_615_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_615_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_615_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_615_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_615_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_616_clock; // @[Decoupled.scala 361:21]
  wire  q_616_reset; // @[Decoupled.scala 361:21]
  wire  q_616_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_616_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_616_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_616_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_616_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_616_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_617_clock; // @[Decoupled.scala 361:21]
  wire  q_617_reset; // @[Decoupled.scala 361:21]
  wire  q_617_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_617_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_617_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_617_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_617_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_617_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_618_clock; // @[Decoupled.scala 361:21]
  wire  q_618_reset; // @[Decoupled.scala 361:21]
  wire  q_618_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_618_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_618_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_618_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_618_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_618_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_619_clock; // @[Decoupled.scala 361:21]
  wire  q_619_reset; // @[Decoupled.scala 361:21]
  wire  q_619_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_619_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_619_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_619_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_619_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_619_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_620_clock; // @[Decoupled.scala 361:21]
  wire  q_620_reset; // @[Decoupled.scala 361:21]
  wire  q_620_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_620_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_620_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_620_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_620_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_620_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_621_clock; // @[Decoupled.scala 361:21]
  wire  q_621_reset; // @[Decoupled.scala 361:21]
  wire  q_621_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_621_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_621_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_621_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_621_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_621_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_622_clock; // @[Decoupled.scala 361:21]
  wire  q_622_reset; // @[Decoupled.scala 361:21]
  wire  q_622_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_622_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_622_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_622_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_622_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_622_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_623_clock; // @[Decoupled.scala 361:21]
  wire  q_623_reset; // @[Decoupled.scala 361:21]
  wire  q_623_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_623_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_623_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_623_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_623_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_623_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_624_clock; // @[Decoupled.scala 361:21]
  wire  q_624_reset; // @[Decoupled.scala 361:21]
  wire  q_624_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_624_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_624_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_624_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_624_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_624_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_625_clock; // @[Decoupled.scala 361:21]
  wire  q_625_reset; // @[Decoupled.scala 361:21]
  wire  q_625_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_625_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_625_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_625_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_625_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_625_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_626_clock; // @[Decoupled.scala 361:21]
  wire  q_626_reset; // @[Decoupled.scala 361:21]
  wire  q_626_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_626_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_626_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_626_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_626_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_626_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_627_clock; // @[Decoupled.scala 361:21]
  wire  q_627_reset; // @[Decoupled.scala 361:21]
  wire  q_627_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_627_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_627_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_627_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_627_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_627_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_628_clock; // @[Decoupled.scala 361:21]
  wire  q_628_reset; // @[Decoupled.scala 361:21]
  wire  q_628_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_628_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_628_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_628_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_628_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_628_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_629_clock; // @[Decoupled.scala 361:21]
  wire  q_629_reset; // @[Decoupled.scala 361:21]
  wire  q_629_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_629_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_629_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_629_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_629_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_629_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_630_clock; // @[Decoupled.scala 361:21]
  wire  q_630_reset; // @[Decoupled.scala 361:21]
  wire  q_630_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_630_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_630_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_630_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_630_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_630_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_631_clock; // @[Decoupled.scala 361:21]
  wire  q_631_reset; // @[Decoupled.scala 361:21]
  wire  q_631_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_631_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_631_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_631_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_631_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_631_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_632_clock; // @[Decoupled.scala 361:21]
  wire  q_632_reset; // @[Decoupled.scala 361:21]
  wire  q_632_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_632_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_632_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_632_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_632_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_632_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_633_clock; // @[Decoupled.scala 361:21]
  wire  q_633_reset; // @[Decoupled.scala 361:21]
  wire  q_633_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_633_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_633_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_633_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_633_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_633_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_634_clock; // @[Decoupled.scala 361:21]
  wire  q_634_reset; // @[Decoupled.scala 361:21]
  wire  q_634_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_634_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_634_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_634_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_634_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_634_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_635_clock; // @[Decoupled.scala 361:21]
  wire  q_635_reset; // @[Decoupled.scala 361:21]
  wire  q_635_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_635_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_635_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_635_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_635_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_635_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_636_clock; // @[Decoupled.scala 361:21]
  wire  q_636_reset; // @[Decoupled.scala 361:21]
  wire  q_636_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_636_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_636_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_636_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_636_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_636_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_637_clock; // @[Decoupled.scala 361:21]
  wire  q_637_reset; // @[Decoupled.scala 361:21]
  wire  q_637_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_637_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_637_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_637_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_637_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_637_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_638_clock; // @[Decoupled.scala 361:21]
  wire  q_638_reset; // @[Decoupled.scala 361:21]
  wire  q_638_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_638_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_638_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_638_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_638_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_638_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_639_clock; // @[Decoupled.scala 361:21]
  wire  q_639_reset; // @[Decoupled.scala 361:21]
  wire  q_639_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_639_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_639_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_639_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_639_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_639_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_640_clock; // @[Decoupled.scala 361:21]
  wire  q_640_reset; // @[Decoupled.scala 361:21]
  wire  q_640_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_640_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_640_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_640_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_640_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_640_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_641_clock; // @[Decoupled.scala 361:21]
  wire  q_641_reset; // @[Decoupled.scala 361:21]
  wire  q_641_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_641_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_641_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_641_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_641_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_641_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_642_clock; // @[Decoupled.scala 361:21]
  wire  q_642_reset; // @[Decoupled.scala 361:21]
  wire  q_642_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_642_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_642_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_642_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_642_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_642_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_643_clock; // @[Decoupled.scala 361:21]
  wire  q_643_reset; // @[Decoupled.scala 361:21]
  wire  q_643_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_643_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_643_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_643_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_643_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_643_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_644_clock; // @[Decoupled.scala 361:21]
  wire  q_644_reset; // @[Decoupled.scala 361:21]
  wire  q_644_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_644_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_644_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_644_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_644_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_644_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_645_clock; // @[Decoupled.scala 361:21]
  wire  q_645_reset; // @[Decoupled.scala 361:21]
  wire  q_645_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_645_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_645_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_645_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_645_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_645_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_646_clock; // @[Decoupled.scala 361:21]
  wire  q_646_reset; // @[Decoupled.scala 361:21]
  wire  q_646_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_646_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_646_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_646_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_646_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_646_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_647_clock; // @[Decoupled.scala 361:21]
  wire  q_647_reset; // @[Decoupled.scala 361:21]
  wire  q_647_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_647_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_647_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_647_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_647_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_647_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_648_clock; // @[Decoupled.scala 361:21]
  wire  q_648_reset; // @[Decoupled.scala 361:21]
  wire  q_648_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_648_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_648_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_648_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_648_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_648_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_649_clock; // @[Decoupled.scala 361:21]
  wire  q_649_reset; // @[Decoupled.scala 361:21]
  wire  q_649_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_649_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_649_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_649_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_649_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_649_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_650_clock; // @[Decoupled.scala 361:21]
  wire  q_650_reset; // @[Decoupled.scala 361:21]
  wire  q_650_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_650_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_650_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_650_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_650_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_650_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_651_clock; // @[Decoupled.scala 361:21]
  wire  q_651_reset; // @[Decoupled.scala 361:21]
  wire  q_651_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_651_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_651_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_651_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_651_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_651_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_652_clock; // @[Decoupled.scala 361:21]
  wire  q_652_reset; // @[Decoupled.scala 361:21]
  wire  q_652_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_652_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_652_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_652_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_652_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_652_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_653_clock; // @[Decoupled.scala 361:21]
  wire  q_653_reset; // @[Decoupled.scala 361:21]
  wire  q_653_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_653_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_653_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_653_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_653_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_653_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_654_clock; // @[Decoupled.scala 361:21]
  wire  q_654_reset; // @[Decoupled.scala 361:21]
  wire  q_654_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_654_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_654_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_654_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_654_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_654_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_655_clock; // @[Decoupled.scala 361:21]
  wire  q_655_reset; // @[Decoupled.scala 361:21]
  wire  q_655_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_655_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_655_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_655_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_655_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_655_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_656_clock; // @[Decoupled.scala 361:21]
  wire  q_656_reset; // @[Decoupled.scala 361:21]
  wire  q_656_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_656_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_656_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_656_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_656_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_656_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_657_clock; // @[Decoupled.scala 361:21]
  wire  q_657_reset; // @[Decoupled.scala 361:21]
  wire  q_657_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_657_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_657_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_657_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_657_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_657_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_658_clock; // @[Decoupled.scala 361:21]
  wire  q_658_reset; // @[Decoupled.scala 361:21]
  wire  q_658_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_658_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_658_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_658_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_658_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_658_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_659_clock; // @[Decoupled.scala 361:21]
  wire  q_659_reset; // @[Decoupled.scala 361:21]
  wire  q_659_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_659_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_659_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_659_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_659_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_659_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_660_clock; // @[Decoupled.scala 361:21]
  wire  q_660_reset; // @[Decoupled.scala 361:21]
  wire  q_660_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_660_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_660_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_660_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_660_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_660_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_661_clock; // @[Decoupled.scala 361:21]
  wire  q_661_reset; // @[Decoupled.scala 361:21]
  wire  q_661_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_661_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_661_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_661_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_661_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_661_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_662_clock; // @[Decoupled.scala 361:21]
  wire  q_662_reset; // @[Decoupled.scala 361:21]
  wire  q_662_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_662_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_662_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_662_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_662_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_662_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_663_clock; // @[Decoupled.scala 361:21]
  wire  q_663_reset; // @[Decoupled.scala 361:21]
  wire  q_663_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_663_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_663_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_663_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_663_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_663_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_664_clock; // @[Decoupled.scala 361:21]
  wire  q_664_reset; // @[Decoupled.scala 361:21]
  wire  q_664_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_664_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_664_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_664_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_664_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_664_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_665_clock; // @[Decoupled.scala 361:21]
  wire  q_665_reset; // @[Decoupled.scala 361:21]
  wire  q_665_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_665_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_665_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_665_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_665_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_665_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_666_clock; // @[Decoupled.scala 361:21]
  wire  q_666_reset; // @[Decoupled.scala 361:21]
  wire  q_666_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_666_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_666_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_666_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_666_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_666_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_667_clock; // @[Decoupled.scala 361:21]
  wire  q_667_reset; // @[Decoupled.scala 361:21]
  wire  q_667_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_667_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_667_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_667_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_667_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_667_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_668_clock; // @[Decoupled.scala 361:21]
  wire  q_668_reset; // @[Decoupled.scala 361:21]
  wire  q_668_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_668_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_668_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_668_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_668_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_668_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_669_clock; // @[Decoupled.scala 361:21]
  wire  q_669_reset; // @[Decoupled.scala 361:21]
  wire  q_669_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_669_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_669_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_669_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_669_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_669_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_670_clock; // @[Decoupled.scala 361:21]
  wire  q_670_reset; // @[Decoupled.scala 361:21]
  wire  q_670_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_670_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_670_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_670_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_670_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_670_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_671_clock; // @[Decoupled.scala 361:21]
  wire  q_671_reset; // @[Decoupled.scala 361:21]
  wire  q_671_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_671_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_671_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_671_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_671_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_671_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_672_clock; // @[Decoupled.scala 361:21]
  wire  q_672_reset; // @[Decoupled.scala 361:21]
  wire  q_672_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_672_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_672_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_672_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_672_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_672_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_673_clock; // @[Decoupled.scala 361:21]
  wire  q_673_reset; // @[Decoupled.scala 361:21]
  wire  q_673_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_673_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_673_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_673_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_673_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_673_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_674_clock; // @[Decoupled.scala 361:21]
  wire  q_674_reset; // @[Decoupled.scala 361:21]
  wire  q_674_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_674_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_674_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_674_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_674_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_674_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_675_clock; // @[Decoupled.scala 361:21]
  wire  q_675_reset; // @[Decoupled.scala 361:21]
  wire  q_675_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_675_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_675_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_675_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_675_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_675_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_676_clock; // @[Decoupled.scala 361:21]
  wire  q_676_reset; // @[Decoupled.scala 361:21]
  wire  q_676_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_676_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_676_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_676_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_676_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_676_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_677_clock; // @[Decoupled.scala 361:21]
  wire  q_677_reset; // @[Decoupled.scala 361:21]
  wire  q_677_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_677_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_677_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_677_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_677_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_677_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_678_clock; // @[Decoupled.scala 361:21]
  wire  q_678_reset; // @[Decoupled.scala 361:21]
  wire  q_678_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_678_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_678_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_678_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_678_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_678_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_679_clock; // @[Decoupled.scala 361:21]
  wire  q_679_reset; // @[Decoupled.scala 361:21]
  wire  q_679_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_679_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_679_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_679_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_679_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_679_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_680_clock; // @[Decoupled.scala 361:21]
  wire  q_680_reset; // @[Decoupled.scala 361:21]
  wire  q_680_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_680_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_680_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_680_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_680_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_680_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_681_clock; // @[Decoupled.scala 361:21]
  wire  q_681_reset; // @[Decoupled.scala 361:21]
  wire  q_681_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_681_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_681_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_681_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_681_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_681_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_682_clock; // @[Decoupled.scala 361:21]
  wire  q_682_reset; // @[Decoupled.scala 361:21]
  wire  q_682_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_682_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_682_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_682_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_682_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_682_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_683_clock; // @[Decoupled.scala 361:21]
  wire  q_683_reset; // @[Decoupled.scala 361:21]
  wire  q_683_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_683_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_683_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_683_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_683_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_683_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_684_clock; // @[Decoupled.scala 361:21]
  wire  q_684_reset; // @[Decoupled.scala 361:21]
  wire  q_684_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_684_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_684_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_684_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_684_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_684_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_685_clock; // @[Decoupled.scala 361:21]
  wire  q_685_reset; // @[Decoupled.scala 361:21]
  wire  q_685_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_685_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_685_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_685_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_685_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_685_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_686_clock; // @[Decoupled.scala 361:21]
  wire  q_686_reset; // @[Decoupled.scala 361:21]
  wire  q_686_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_686_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_686_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_686_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_686_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_686_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_687_clock; // @[Decoupled.scala 361:21]
  wire  q_687_reset; // @[Decoupled.scala 361:21]
  wire  q_687_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_687_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_687_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_687_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_687_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_687_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_688_clock; // @[Decoupled.scala 361:21]
  wire  q_688_reset; // @[Decoupled.scala 361:21]
  wire  q_688_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_688_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_688_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_688_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_688_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_688_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_689_clock; // @[Decoupled.scala 361:21]
  wire  q_689_reset; // @[Decoupled.scala 361:21]
  wire  q_689_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_689_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_689_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_689_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_689_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_689_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_690_clock; // @[Decoupled.scala 361:21]
  wire  q_690_reset; // @[Decoupled.scala 361:21]
  wire  q_690_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_690_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_690_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_690_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_690_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_690_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_691_clock; // @[Decoupled.scala 361:21]
  wire  q_691_reset; // @[Decoupled.scala 361:21]
  wire  q_691_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_691_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_691_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_691_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_691_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_691_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_692_clock; // @[Decoupled.scala 361:21]
  wire  q_692_reset; // @[Decoupled.scala 361:21]
  wire  q_692_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_692_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_692_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_692_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_692_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_692_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_693_clock; // @[Decoupled.scala 361:21]
  wire  q_693_reset; // @[Decoupled.scala 361:21]
  wire  q_693_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_693_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_693_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_693_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_693_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_693_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_694_clock; // @[Decoupled.scala 361:21]
  wire  q_694_reset; // @[Decoupled.scala 361:21]
  wire  q_694_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_694_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_694_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_694_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_694_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_694_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_695_clock; // @[Decoupled.scala 361:21]
  wire  q_695_reset; // @[Decoupled.scala 361:21]
  wire  q_695_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_695_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_695_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_695_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_695_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_695_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_696_clock; // @[Decoupled.scala 361:21]
  wire  q_696_reset; // @[Decoupled.scala 361:21]
  wire  q_696_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_696_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_696_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_696_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_696_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_696_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_697_clock; // @[Decoupled.scala 361:21]
  wire  q_697_reset; // @[Decoupled.scala 361:21]
  wire  q_697_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_697_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_697_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_697_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_697_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_697_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_698_clock; // @[Decoupled.scala 361:21]
  wire  q_698_reset; // @[Decoupled.scala 361:21]
  wire  q_698_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_698_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_698_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_698_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_698_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_698_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_699_clock; // @[Decoupled.scala 361:21]
  wire  q_699_reset; // @[Decoupled.scala 361:21]
  wire  q_699_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_699_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_699_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_699_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_699_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_699_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_700_clock; // @[Decoupled.scala 361:21]
  wire  q_700_reset; // @[Decoupled.scala 361:21]
  wire  q_700_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_700_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_700_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_700_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_700_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_700_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_701_clock; // @[Decoupled.scala 361:21]
  wire  q_701_reset; // @[Decoupled.scala 361:21]
  wire  q_701_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_701_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_701_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_701_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_701_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_701_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_702_clock; // @[Decoupled.scala 361:21]
  wire  q_702_reset; // @[Decoupled.scala 361:21]
  wire  q_702_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_702_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_702_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_702_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_702_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_702_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_703_clock; // @[Decoupled.scala 361:21]
  wire  q_703_reset; // @[Decoupled.scala 361:21]
  wire  q_703_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_703_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_703_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_703_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_703_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_703_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_704_clock; // @[Decoupled.scala 361:21]
  wire  q_704_reset; // @[Decoupled.scala 361:21]
  wire  q_704_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_704_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_704_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_704_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_704_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_704_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_705_clock; // @[Decoupled.scala 361:21]
  wire  q_705_reset; // @[Decoupled.scala 361:21]
  wire  q_705_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_705_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_705_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_705_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_705_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_705_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_706_clock; // @[Decoupled.scala 361:21]
  wire  q_706_reset; // @[Decoupled.scala 361:21]
  wire  q_706_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_706_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_706_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_706_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_706_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_706_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_707_clock; // @[Decoupled.scala 361:21]
  wire  q_707_reset; // @[Decoupled.scala 361:21]
  wire  q_707_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_707_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_707_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_707_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_707_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_707_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_708_clock; // @[Decoupled.scala 361:21]
  wire  q_708_reset; // @[Decoupled.scala 361:21]
  wire  q_708_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_708_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_708_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_708_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_708_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_708_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_709_clock; // @[Decoupled.scala 361:21]
  wire  q_709_reset; // @[Decoupled.scala 361:21]
  wire  q_709_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_709_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_709_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_709_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_709_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_709_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_710_clock; // @[Decoupled.scala 361:21]
  wire  q_710_reset; // @[Decoupled.scala 361:21]
  wire  q_710_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_710_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_710_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_710_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_710_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_710_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_711_clock; // @[Decoupled.scala 361:21]
  wire  q_711_reset; // @[Decoupled.scala 361:21]
  wire  q_711_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_711_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_711_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_711_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_711_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_711_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_712_clock; // @[Decoupled.scala 361:21]
  wire  q_712_reset; // @[Decoupled.scala 361:21]
  wire  q_712_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_712_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_712_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_712_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_712_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_712_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_713_clock; // @[Decoupled.scala 361:21]
  wire  q_713_reset; // @[Decoupled.scala 361:21]
  wire  q_713_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_713_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_713_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_713_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_713_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_713_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_714_clock; // @[Decoupled.scala 361:21]
  wire  q_714_reset; // @[Decoupled.scala 361:21]
  wire  q_714_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_714_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_714_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_714_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_714_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_714_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_715_clock; // @[Decoupled.scala 361:21]
  wire  q_715_reset; // @[Decoupled.scala 361:21]
  wire  q_715_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_715_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_715_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_715_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_715_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_715_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_716_clock; // @[Decoupled.scala 361:21]
  wire  q_716_reset; // @[Decoupled.scala 361:21]
  wire  q_716_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_716_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_716_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_716_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_716_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_716_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_717_clock; // @[Decoupled.scala 361:21]
  wire  q_717_reset; // @[Decoupled.scala 361:21]
  wire  q_717_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_717_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_717_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_717_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_717_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_717_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_718_clock; // @[Decoupled.scala 361:21]
  wire  q_718_reset; // @[Decoupled.scala 361:21]
  wire  q_718_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_718_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_718_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_718_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_718_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_718_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_719_clock; // @[Decoupled.scala 361:21]
  wire  q_719_reset; // @[Decoupled.scala 361:21]
  wire  q_719_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_719_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_719_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_719_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_719_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_719_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_720_clock; // @[Decoupled.scala 361:21]
  wire  q_720_reset; // @[Decoupled.scala 361:21]
  wire  q_720_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_720_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_720_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_720_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_720_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_720_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_721_clock; // @[Decoupled.scala 361:21]
  wire  q_721_reset; // @[Decoupled.scala 361:21]
  wire  q_721_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_721_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_721_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_721_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_721_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_721_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_722_clock; // @[Decoupled.scala 361:21]
  wire  q_722_reset; // @[Decoupled.scala 361:21]
  wire  q_722_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_722_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_722_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_722_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_722_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_722_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_723_clock; // @[Decoupled.scala 361:21]
  wire  q_723_reset; // @[Decoupled.scala 361:21]
  wire  q_723_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_723_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_723_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_723_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_723_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_723_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_724_clock; // @[Decoupled.scala 361:21]
  wire  q_724_reset; // @[Decoupled.scala 361:21]
  wire  q_724_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_724_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_724_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_724_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_724_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_724_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_725_clock; // @[Decoupled.scala 361:21]
  wire  q_725_reset; // @[Decoupled.scala 361:21]
  wire  q_725_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_725_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_725_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_725_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_725_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_725_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_726_clock; // @[Decoupled.scala 361:21]
  wire  q_726_reset; // @[Decoupled.scala 361:21]
  wire  q_726_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_726_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_726_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_726_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_726_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_726_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_727_clock; // @[Decoupled.scala 361:21]
  wire  q_727_reset; // @[Decoupled.scala 361:21]
  wire  q_727_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_727_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_727_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_727_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_727_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_727_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_728_clock; // @[Decoupled.scala 361:21]
  wire  q_728_reset; // @[Decoupled.scala 361:21]
  wire  q_728_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_728_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_728_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_728_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_728_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_728_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_729_clock; // @[Decoupled.scala 361:21]
  wire  q_729_reset; // @[Decoupled.scala 361:21]
  wire  q_729_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_729_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_729_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_729_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_729_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_729_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_730_clock; // @[Decoupled.scala 361:21]
  wire  q_730_reset; // @[Decoupled.scala 361:21]
  wire  q_730_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_730_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_730_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_730_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_730_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_730_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_731_clock; // @[Decoupled.scala 361:21]
  wire  q_731_reset; // @[Decoupled.scala 361:21]
  wire  q_731_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_731_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_731_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_731_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_731_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_731_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_732_clock; // @[Decoupled.scala 361:21]
  wire  q_732_reset; // @[Decoupled.scala 361:21]
  wire  q_732_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_732_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_732_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_732_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_732_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_732_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_733_clock; // @[Decoupled.scala 361:21]
  wire  q_733_reset; // @[Decoupled.scala 361:21]
  wire  q_733_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_733_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_733_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_733_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_733_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_733_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_734_clock; // @[Decoupled.scala 361:21]
  wire  q_734_reset; // @[Decoupled.scala 361:21]
  wire  q_734_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_734_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_734_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_734_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_734_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_734_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_735_clock; // @[Decoupled.scala 361:21]
  wire  q_735_reset; // @[Decoupled.scala 361:21]
  wire  q_735_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_735_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_735_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_735_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_735_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_735_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_736_clock; // @[Decoupled.scala 361:21]
  wire  q_736_reset; // @[Decoupled.scala 361:21]
  wire  q_736_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_736_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_736_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_736_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_736_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_736_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_737_clock; // @[Decoupled.scala 361:21]
  wire  q_737_reset; // @[Decoupled.scala 361:21]
  wire  q_737_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_737_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_737_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_737_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_737_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_737_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_738_clock; // @[Decoupled.scala 361:21]
  wire  q_738_reset; // @[Decoupled.scala 361:21]
  wire  q_738_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_738_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_738_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_738_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_738_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_738_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_739_clock; // @[Decoupled.scala 361:21]
  wire  q_739_reset; // @[Decoupled.scala 361:21]
  wire  q_739_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_739_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_739_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_739_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_739_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_739_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_740_clock; // @[Decoupled.scala 361:21]
  wire  q_740_reset; // @[Decoupled.scala 361:21]
  wire  q_740_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_740_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_740_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_740_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_740_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_740_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_741_clock; // @[Decoupled.scala 361:21]
  wire  q_741_reset; // @[Decoupled.scala 361:21]
  wire  q_741_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_741_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_741_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_741_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_741_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_741_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_742_clock; // @[Decoupled.scala 361:21]
  wire  q_742_reset; // @[Decoupled.scala 361:21]
  wire  q_742_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_742_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_742_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_742_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_742_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_742_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_743_clock; // @[Decoupled.scala 361:21]
  wire  q_743_reset; // @[Decoupled.scala 361:21]
  wire  q_743_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_743_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_743_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_743_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_743_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_743_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_744_clock; // @[Decoupled.scala 361:21]
  wire  q_744_reset; // @[Decoupled.scala 361:21]
  wire  q_744_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_744_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_744_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_744_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_744_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_744_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_745_clock; // @[Decoupled.scala 361:21]
  wire  q_745_reset; // @[Decoupled.scala 361:21]
  wire  q_745_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_745_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_745_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_745_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_745_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_745_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_746_clock; // @[Decoupled.scala 361:21]
  wire  q_746_reset; // @[Decoupled.scala 361:21]
  wire  q_746_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_746_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_746_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_746_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_746_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_746_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_747_clock; // @[Decoupled.scala 361:21]
  wire  q_747_reset; // @[Decoupled.scala 361:21]
  wire  q_747_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_747_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_747_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_747_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_747_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_747_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_748_clock; // @[Decoupled.scala 361:21]
  wire  q_748_reset; // @[Decoupled.scala 361:21]
  wire  q_748_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_748_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_748_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_748_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_748_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_748_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_749_clock; // @[Decoupled.scala 361:21]
  wire  q_749_reset; // @[Decoupled.scala 361:21]
  wire  q_749_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_749_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_749_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_749_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_749_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_749_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_750_clock; // @[Decoupled.scala 361:21]
  wire  q_750_reset; // @[Decoupled.scala 361:21]
  wire  q_750_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_750_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_750_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_750_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_750_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_750_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_751_clock; // @[Decoupled.scala 361:21]
  wire  q_751_reset; // @[Decoupled.scala 361:21]
  wire  q_751_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_751_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_751_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_751_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_751_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_751_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_752_clock; // @[Decoupled.scala 361:21]
  wire  q_752_reset; // @[Decoupled.scala 361:21]
  wire  q_752_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_752_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_752_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_752_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_752_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_752_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_753_clock; // @[Decoupled.scala 361:21]
  wire  q_753_reset; // @[Decoupled.scala 361:21]
  wire  q_753_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_753_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_753_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_753_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_753_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_753_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_754_clock; // @[Decoupled.scala 361:21]
  wire  q_754_reset; // @[Decoupled.scala 361:21]
  wire  q_754_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_754_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_754_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_754_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_754_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_754_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_755_clock; // @[Decoupled.scala 361:21]
  wire  q_755_reset; // @[Decoupled.scala 361:21]
  wire  q_755_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_755_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_755_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_755_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_755_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_755_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_756_clock; // @[Decoupled.scala 361:21]
  wire  q_756_reset; // @[Decoupled.scala 361:21]
  wire  q_756_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_756_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_756_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_756_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_756_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_756_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_757_clock; // @[Decoupled.scala 361:21]
  wire  q_757_reset; // @[Decoupled.scala 361:21]
  wire  q_757_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_757_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_757_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_757_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_757_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_757_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_758_clock; // @[Decoupled.scala 361:21]
  wire  q_758_reset; // @[Decoupled.scala 361:21]
  wire  q_758_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_758_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_758_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_758_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_758_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_758_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_759_clock; // @[Decoupled.scala 361:21]
  wire  q_759_reset; // @[Decoupled.scala 361:21]
  wire  q_759_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_759_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_759_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_759_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_759_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_759_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_760_clock; // @[Decoupled.scala 361:21]
  wire  q_760_reset; // @[Decoupled.scala 361:21]
  wire  q_760_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_760_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_760_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_760_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_760_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_760_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_761_clock; // @[Decoupled.scala 361:21]
  wire  q_761_reset; // @[Decoupled.scala 361:21]
  wire  q_761_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_761_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_761_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_761_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_761_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_761_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_762_clock; // @[Decoupled.scala 361:21]
  wire  q_762_reset; // @[Decoupled.scala 361:21]
  wire  q_762_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_762_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_762_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_762_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_762_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_762_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_763_clock; // @[Decoupled.scala 361:21]
  wire  q_763_reset; // @[Decoupled.scala 361:21]
  wire  q_763_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_763_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_763_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_763_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_763_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_763_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_764_clock; // @[Decoupled.scala 361:21]
  wire  q_764_reset; // @[Decoupled.scala 361:21]
  wire  q_764_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_764_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_764_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_764_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_764_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_764_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_765_clock; // @[Decoupled.scala 361:21]
  wire  q_765_reset; // @[Decoupled.scala 361:21]
  wire  q_765_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_765_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_765_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_765_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_765_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_765_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_766_clock; // @[Decoupled.scala 361:21]
  wire  q_766_reset; // @[Decoupled.scala 361:21]
  wire  q_766_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_766_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_766_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_766_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_766_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_766_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  q_767_clock; // @[Decoupled.scala 361:21]
  wire  q_767_reset; // @[Decoupled.scala 361:21]
  wire  q_767_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  q_767_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_767_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  q_767_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  q_767_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] q_767_io_deq_bits; // @[Decoupled.scala 361:21]
  ProcessingElement cols_0_0 ( // @[Stab.scala 85:60]
    .clock(cols_0_0_clock),
    .reset(cols_0_0_reset),
    .io_left_in_ready(cols_0_0_io_left_in_ready),
    .io_left_in_valid(cols_0_0_io_left_in_valid),
    .io_left_in_bits(cols_0_0_io_left_in_bits),
    .io_top_in_ready(cols_0_0_io_top_in_ready),
    .io_top_in_valid(cols_0_0_io_top_in_valid),
    .io_top_in_bits(cols_0_0_io_top_in_bits),
    .io_sum_ready(cols_0_0_io_sum_ready),
    .io_sum_valid(cols_0_0_io_sum_valid),
    .io_sum_bits(cols_0_0_io_sum_bits),
    .io_right_out_ready(cols_0_0_io_right_out_ready),
    .io_right_out_valid(cols_0_0_io_right_out_valid),
    .io_right_out_bits(cols_0_0_io_right_out_bits),
    .io_bottom_out_ready(cols_0_0_io_bottom_out_ready),
    .io_bottom_out_valid(cols_0_0_io_bottom_out_valid),
    .io_bottom_out_bits(cols_0_0_io_bottom_out_bits)
  );
  ProcessingElement cols_1_0 ( // @[Stab.scala 85:60]
    .clock(cols_1_0_clock),
    .reset(cols_1_0_reset),
    .io_left_in_ready(cols_1_0_io_left_in_ready),
    .io_left_in_valid(cols_1_0_io_left_in_valid),
    .io_left_in_bits(cols_1_0_io_left_in_bits),
    .io_top_in_ready(cols_1_0_io_top_in_ready),
    .io_top_in_valid(cols_1_0_io_top_in_valid),
    .io_top_in_bits(cols_1_0_io_top_in_bits),
    .io_sum_ready(cols_1_0_io_sum_ready),
    .io_sum_valid(cols_1_0_io_sum_valid),
    .io_sum_bits(cols_1_0_io_sum_bits),
    .io_right_out_ready(cols_1_0_io_right_out_ready),
    .io_right_out_valid(cols_1_0_io_right_out_valid),
    .io_right_out_bits(cols_1_0_io_right_out_bits),
    .io_bottom_out_ready(cols_1_0_io_bottom_out_ready),
    .io_bottom_out_valid(cols_1_0_io_bottom_out_valid),
    .io_bottom_out_bits(cols_1_0_io_bottom_out_bits)
  );
  ProcessingElement cols_2_0 ( // @[Stab.scala 85:60]
    .clock(cols_2_0_clock),
    .reset(cols_2_0_reset),
    .io_left_in_ready(cols_2_0_io_left_in_ready),
    .io_left_in_valid(cols_2_0_io_left_in_valid),
    .io_left_in_bits(cols_2_0_io_left_in_bits),
    .io_top_in_ready(cols_2_0_io_top_in_ready),
    .io_top_in_valid(cols_2_0_io_top_in_valid),
    .io_top_in_bits(cols_2_0_io_top_in_bits),
    .io_sum_ready(cols_2_0_io_sum_ready),
    .io_sum_valid(cols_2_0_io_sum_valid),
    .io_sum_bits(cols_2_0_io_sum_bits),
    .io_right_out_ready(cols_2_0_io_right_out_ready),
    .io_right_out_valid(cols_2_0_io_right_out_valid),
    .io_right_out_bits(cols_2_0_io_right_out_bits),
    .io_bottom_out_ready(cols_2_0_io_bottom_out_ready),
    .io_bottom_out_valid(cols_2_0_io_bottom_out_valid),
    .io_bottom_out_bits(cols_2_0_io_bottom_out_bits)
  );
  ProcessingElement cols_3_0 ( // @[Stab.scala 85:60]
    .clock(cols_3_0_clock),
    .reset(cols_3_0_reset),
    .io_left_in_ready(cols_3_0_io_left_in_ready),
    .io_left_in_valid(cols_3_0_io_left_in_valid),
    .io_left_in_bits(cols_3_0_io_left_in_bits),
    .io_top_in_ready(cols_3_0_io_top_in_ready),
    .io_top_in_valid(cols_3_0_io_top_in_valid),
    .io_top_in_bits(cols_3_0_io_top_in_bits),
    .io_sum_ready(cols_3_0_io_sum_ready),
    .io_sum_valid(cols_3_0_io_sum_valid),
    .io_sum_bits(cols_3_0_io_sum_bits),
    .io_right_out_ready(cols_3_0_io_right_out_ready),
    .io_right_out_valid(cols_3_0_io_right_out_valid),
    .io_right_out_bits(cols_3_0_io_right_out_bits),
    .io_bottom_out_ready(cols_3_0_io_bottom_out_ready),
    .io_bottom_out_valid(cols_3_0_io_bottom_out_valid),
    .io_bottom_out_bits(cols_3_0_io_bottom_out_bits)
  );
  ProcessingElement cols_4_0 ( // @[Stab.scala 85:60]
    .clock(cols_4_0_clock),
    .reset(cols_4_0_reset),
    .io_left_in_ready(cols_4_0_io_left_in_ready),
    .io_left_in_valid(cols_4_0_io_left_in_valid),
    .io_left_in_bits(cols_4_0_io_left_in_bits),
    .io_top_in_ready(cols_4_0_io_top_in_ready),
    .io_top_in_valid(cols_4_0_io_top_in_valid),
    .io_top_in_bits(cols_4_0_io_top_in_bits),
    .io_sum_ready(cols_4_0_io_sum_ready),
    .io_sum_valid(cols_4_0_io_sum_valid),
    .io_sum_bits(cols_4_0_io_sum_bits),
    .io_right_out_ready(cols_4_0_io_right_out_ready),
    .io_right_out_valid(cols_4_0_io_right_out_valid),
    .io_right_out_bits(cols_4_0_io_right_out_bits),
    .io_bottom_out_ready(cols_4_0_io_bottom_out_ready),
    .io_bottom_out_valid(cols_4_0_io_bottom_out_valid),
    .io_bottom_out_bits(cols_4_0_io_bottom_out_bits)
  );
  ProcessingElement cols_5_0 ( // @[Stab.scala 85:60]
    .clock(cols_5_0_clock),
    .reset(cols_5_0_reset),
    .io_left_in_ready(cols_5_0_io_left_in_ready),
    .io_left_in_valid(cols_5_0_io_left_in_valid),
    .io_left_in_bits(cols_5_0_io_left_in_bits),
    .io_top_in_ready(cols_5_0_io_top_in_ready),
    .io_top_in_valid(cols_5_0_io_top_in_valid),
    .io_top_in_bits(cols_5_0_io_top_in_bits),
    .io_sum_ready(cols_5_0_io_sum_ready),
    .io_sum_valid(cols_5_0_io_sum_valid),
    .io_sum_bits(cols_5_0_io_sum_bits),
    .io_right_out_ready(cols_5_0_io_right_out_ready),
    .io_right_out_valid(cols_5_0_io_right_out_valid),
    .io_right_out_bits(cols_5_0_io_right_out_bits),
    .io_bottom_out_ready(cols_5_0_io_bottom_out_ready),
    .io_bottom_out_valid(cols_5_0_io_bottom_out_valid),
    .io_bottom_out_bits(cols_5_0_io_bottom_out_bits)
  );
  ProcessingElement cols_6_0 ( // @[Stab.scala 85:60]
    .clock(cols_6_0_clock),
    .reset(cols_6_0_reset),
    .io_left_in_ready(cols_6_0_io_left_in_ready),
    .io_left_in_valid(cols_6_0_io_left_in_valid),
    .io_left_in_bits(cols_6_0_io_left_in_bits),
    .io_top_in_ready(cols_6_0_io_top_in_ready),
    .io_top_in_valid(cols_6_0_io_top_in_valid),
    .io_top_in_bits(cols_6_0_io_top_in_bits),
    .io_sum_ready(cols_6_0_io_sum_ready),
    .io_sum_valid(cols_6_0_io_sum_valid),
    .io_sum_bits(cols_6_0_io_sum_bits),
    .io_right_out_ready(cols_6_0_io_right_out_ready),
    .io_right_out_valid(cols_6_0_io_right_out_valid),
    .io_right_out_bits(cols_6_0_io_right_out_bits),
    .io_bottom_out_ready(cols_6_0_io_bottom_out_ready),
    .io_bottom_out_valid(cols_6_0_io_bottom_out_valid),
    .io_bottom_out_bits(cols_6_0_io_bottom_out_bits)
  );
  ProcessingElement cols_7_0 ( // @[Stab.scala 85:60]
    .clock(cols_7_0_clock),
    .reset(cols_7_0_reset),
    .io_left_in_ready(cols_7_0_io_left_in_ready),
    .io_left_in_valid(cols_7_0_io_left_in_valid),
    .io_left_in_bits(cols_7_0_io_left_in_bits),
    .io_top_in_ready(cols_7_0_io_top_in_ready),
    .io_top_in_valid(cols_7_0_io_top_in_valid),
    .io_top_in_bits(cols_7_0_io_top_in_bits),
    .io_sum_ready(cols_7_0_io_sum_ready),
    .io_sum_valid(cols_7_0_io_sum_valid),
    .io_sum_bits(cols_7_0_io_sum_bits),
    .io_right_out_ready(cols_7_0_io_right_out_ready),
    .io_right_out_valid(cols_7_0_io_right_out_valid),
    .io_right_out_bits(cols_7_0_io_right_out_bits),
    .io_bottom_out_ready(cols_7_0_io_bottom_out_ready),
    .io_bottom_out_valid(cols_7_0_io_bottom_out_valid),
    .io_bottom_out_bits(cols_7_0_io_bottom_out_bits)
  );
  ProcessingElement cols_8_0 ( // @[Stab.scala 85:60]
    .clock(cols_8_0_clock),
    .reset(cols_8_0_reset),
    .io_left_in_ready(cols_8_0_io_left_in_ready),
    .io_left_in_valid(cols_8_0_io_left_in_valid),
    .io_left_in_bits(cols_8_0_io_left_in_bits),
    .io_top_in_ready(cols_8_0_io_top_in_ready),
    .io_top_in_valid(cols_8_0_io_top_in_valid),
    .io_top_in_bits(cols_8_0_io_top_in_bits),
    .io_sum_ready(cols_8_0_io_sum_ready),
    .io_sum_valid(cols_8_0_io_sum_valid),
    .io_sum_bits(cols_8_0_io_sum_bits),
    .io_right_out_ready(cols_8_0_io_right_out_ready),
    .io_right_out_valid(cols_8_0_io_right_out_valid),
    .io_right_out_bits(cols_8_0_io_right_out_bits),
    .io_bottom_out_ready(cols_8_0_io_bottom_out_ready),
    .io_bottom_out_valid(cols_8_0_io_bottom_out_valid),
    .io_bottom_out_bits(cols_8_0_io_bottom_out_bits)
  );
  ProcessingElement cols_9_0 ( // @[Stab.scala 85:60]
    .clock(cols_9_0_clock),
    .reset(cols_9_0_reset),
    .io_left_in_ready(cols_9_0_io_left_in_ready),
    .io_left_in_valid(cols_9_0_io_left_in_valid),
    .io_left_in_bits(cols_9_0_io_left_in_bits),
    .io_top_in_ready(cols_9_0_io_top_in_ready),
    .io_top_in_valid(cols_9_0_io_top_in_valid),
    .io_top_in_bits(cols_9_0_io_top_in_bits),
    .io_sum_ready(cols_9_0_io_sum_ready),
    .io_sum_valid(cols_9_0_io_sum_valid),
    .io_sum_bits(cols_9_0_io_sum_bits),
    .io_right_out_ready(cols_9_0_io_right_out_ready),
    .io_right_out_valid(cols_9_0_io_right_out_valid),
    .io_right_out_bits(cols_9_0_io_right_out_bits),
    .io_bottom_out_ready(cols_9_0_io_bottom_out_ready),
    .io_bottom_out_valid(cols_9_0_io_bottom_out_valid),
    .io_bottom_out_bits(cols_9_0_io_bottom_out_bits)
  );
  ProcessingElement cols_10_0 ( // @[Stab.scala 85:60]
    .clock(cols_10_0_clock),
    .reset(cols_10_0_reset),
    .io_left_in_ready(cols_10_0_io_left_in_ready),
    .io_left_in_valid(cols_10_0_io_left_in_valid),
    .io_left_in_bits(cols_10_0_io_left_in_bits),
    .io_top_in_ready(cols_10_0_io_top_in_ready),
    .io_top_in_valid(cols_10_0_io_top_in_valid),
    .io_top_in_bits(cols_10_0_io_top_in_bits),
    .io_sum_ready(cols_10_0_io_sum_ready),
    .io_sum_valid(cols_10_0_io_sum_valid),
    .io_sum_bits(cols_10_0_io_sum_bits),
    .io_right_out_ready(cols_10_0_io_right_out_ready),
    .io_right_out_valid(cols_10_0_io_right_out_valid),
    .io_right_out_bits(cols_10_0_io_right_out_bits),
    .io_bottom_out_ready(cols_10_0_io_bottom_out_ready),
    .io_bottom_out_valid(cols_10_0_io_bottom_out_valid),
    .io_bottom_out_bits(cols_10_0_io_bottom_out_bits)
  );
  ProcessingElement cols_11_0 ( // @[Stab.scala 85:60]
    .clock(cols_11_0_clock),
    .reset(cols_11_0_reset),
    .io_left_in_ready(cols_11_0_io_left_in_ready),
    .io_left_in_valid(cols_11_0_io_left_in_valid),
    .io_left_in_bits(cols_11_0_io_left_in_bits),
    .io_top_in_ready(cols_11_0_io_top_in_ready),
    .io_top_in_valid(cols_11_0_io_top_in_valid),
    .io_top_in_bits(cols_11_0_io_top_in_bits),
    .io_sum_ready(cols_11_0_io_sum_ready),
    .io_sum_valid(cols_11_0_io_sum_valid),
    .io_sum_bits(cols_11_0_io_sum_bits),
    .io_right_out_ready(cols_11_0_io_right_out_ready),
    .io_right_out_valid(cols_11_0_io_right_out_valid),
    .io_right_out_bits(cols_11_0_io_right_out_bits),
    .io_bottom_out_ready(cols_11_0_io_bottom_out_ready),
    .io_bottom_out_valid(cols_11_0_io_bottom_out_valid),
    .io_bottom_out_bits(cols_11_0_io_bottom_out_bits)
  );
  ProcessingElement cols_12_0 ( // @[Stab.scala 85:60]
    .clock(cols_12_0_clock),
    .reset(cols_12_0_reset),
    .io_left_in_ready(cols_12_0_io_left_in_ready),
    .io_left_in_valid(cols_12_0_io_left_in_valid),
    .io_left_in_bits(cols_12_0_io_left_in_bits),
    .io_top_in_ready(cols_12_0_io_top_in_ready),
    .io_top_in_valid(cols_12_0_io_top_in_valid),
    .io_top_in_bits(cols_12_0_io_top_in_bits),
    .io_sum_ready(cols_12_0_io_sum_ready),
    .io_sum_valid(cols_12_0_io_sum_valid),
    .io_sum_bits(cols_12_0_io_sum_bits),
    .io_right_out_ready(cols_12_0_io_right_out_ready),
    .io_right_out_valid(cols_12_0_io_right_out_valid),
    .io_right_out_bits(cols_12_0_io_right_out_bits),
    .io_bottom_out_ready(cols_12_0_io_bottom_out_ready),
    .io_bottom_out_valid(cols_12_0_io_bottom_out_valid),
    .io_bottom_out_bits(cols_12_0_io_bottom_out_bits)
  );
  ProcessingElement cols_13_0 ( // @[Stab.scala 85:60]
    .clock(cols_13_0_clock),
    .reset(cols_13_0_reset),
    .io_left_in_ready(cols_13_0_io_left_in_ready),
    .io_left_in_valid(cols_13_0_io_left_in_valid),
    .io_left_in_bits(cols_13_0_io_left_in_bits),
    .io_top_in_ready(cols_13_0_io_top_in_ready),
    .io_top_in_valid(cols_13_0_io_top_in_valid),
    .io_top_in_bits(cols_13_0_io_top_in_bits),
    .io_sum_ready(cols_13_0_io_sum_ready),
    .io_sum_valid(cols_13_0_io_sum_valid),
    .io_sum_bits(cols_13_0_io_sum_bits),
    .io_right_out_ready(cols_13_0_io_right_out_ready),
    .io_right_out_valid(cols_13_0_io_right_out_valid),
    .io_right_out_bits(cols_13_0_io_right_out_bits),
    .io_bottom_out_ready(cols_13_0_io_bottom_out_ready),
    .io_bottom_out_valid(cols_13_0_io_bottom_out_valid),
    .io_bottom_out_bits(cols_13_0_io_bottom_out_bits)
  );
  ProcessingElement cols_14_0 ( // @[Stab.scala 85:60]
    .clock(cols_14_0_clock),
    .reset(cols_14_0_reset),
    .io_left_in_ready(cols_14_0_io_left_in_ready),
    .io_left_in_valid(cols_14_0_io_left_in_valid),
    .io_left_in_bits(cols_14_0_io_left_in_bits),
    .io_top_in_ready(cols_14_0_io_top_in_ready),
    .io_top_in_valid(cols_14_0_io_top_in_valid),
    .io_top_in_bits(cols_14_0_io_top_in_bits),
    .io_sum_ready(cols_14_0_io_sum_ready),
    .io_sum_valid(cols_14_0_io_sum_valid),
    .io_sum_bits(cols_14_0_io_sum_bits),
    .io_right_out_ready(cols_14_0_io_right_out_ready),
    .io_right_out_valid(cols_14_0_io_right_out_valid),
    .io_right_out_bits(cols_14_0_io_right_out_bits),
    .io_bottom_out_ready(cols_14_0_io_bottom_out_ready),
    .io_bottom_out_valid(cols_14_0_io_bottom_out_valid),
    .io_bottom_out_bits(cols_14_0_io_bottom_out_bits)
  );
  ProcessingElement cols_15_0 ( // @[Stab.scala 85:60]
    .clock(cols_15_0_clock),
    .reset(cols_15_0_reset),
    .io_left_in_ready(cols_15_0_io_left_in_ready),
    .io_left_in_valid(cols_15_0_io_left_in_valid),
    .io_left_in_bits(cols_15_0_io_left_in_bits),
    .io_top_in_ready(cols_15_0_io_top_in_ready),
    .io_top_in_valid(cols_15_0_io_top_in_valid),
    .io_top_in_bits(cols_15_0_io_top_in_bits),
    .io_sum_ready(cols_15_0_io_sum_ready),
    .io_sum_valid(cols_15_0_io_sum_valid),
    .io_sum_bits(cols_15_0_io_sum_bits),
    .io_right_out_ready(cols_15_0_io_right_out_ready),
    .io_right_out_valid(cols_15_0_io_right_out_valid),
    .io_right_out_bits(cols_15_0_io_right_out_bits),
    .io_bottom_out_ready(cols_15_0_io_bottom_out_ready),
    .io_bottom_out_valid(cols_15_0_io_bottom_out_valid),
    .io_bottom_out_bits(cols_15_0_io_bottom_out_bits)
  );
  ProcessingElement cols_0_1 ( // @[Stab.scala 85:60]
    .clock(cols_0_1_clock),
    .reset(cols_0_1_reset),
    .io_left_in_ready(cols_0_1_io_left_in_ready),
    .io_left_in_valid(cols_0_1_io_left_in_valid),
    .io_left_in_bits(cols_0_1_io_left_in_bits),
    .io_top_in_ready(cols_0_1_io_top_in_ready),
    .io_top_in_valid(cols_0_1_io_top_in_valid),
    .io_top_in_bits(cols_0_1_io_top_in_bits),
    .io_sum_ready(cols_0_1_io_sum_ready),
    .io_sum_valid(cols_0_1_io_sum_valid),
    .io_sum_bits(cols_0_1_io_sum_bits),
    .io_right_out_ready(cols_0_1_io_right_out_ready),
    .io_right_out_valid(cols_0_1_io_right_out_valid),
    .io_right_out_bits(cols_0_1_io_right_out_bits),
    .io_bottom_out_ready(cols_0_1_io_bottom_out_ready),
    .io_bottom_out_valid(cols_0_1_io_bottom_out_valid),
    .io_bottom_out_bits(cols_0_1_io_bottom_out_bits)
  );
  ProcessingElement cols_1_1 ( // @[Stab.scala 85:60]
    .clock(cols_1_1_clock),
    .reset(cols_1_1_reset),
    .io_left_in_ready(cols_1_1_io_left_in_ready),
    .io_left_in_valid(cols_1_1_io_left_in_valid),
    .io_left_in_bits(cols_1_1_io_left_in_bits),
    .io_top_in_ready(cols_1_1_io_top_in_ready),
    .io_top_in_valid(cols_1_1_io_top_in_valid),
    .io_top_in_bits(cols_1_1_io_top_in_bits),
    .io_sum_ready(cols_1_1_io_sum_ready),
    .io_sum_valid(cols_1_1_io_sum_valid),
    .io_sum_bits(cols_1_1_io_sum_bits),
    .io_right_out_ready(cols_1_1_io_right_out_ready),
    .io_right_out_valid(cols_1_1_io_right_out_valid),
    .io_right_out_bits(cols_1_1_io_right_out_bits),
    .io_bottom_out_ready(cols_1_1_io_bottom_out_ready),
    .io_bottom_out_valid(cols_1_1_io_bottom_out_valid),
    .io_bottom_out_bits(cols_1_1_io_bottom_out_bits)
  );
  ProcessingElement cols_2_1 ( // @[Stab.scala 85:60]
    .clock(cols_2_1_clock),
    .reset(cols_2_1_reset),
    .io_left_in_ready(cols_2_1_io_left_in_ready),
    .io_left_in_valid(cols_2_1_io_left_in_valid),
    .io_left_in_bits(cols_2_1_io_left_in_bits),
    .io_top_in_ready(cols_2_1_io_top_in_ready),
    .io_top_in_valid(cols_2_1_io_top_in_valid),
    .io_top_in_bits(cols_2_1_io_top_in_bits),
    .io_sum_ready(cols_2_1_io_sum_ready),
    .io_sum_valid(cols_2_1_io_sum_valid),
    .io_sum_bits(cols_2_1_io_sum_bits),
    .io_right_out_ready(cols_2_1_io_right_out_ready),
    .io_right_out_valid(cols_2_1_io_right_out_valid),
    .io_right_out_bits(cols_2_1_io_right_out_bits),
    .io_bottom_out_ready(cols_2_1_io_bottom_out_ready),
    .io_bottom_out_valid(cols_2_1_io_bottom_out_valid),
    .io_bottom_out_bits(cols_2_1_io_bottom_out_bits)
  );
  ProcessingElement cols_3_1 ( // @[Stab.scala 85:60]
    .clock(cols_3_1_clock),
    .reset(cols_3_1_reset),
    .io_left_in_ready(cols_3_1_io_left_in_ready),
    .io_left_in_valid(cols_3_1_io_left_in_valid),
    .io_left_in_bits(cols_3_1_io_left_in_bits),
    .io_top_in_ready(cols_3_1_io_top_in_ready),
    .io_top_in_valid(cols_3_1_io_top_in_valid),
    .io_top_in_bits(cols_3_1_io_top_in_bits),
    .io_sum_ready(cols_3_1_io_sum_ready),
    .io_sum_valid(cols_3_1_io_sum_valid),
    .io_sum_bits(cols_3_1_io_sum_bits),
    .io_right_out_ready(cols_3_1_io_right_out_ready),
    .io_right_out_valid(cols_3_1_io_right_out_valid),
    .io_right_out_bits(cols_3_1_io_right_out_bits),
    .io_bottom_out_ready(cols_3_1_io_bottom_out_ready),
    .io_bottom_out_valid(cols_3_1_io_bottom_out_valid),
    .io_bottom_out_bits(cols_3_1_io_bottom_out_bits)
  );
  ProcessingElement cols_4_1 ( // @[Stab.scala 85:60]
    .clock(cols_4_1_clock),
    .reset(cols_4_1_reset),
    .io_left_in_ready(cols_4_1_io_left_in_ready),
    .io_left_in_valid(cols_4_1_io_left_in_valid),
    .io_left_in_bits(cols_4_1_io_left_in_bits),
    .io_top_in_ready(cols_4_1_io_top_in_ready),
    .io_top_in_valid(cols_4_1_io_top_in_valid),
    .io_top_in_bits(cols_4_1_io_top_in_bits),
    .io_sum_ready(cols_4_1_io_sum_ready),
    .io_sum_valid(cols_4_1_io_sum_valid),
    .io_sum_bits(cols_4_1_io_sum_bits),
    .io_right_out_ready(cols_4_1_io_right_out_ready),
    .io_right_out_valid(cols_4_1_io_right_out_valid),
    .io_right_out_bits(cols_4_1_io_right_out_bits),
    .io_bottom_out_ready(cols_4_1_io_bottom_out_ready),
    .io_bottom_out_valid(cols_4_1_io_bottom_out_valid),
    .io_bottom_out_bits(cols_4_1_io_bottom_out_bits)
  );
  ProcessingElement cols_5_1 ( // @[Stab.scala 85:60]
    .clock(cols_5_1_clock),
    .reset(cols_5_1_reset),
    .io_left_in_ready(cols_5_1_io_left_in_ready),
    .io_left_in_valid(cols_5_1_io_left_in_valid),
    .io_left_in_bits(cols_5_1_io_left_in_bits),
    .io_top_in_ready(cols_5_1_io_top_in_ready),
    .io_top_in_valid(cols_5_1_io_top_in_valid),
    .io_top_in_bits(cols_5_1_io_top_in_bits),
    .io_sum_ready(cols_5_1_io_sum_ready),
    .io_sum_valid(cols_5_1_io_sum_valid),
    .io_sum_bits(cols_5_1_io_sum_bits),
    .io_right_out_ready(cols_5_1_io_right_out_ready),
    .io_right_out_valid(cols_5_1_io_right_out_valid),
    .io_right_out_bits(cols_5_1_io_right_out_bits),
    .io_bottom_out_ready(cols_5_1_io_bottom_out_ready),
    .io_bottom_out_valid(cols_5_1_io_bottom_out_valid),
    .io_bottom_out_bits(cols_5_1_io_bottom_out_bits)
  );
  ProcessingElement cols_6_1 ( // @[Stab.scala 85:60]
    .clock(cols_6_1_clock),
    .reset(cols_6_1_reset),
    .io_left_in_ready(cols_6_1_io_left_in_ready),
    .io_left_in_valid(cols_6_1_io_left_in_valid),
    .io_left_in_bits(cols_6_1_io_left_in_bits),
    .io_top_in_ready(cols_6_1_io_top_in_ready),
    .io_top_in_valid(cols_6_1_io_top_in_valid),
    .io_top_in_bits(cols_6_1_io_top_in_bits),
    .io_sum_ready(cols_6_1_io_sum_ready),
    .io_sum_valid(cols_6_1_io_sum_valid),
    .io_sum_bits(cols_6_1_io_sum_bits),
    .io_right_out_ready(cols_6_1_io_right_out_ready),
    .io_right_out_valid(cols_6_1_io_right_out_valid),
    .io_right_out_bits(cols_6_1_io_right_out_bits),
    .io_bottom_out_ready(cols_6_1_io_bottom_out_ready),
    .io_bottom_out_valid(cols_6_1_io_bottom_out_valid),
    .io_bottom_out_bits(cols_6_1_io_bottom_out_bits)
  );
  ProcessingElement cols_7_1 ( // @[Stab.scala 85:60]
    .clock(cols_7_1_clock),
    .reset(cols_7_1_reset),
    .io_left_in_ready(cols_7_1_io_left_in_ready),
    .io_left_in_valid(cols_7_1_io_left_in_valid),
    .io_left_in_bits(cols_7_1_io_left_in_bits),
    .io_top_in_ready(cols_7_1_io_top_in_ready),
    .io_top_in_valid(cols_7_1_io_top_in_valid),
    .io_top_in_bits(cols_7_1_io_top_in_bits),
    .io_sum_ready(cols_7_1_io_sum_ready),
    .io_sum_valid(cols_7_1_io_sum_valid),
    .io_sum_bits(cols_7_1_io_sum_bits),
    .io_right_out_ready(cols_7_1_io_right_out_ready),
    .io_right_out_valid(cols_7_1_io_right_out_valid),
    .io_right_out_bits(cols_7_1_io_right_out_bits),
    .io_bottom_out_ready(cols_7_1_io_bottom_out_ready),
    .io_bottom_out_valid(cols_7_1_io_bottom_out_valid),
    .io_bottom_out_bits(cols_7_1_io_bottom_out_bits)
  );
  ProcessingElement cols_8_1 ( // @[Stab.scala 85:60]
    .clock(cols_8_1_clock),
    .reset(cols_8_1_reset),
    .io_left_in_ready(cols_8_1_io_left_in_ready),
    .io_left_in_valid(cols_8_1_io_left_in_valid),
    .io_left_in_bits(cols_8_1_io_left_in_bits),
    .io_top_in_ready(cols_8_1_io_top_in_ready),
    .io_top_in_valid(cols_8_1_io_top_in_valid),
    .io_top_in_bits(cols_8_1_io_top_in_bits),
    .io_sum_ready(cols_8_1_io_sum_ready),
    .io_sum_valid(cols_8_1_io_sum_valid),
    .io_sum_bits(cols_8_1_io_sum_bits),
    .io_right_out_ready(cols_8_1_io_right_out_ready),
    .io_right_out_valid(cols_8_1_io_right_out_valid),
    .io_right_out_bits(cols_8_1_io_right_out_bits),
    .io_bottom_out_ready(cols_8_1_io_bottom_out_ready),
    .io_bottom_out_valid(cols_8_1_io_bottom_out_valid),
    .io_bottom_out_bits(cols_8_1_io_bottom_out_bits)
  );
  ProcessingElement cols_9_1 ( // @[Stab.scala 85:60]
    .clock(cols_9_1_clock),
    .reset(cols_9_1_reset),
    .io_left_in_ready(cols_9_1_io_left_in_ready),
    .io_left_in_valid(cols_9_1_io_left_in_valid),
    .io_left_in_bits(cols_9_1_io_left_in_bits),
    .io_top_in_ready(cols_9_1_io_top_in_ready),
    .io_top_in_valid(cols_9_1_io_top_in_valid),
    .io_top_in_bits(cols_9_1_io_top_in_bits),
    .io_sum_ready(cols_9_1_io_sum_ready),
    .io_sum_valid(cols_9_1_io_sum_valid),
    .io_sum_bits(cols_9_1_io_sum_bits),
    .io_right_out_ready(cols_9_1_io_right_out_ready),
    .io_right_out_valid(cols_9_1_io_right_out_valid),
    .io_right_out_bits(cols_9_1_io_right_out_bits),
    .io_bottom_out_ready(cols_9_1_io_bottom_out_ready),
    .io_bottom_out_valid(cols_9_1_io_bottom_out_valid),
    .io_bottom_out_bits(cols_9_1_io_bottom_out_bits)
  );
  ProcessingElement cols_10_1 ( // @[Stab.scala 85:60]
    .clock(cols_10_1_clock),
    .reset(cols_10_1_reset),
    .io_left_in_ready(cols_10_1_io_left_in_ready),
    .io_left_in_valid(cols_10_1_io_left_in_valid),
    .io_left_in_bits(cols_10_1_io_left_in_bits),
    .io_top_in_ready(cols_10_1_io_top_in_ready),
    .io_top_in_valid(cols_10_1_io_top_in_valid),
    .io_top_in_bits(cols_10_1_io_top_in_bits),
    .io_sum_ready(cols_10_1_io_sum_ready),
    .io_sum_valid(cols_10_1_io_sum_valid),
    .io_sum_bits(cols_10_1_io_sum_bits),
    .io_right_out_ready(cols_10_1_io_right_out_ready),
    .io_right_out_valid(cols_10_1_io_right_out_valid),
    .io_right_out_bits(cols_10_1_io_right_out_bits),
    .io_bottom_out_ready(cols_10_1_io_bottom_out_ready),
    .io_bottom_out_valid(cols_10_1_io_bottom_out_valid),
    .io_bottom_out_bits(cols_10_1_io_bottom_out_bits)
  );
  ProcessingElement cols_11_1 ( // @[Stab.scala 85:60]
    .clock(cols_11_1_clock),
    .reset(cols_11_1_reset),
    .io_left_in_ready(cols_11_1_io_left_in_ready),
    .io_left_in_valid(cols_11_1_io_left_in_valid),
    .io_left_in_bits(cols_11_1_io_left_in_bits),
    .io_top_in_ready(cols_11_1_io_top_in_ready),
    .io_top_in_valid(cols_11_1_io_top_in_valid),
    .io_top_in_bits(cols_11_1_io_top_in_bits),
    .io_sum_ready(cols_11_1_io_sum_ready),
    .io_sum_valid(cols_11_1_io_sum_valid),
    .io_sum_bits(cols_11_1_io_sum_bits),
    .io_right_out_ready(cols_11_1_io_right_out_ready),
    .io_right_out_valid(cols_11_1_io_right_out_valid),
    .io_right_out_bits(cols_11_1_io_right_out_bits),
    .io_bottom_out_ready(cols_11_1_io_bottom_out_ready),
    .io_bottom_out_valid(cols_11_1_io_bottom_out_valid),
    .io_bottom_out_bits(cols_11_1_io_bottom_out_bits)
  );
  ProcessingElement cols_12_1 ( // @[Stab.scala 85:60]
    .clock(cols_12_1_clock),
    .reset(cols_12_1_reset),
    .io_left_in_ready(cols_12_1_io_left_in_ready),
    .io_left_in_valid(cols_12_1_io_left_in_valid),
    .io_left_in_bits(cols_12_1_io_left_in_bits),
    .io_top_in_ready(cols_12_1_io_top_in_ready),
    .io_top_in_valid(cols_12_1_io_top_in_valid),
    .io_top_in_bits(cols_12_1_io_top_in_bits),
    .io_sum_ready(cols_12_1_io_sum_ready),
    .io_sum_valid(cols_12_1_io_sum_valid),
    .io_sum_bits(cols_12_1_io_sum_bits),
    .io_right_out_ready(cols_12_1_io_right_out_ready),
    .io_right_out_valid(cols_12_1_io_right_out_valid),
    .io_right_out_bits(cols_12_1_io_right_out_bits),
    .io_bottom_out_ready(cols_12_1_io_bottom_out_ready),
    .io_bottom_out_valid(cols_12_1_io_bottom_out_valid),
    .io_bottom_out_bits(cols_12_1_io_bottom_out_bits)
  );
  ProcessingElement cols_13_1 ( // @[Stab.scala 85:60]
    .clock(cols_13_1_clock),
    .reset(cols_13_1_reset),
    .io_left_in_ready(cols_13_1_io_left_in_ready),
    .io_left_in_valid(cols_13_1_io_left_in_valid),
    .io_left_in_bits(cols_13_1_io_left_in_bits),
    .io_top_in_ready(cols_13_1_io_top_in_ready),
    .io_top_in_valid(cols_13_1_io_top_in_valid),
    .io_top_in_bits(cols_13_1_io_top_in_bits),
    .io_sum_ready(cols_13_1_io_sum_ready),
    .io_sum_valid(cols_13_1_io_sum_valid),
    .io_sum_bits(cols_13_1_io_sum_bits),
    .io_right_out_ready(cols_13_1_io_right_out_ready),
    .io_right_out_valid(cols_13_1_io_right_out_valid),
    .io_right_out_bits(cols_13_1_io_right_out_bits),
    .io_bottom_out_ready(cols_13_1_io_bottom_out_ready),
    .io_bottom_out_valid(cols_13_1_io_bottom_out_valid),
    .io_bottom_out_bits(cols_13_1_io_bottom_out_bits)
  );
  ProcessingElement cols_14_1 ( // @[Stab.scala 85:60]
    .clock(cols_14_1_clock),
    .reset(cols_14_1_reset),
    .io_left_in_ready(cols_14_1_io_left_in_ready),
    .io_left_in_valid(cols_14_1_io_left_in_valid),
    .io_left_in_bits(cols_14_1_io_left_in_bits),
    .io_top_in_ready(cols_14_1_io_top_in_ready),
    .io_top_in_valid(cols_14_1_io_top_in_valid),
    .io_top_in_bits(cols_14_1_io_top_in_bits),
    .io_sum_ready(cols_14_1_io_sum_ready),
    .io_sum_valid(cols_14_1_io_sum_valid),
    .io_sum_bits(cols_14_1_io_sum_bits),
    .io_right_out_ready(cols_14_1_io_right_out_ready),
    .io_right_out_valid(cols_14_1_io_right_out_valid),
    .io_right_out_bits(cols_14_1_io_right_out_bits),
    .io_bottom_out_ready(cols_14_1_io_bottom_out_ready),
    .io_bottom_out_valid(cols_14_1_io_bottom_out_valid),
    .io_bottom_out_bits(cols_14_1_io_bottom_out_bits)
  );
  ProcessingElement cols_15_1 ( // @[Stab.scala 85:60]
    .clock(cols_15_1_clock),
    .reset(cols_15_1_reset),
    .io_left_in_ready(cols_15_1_io_left_in_ready),
    .io_left_in_valid(cols_15_1_io_left_in_valid),
    .io_left_in_bits(cols_15_1_io_left_in_bits),
    .io_top_in_ready(cols_15_1_io_top_in_ready),
    .io_top_in_valid(cols_15_1_io_top_in_valid),
    .io_top_in_bits(cols_15_1_io_top_in_bits),
    .io_sum_ready(cols_15_1_io_sum_ready),
    .io_sum_valid(cols_15_1_io_sum_valid),
    .io_sum_bits(cols_15_1_io_sum_bits),
    .io_right_out_ready(cols_15_1_io_right_out_ready),
    .io_right_out_valid(cols_15_1_io_right_out_valid),
    .io_right_out_bits(cols_15_1_io_right_out_bits),
    .io_bottom_out_ready(cols_15_1_io_bottom_out_ready),
    .io_bottom_out_valid(cols_15_1_io_bottom_out_valid),
    .io_bottom_out_bits(cols_15_1_io_bottom_out_bits)
  );
  ProcessingElement cols_0_2 ( // @[Stab.scala 85:60]
    .clock(cols_0_2_clock),
    .reset(cols_0_2_reset),
    .io_left_in_ready(cols_0_2_io_left_in_ready),
    .io_left_in_valid(cols_0_2_io_left_in_valid),
    .io_left_in_bits(cols_0_2_io_left_in_bits),
    .io_top_in_ready(cols_0_2_io_top_in_ready),
    .io_top_in_valid(cols_0_2_io_top_in_valid),
    .io_top_in_bits(cols_0_2_io_top_in_bits),
    .io_sum_ready(cols_0_2_io_sum_ready),
    .io_sum_valid(cols_0_2_io_sum_valid),
    .io_sum_bits(cols_0_2_io_sum_bits),
    .io_right_out_ready(cols_0_2_io_right_out_ready),
    .io_right_out_valid(cols_0_2_io_right_out_valid),
    .io_right_out_bits(cols_0_2_io_right_out_bits),
    .io_bottom_out_ready(cols_0_2_io_bottom_out_ready),
    .io_bottom_out_valid(cols_0_2_io_bottom_out_valid),
    .io_bottom_out_bits(cols_0_2_io_bottom_out_bits)
  );
  ProcessingElement cols_1_2 ( // @[Stab.scala 85:60]
    .clock(cols_1_2_clock),
    .reset(cols_1_2_reset),
    .io_left_in_ready(cols_1_2_io_left_in_ready),
    .io_left_in_valid(cols_1_2_io_left_in_valid),
    .io_left_in_bits(cols_1_2_io_left_in_bits),
    .io_top_in_ready(cols_1_2_io_top_in_ready),
    .io_top_in_valid(cols_1_2_io_top_in_valid),
    .io_top_in_bits(cols_1_2_io_top_in_bits),
    .io_sum_ready(cols_1_2_io_sum_ready),
    .io_sum_valid(cols_1_2_io_sum_valid),
    .io_sum_bits(cols_1_2_io_sum_bits),
    .io_right_out_ready(cols_1_2_io_right_out_ready),
    .io_right_out_valid(cols_1_2_io_right_out_valid),
    .io_right_out_bits(cols_1_2_io_right_out_bits),
    .io_bottom_out_ready(cols_1_2_io_bottom_out_ready),
    .io_bottom_out_valid(cols_1_2_io_bottom_out_valid),
    .io_bottom_out_bits(cols_1_2_io_bottom_out_bits)
  );
  ProcessingElement cols_2_2 ( // @[Stab.scala 85:60]
    .clock(cols_2_2_clock),
    .reset(cols_2_2_reset),
    .io_left_in_ready(cols_2_2_io_left_in_ready),
    .io_left_in_valid(cols_2_2_io_left_in_valid),
    .io_left_in_bits(cols_2_2_io_left_in_bits),
    .io_top_in_ready(cols_2_2_io_top_in_ready),
    .io_top_in_valid(cols_2_2_io_top_in_valid),
    .io_top_in_bits(cols_2_2_io_top_in_bits),
    .io_sum_ready(cols_2_2_io_sum_ready),
    .io_sum_valid(cols_2_2_io_sum_valid),
    .io_sum_bits(cols_2_2_io_sum_bits),
    .io_right_out_ready(cols_2_2_io_right_out_ready),
    .io_right_out_valid(cols_2_2_io_right_out_valid),
    .io_right_out_bits(cols_2_2_io_right_out_bits),
    .io_bottom_out_ready(cols_2_2_io_bottom_out_ready),
    .io_bottom_out_valid(cols_2_2_io_bottom_out_valid),
    .io_bottom_out_bits(cols_2_2_io_bottom_out_bits)
  );
  ProcessingElement cols_3_2 ( // @[Stab.scala 85:60]
    .clock(cols_3_2_clock),
    .reset(cols_3_2_reset),
    .io_left_in_ready(cols_3_2_io_left_in_ready),
    .io_left_in_valid(cols_3_2_io_left_in_valid),
    .io_left_in_bits(cols_3_2_io_left_in_bits),
    .io_top_in_ready(cols_3_2_io_top_in_ready),
    .io_top_in_valid(cols_3_2_io_top_in_valid),
    .io_top_in_bits(cols_3_2_io_top_in_bits),
    .io_sum_ready(cols_3_2_io_sum_ready),
    .io_sum_valid(cols_3_2_io_sum_valid),
    .io_sum_bits(cols_3_2_io_sum_bits),
    .io_right_out_ready(cols_3_2_io_right_out_ready),
    .io_right_out_valid(cols_3_2_io_right_out_valid),
    .io_right_out_bits(cols_3_2_io_right_out_bits),
    .io_bottom_out_ready(cols_3_2_io_bottom_out_ready),
    .io_bottom_out_valid(cols_3_2_io_bottom_out_valid),
    .io_bottom_out_bits(cols_3_2_io_bottom_out_bits)
  );
  ProcessingElement cols_4_2 ( // @[Stab.scala 85:60]
    .clock(cols_4_2_clock),
    .reset(cols_4_2_reset),
    .io_left_in_ready(cols_4_2_io_left_in_ready),
    .io_left_in_valid(cols_4_2_io_left_in_valid),
    .io_left_in_bits(cols_4_2_io_left_in_bits),
    .io_top_in_ready(cols_4_2_io_top_in_ready),
    .io_top_in_valid(cols_4_2_io_top_in_valid),
    .io_top_in_bits(cols_4_2_io_top_in_bits),
    .io_sum_ready(cols_4_2_io_sum_ready),
    .io_sum_valid(cols_4_2_io_sum_valid),
    .io_sum_bits(cols_4_2_io_sum_bits),
    .io_right_out_ready(cols_4_2_io_right_out_ready),
    .io_right_out_valid(cols_4_2_io_right_out_valid),
    .io_right_out_bits(cols_4_2_io_right_out_bits),
    .io_bottom_out_ready(cols_4_2_io_bottom_out_ready),
    .io_bottom_out_valid(cols_4_2_io_bottom_out_valid),
    .io_bottom_out_bits(cols_4_2_io_bottom_out_bits)
  );
  ProcessingElement cols_5_2 ( // @[Stab.scala 85:60]
    .clock(cols_5_2_clock),
    .reset(cols_5_2_reset),
    .io_left_in_ready(cols_5_2_io_left_in_ready),
    .io_left_in_valid(cols_5_2_io_left_in_valid),
    .io_left_in_bits(cols_5_2_io_left_in_bits),
    .io_top_in_ready(cols_5_2_io_top_in_ready),
    .io_top_in_valid(cols_5_2_io_top_in_valid),
    .io_top_in_bits(cols_5_2_io_top_in_bits),
    .io_sum_ready(cols_5_2_io_sum_ready),
    .io_sum_valid(cols_5_2_io_sum_valid),
    .io_sum_bits(cols_5_2_io_sum_bits),
    .io_right_out_ready(cols_5_2_io_right_out_ready),
    .io_right_out_valid(cols_5_2_io_right_out_valid),
    .io_right_out_bits(cols_5_2_io_right_out_bits),
    .io_bottom_out_ready(cols_5_2_io_bottom_out_ready),
    .io_bottom_out_valid(cols_5_2_io_bottom_out_valid),
    .io_bottom_out_bits(cols_5_2_io_bottom_out_bits)
  );
  ProcessingElement cols_6_2 ( // @[Stab.scala 85:60]
    .clock(cols_6_2_clock),
    .reset(cols_6_2_reset),
    .io_left_in_ready(cols_6_2_io_left_in_ready),
    .io_left_in_valid(cols_6_2_io_left_in_valid),
    .io_left_in_bits(cols_6_2_io_left_in_bits),
    .io_top_in_ready(cols_6_2_io_top_in_ready),
    .io_top_in_valid(cols_6_2_io_top_in_valid),
    .io_top_in_bits(cols_6_2_io_top_in_bits),
    .io_sum_ready(cols_6_2_io_sum_ready),
    .io_sum_valid(cols_6_2_io_sum_valid),
    .io_sum_bits(cols_6_2_io_sum_bits),
    .io_right_out_ready(cols_6_2_io_right_out_ready),
    .io_right_out_valid(cols_6_2_io_right_out_valid),
    .io_right_out_bits(cols_6_2_io_right_out_bits),
    .io_bottom_out_ready(cols_6_2_io_bottom_out_ready),
    .io_bottom_out_valid(cols_6_2_io_bottom_out_valid),
    .io_bottom_out_bits(cols_6_2_io_bottom_out_bits)
  );
  ProcessingElement cols_7_2 ( // @[Stab.scala 85:60]
    .clock(cols_7_2_clock),
    .reset(cols_7_2_reset),
    .io_left_in_ready(cols_7_2_io_left_in_ready),
    .io_left_in_valid(cols_7_2_io_left_in_valid),
    .io_left_in_bits(cols_7_2_io_left_in_bits),
    .io_top_in_ready(cols_7_2_io_top_in_ready),
    .io_top_in_valid(cols_7_2_io_top_in_valid),
    .io_top_in_bits(cols_7_2_io_top_in_bits),
    .io_sum_ready(cols_7_2_io_sum_ready),
    .io_sum_valid(cols_7_2_io_sum_valid),
    .io_sum_bits(cols_7_2_io_sum_bits),
    .io_right_out_ready(cols_7_2_io_right_out_ready),
    .io_right_out_valid(cols_7_2_io_right_out_valid),
    .io_right_out_bits(cols_7_2_io_right_out_bits),
    .io_bottom_out_ready(cols_7_2_io_bottom_out_ready),
    .io_bottom_out_valid(cols_7_2_io_bottom_out_valid),
    .io_bottom_out_bits(cols_7_2_io_bottom_out_bits)
  );
  ProcessingElement cols_8_2 ( // @[Stab.scala 85:60]
    .clock(cols_8_2_clock),
    .reset(cols_8_2_reset),
    .io_left_in_ready(cols_8_2_io_left_in_ready),
    .io_left_in_valid(cols_8_2_io_left_in_valid),
    .io_left_in_bits(cols_8_2_io_left_in_bits),
    .io_top_in_ready(cols_8_2_io_top_in_ready),
    .io_top_in_valid(cols_8_2_io_top_in_valid),
    .io_top_in_bits(cols_8_2_io_top_in_bits),
    .io_sum_ready(cols_8_2_io_sum_ready),
    .io_sum_valid(cols_8_2_io_sum_valid),
    .io_sum_bits(cols_8_2_io_sum_bits),
    .io_right_out_ready(cols_8_2_io_right_out_ready),
    .io_right_out_valid(cols_8_2_io_right_out_valid),
    .io_right_out_bits(cols_8_2_io_right_out_bits),
    .io_bottom_out_ready(cols_8_2_io_bottom_out_ready),
    .io_bottom_out_valid(cols_8_2_io_bottom_out_valid),
    .io_bottom_out_bits(cols_8_2_io_bottom_out_bits)
  );
  ProcessingElement cols_9_2 ( // @[Stab.scala 85:60]
    .clock(cols_9_2_clock),
    .reset(cols_9_2_reset),
    .io_left_in_ready(cols_9_2_io_left_in_ready),
    .io_left_in_valid(cols_9_2_io_left_in_valid),
    .io_left_in_bits(cols_9_2_io_left_in_bits),
    .io_top_in_ready(cols_9_2_io_top_in_ready),
    .io_top_in_valid(cols_9_2_io_top_in_valid),
    .io_top_in_bits(cols_9_2_io_top_in_bits),
    .io_sum_ready(cols_9_2_io_sum_ready),
    .io_sum_valid(cols_9_2_io_sum_valid),
    .io_sum_bits(cols_9_2_io_sum_bits),
    .io_right_out_ready(cols_9_2_io_right_out_ready),
    .io_right_out_valid(cols_9_2_io_right_out_valid),
    .io_right_out_bits(cols_9_2_io_right_out_bits),
    .io_bottom_out_ready(cols_9_2_io_bottom_out_ready),
    .io_bottom_out_valid(cols_9_2_io_bottom_out_valid),
    .io_bottom_out_bits(cols_9_2_io_bottom_out_bits)
  );
  ProcessingElement cols_10_2 ( // @[Stab.scala 85:60]
    .clock(cols_10_2_clock),
    .reset(cols_10_2_reset),
    .io_left_in_ready(cols_10_2_io_left_in_ready),
    .io_left_in_valid(cols_10_2_io_left_in_valid),
    .io_left_in_bits(cols_10_2_io_left_in_bits),
    .io_top_in_ready(cols_10_2_io_top_in_ready),
    .io_top_in_valid(cols_10_2_io_top_in_valid),
    .io_top_in_bits(cols_10_2_io_top_in_bits),
    .io_sum_ready(cols_10_2_io_sum_ready),
    .io_sum_valid(cols_10_2_io_sum_valid),
    .io_sum_bits(cols_10_2_io_sum_bits),
    .io_right_out_ready(cols_10_2_io_right_out_ready),
    .io_right_out_valid(cols_10_2_io_right_out_valid),
    .io_right_out_bits(cols_10_2_io_right_out_bits),
    .io_bottom_out_ready(cols_10_2_io_bottom_out_ready),
    .io_bottom_out_valid(cols_10_2_io_bottom_out_valid),
    .io_bottom_out_bits(cols_10_2_io_bottom_out_bits)
  );
  ProcessingElement cols_11_2 ( // @[Stab.scala 85:60]
    .clock(cols_11_2_clock),
    .reset(cols_11_2_reset),
    .io_left_in_ready(cols_11_2_io_left_in_ready),
    .io_left_in_valid(cols_11_2_io_left_in_valid),
    .io_left_in_bits(cols_11_2_io_left_in_bits),
    .io_top_in_ready(cols_11_2_io_top_in_ready),
    .io_top_in_valid(cols_11_2_io_top_in_valid),
    .io_top_in_bits(cols_11_2_io_top_in_bits),
    .io_sum_ready(cols_11_2_io_sum_ready),
    .io_sum_valid(cols_11_2_io_sum_valid),
    .io_sum_bits(cols_11_2_io_sum_bits),
    .io_right_out_ready(cols_11_2_io_right_out_ready),
    .io_right_out_valid(cols_11_2_io_right_out_valid),
    .io_right_out_bits(cols_11_2_io_right_out_bits),
    .io_bottom_out_ready(cols_11_2_io_bottom_out_ready),
    .io_bottom_out_valid(cols_11_2_io_bottom_out_valid),
    .io_bottom_out_bits(cols_11_2_io_bottom_out_bits)
  );
  ProcessingElement cols_12_2 ( // @[Stab.scala 85:60]
    .clock(cols_12_2_clock),
    .reset(cols_12_2_reset),
    .io_left_in_ready(cols_12_2_io_left_in_ready),
    .io_left_in_valid(cols_12_2_io_left_in_valid),
    .io_left_in_bits(cols_12_2_io_left_in_bits),
    .io_top_in_ready(cols_12_2_io_top_in_ready),
    .io_top_in_valid(cols_12_2_io_top_in_valid),
    .io_top_in_bits(cols_12_2_io_top_in_bits),
    .io_sum_ready(cols_12_2_io_sum_ready),
    .io_sum_valid(cols_12_2_io_sum_valid),
    .io_sum_bits(cols_12_2_io_sum_bits),
    .io_right_out_ready(cols_12_2_io_right_out_ready),
    .io_right_out_valid(cols_12_2_io_right_out_valid),
    .io_right_out_bits(cols_12_2_io_right_out_bits),
    .io_bottom_out_ready(cols_12_2_io_bottom_out_ready),
    .io_bottom_out_valid(cols_12_2_io_bottom_out_valid),
    .io_bottom_out_bits(cols_12_2_io_bottom_out_bits)
  );
  ProcessingElement cols_13_2 ( // @[Stab.scala 85:60]
    .clock(cols_13_2_clock),
    .reset(cols_13_2_reset),
    .io_left_in_ready(cols_13_2_io_left_in_ready),
    .io_left_in_valid(cols_13_2_io_left_in_valid),
    .io_left_in_bits(cols_13_2_io_left_in_bits),
    .io_top_in_ready(cols_13_2_io_top_in_ready),
    .io_top_in_valid(cols_13_2_io_top_in_valid),
    .io_top_in_bits(cols_13_2_io_top_in_bits),
    .io_sum_ready(cols_13_2_io_sum_ready),
    .io_sum_valid(cols_13_2_io_sum_valid),
    .io_sum_bits(cols_13_2_io_sum_bits),
    .io_right_out_ready(cols_13_2_io_right_out_ready),
    .io_right_out_valid(cols_13_2_io_right_out_valid),
    .io_right_out_bits(cols_13_2_io_right_out_bits),
    .io_bottom_out_ready(cols_13_2_io_bottom_out_ready),
    .io_bottom_out_valid(cols_13_2_io_bottom_out_valid),
    .io_bottom_out_bits(cols_13_2_io_bottom_out_bits)
  );
  ProcessingElement cols_14_2 ( // @[Stab.scala 85:60]
    .clock(cols_14_2_clock),
    .reset(cols_14_2_reset),
    .io_left_in_ready(cols_14_2_io_left_in_ready),
    .io_left_in_valid(cols_14_2_io_left_in_valid),
    .io_left_in_bits(cols_14_2_io_left_in_bits),
    .io_top_in_ready(cols_14_2_io_top_in_ready),
    .io_top_in_valid(cols_14_2_io_top_in_valid),
    .io_top_in_bits(cols_14_2_io_top_in_bits),
    .io_sum_ready(cols_14_2_io_sum_ready),
    .io_sum_valid(cols_14_2_io_sum_valid),
    .io_sum_bits(cols_14_2_io_sum_bits),
    .io_right_out_ready(cols_14_2_io_right_out_ready),
    .io_right_out_valid(cols_14_2_io_right_out_valid),
    .io_right_out_bits(cols_14_2_io_right_out_bits),
    .io_bottom_out_ready(cols_14_2_io_bottom_out_ready),
    .io_bottom_out_valid(cols_14_2_io_bottom_out_valid),
    .io_bottom_out_bits(cols_14_2_io_bottom_out_bits)
  );
  ProcessingElement cols_15_2 ( // @[Stab.scala 85:60]
    .clock(cols_15_2_clock),
    .reset(cols_15_2_reset),
    .io_left_in_ready(cols_15_2_io_left_in_ready),
    .io_left_in_valid(cols_15_2_io_left_in_valid),
    .io_left_in_bits(cols_15_2_io_left_in_bits),
    .io_top_in_ready(cols_15_2_io_top_in_ready),
    .io_top_in_valid(cols_15_2_io_top_in_valid),
    .io_top_in_bits(cols_15_2_io_top_in_bits),
    .io_sum_ready(cols_15_2_io_sum_ready),
    .io_sum_valid(cols_15_2_io_sum_valid),
    .io_sum_bits(cols_15_2_io_sum_bits),
    .io_right_out_ready(cols_15_2_io_right_out_ready),
    .io_right_out_valid(cols_15_2_io_right_out_valid),
    .io_right_out_bits(cols_15_2_io_right_out_bits),
    .io_bottom_out_ready(cols_15_2_io_bottom_out_ready),
    .io_bottom_out_valid(cols_15_2_io_bottom_out_valid),
    .io_bottom_out_bits(cols_15_2_io_bottom_out_bits)
  );
  ProcessingElement cols_0_3 ( // @[Stab.scala 85:60]
    .clock(cols_0_3_clock),
    .reset(cols_0_3_reset),
    .io_left_in_ready(cols_0_3_io_left_in_ready),
    .io_left_in_valid(cols_0_3_io_left_in_valid),
    .io_left_in_bits(cols_0_3_io_left_in_bits),
    .io_top_in_ready(cols_0_3_io_top_in_ready),
    .io_top_in_valid(cols_0_3_io_top_in_valid),
    .io_top_in_bits(cols_0_3_io_top_in_bits),
    .io_sum_ready(cols_0_3_io_sum_ready),
    .io_sum_valid(cols_0_3_io_sum_valid),
    .io_sum_bits(cols_0_3_io_sum_bits),
    .io_right_out_ready(cols_0_3_io_right_out_ready),
    .io_right_out_valid(cols_0_3_io_right_out_valid),
    .io_right_out_bits(cols_0_3_io_right_out_bits),
    .io_bottom_out_ready(cols_0_3_io_bottom_out_ready),
    .io_bottom_out_valid(cols_0_3_io_bottom_out_valid),
    .io_bottom_out_bits(cols_0_3_io_bottom_out_bits)
  );
  ProcessingElement cols_1_3 ( // @[Stab.scala 85:60]
    .clock(cols_1_3_clock),
    .reset(cols_1_3_reset),
    .io_left_in_ready(cols_1_3_io_left_in_ready),
    .io_left_in_valid(cols_1_3_io_left_in_valid),
    .io_left_in_bits(cols_1_3_io_left_in_bits),
    .io_top_in_ready(cols_1_3_io_top_in_ready),
    .io_top_in_valid(cols_1_3_io_top_in_valid),
    .io_top_in_bits(cols_1_3_io_top_in_bits),
    .io_sum_ready(cols_1_3_io_sum_ready),
    .io_sum_valid(cols_1_3_io_sum_valid),
    .io_sum_bits(cols_1_3_io_sum_bits),
    .io_right_out_ready(cols_1_3_io_right_out_ready),
    .io_right_out_valid(cols_1_3_io_right_out_valid),
    .io_right_out_bits(cols_1_3_io_right_out_bits),
    .io_bottom_out_ready(cols_1_3_io_bottom_out_ready),
    .io_bottom_out_valid(cols_1_3_io_bottom_out_valid),
    .io_bottom_out_bits(cols_1_3_io_bottom_out_bits)
  );
  ProcessingElement cols_2_3 ( // @[Stab.scala 85:60]
    .clock(cols_2_3_clock),
    .reset(cols_2_3_reset),
    .io_left_in_ready(cols_2_3_io_left_in_ready),
    .io_left_in_valid(cols_2_3_io_left_in_valid),
    .io_left_in_bits(cols_2_3_io_left_in_bits),
    .io_top_in_ready(cols_2_3_io_top_in_ready),
    .io_top_in_valid(cols_2_3_io_top_in_valid),
    .io_top_in_bits(cols_2_3_io_top_in_bits),
    .io_sum_ready(cols_2_3_io_sum_ready),
    .io_sum_valid(cols_2_3_io_sum_valid),
    .io_sum_bits(cols_2_3_io_sum_bits),
    .io_right_out_ready(cols_2_3_io_right_out_ready),
    .io_right_out_valid(cols_2_3_io_right_out_valid),
    .io_right_out_bits(cols_2_3_io_right_out_bits),
    .io_bottom_out_ready(cols_2_3_io_bottom_out_ready),
    .io_bottom_out_valid(cols_2_3_io_bottom_out_valid),
    .io_bottom_out_bits(cols_2_3_io_bottom_out_bits)
  );
  ProcessingElement cols_3_3 ( // @[Stab.scala 85:60]
    .clock(cols_3_3_clock),
    .reset(cols_3_3_reset),
    .io_left_in_ready(cols_3_3_io_left_in_ready),
    .io_left_in_valid(cols_3_3_io_left_in_valid),
    .io_left_in_bits(cols_3_3_io_left_in_bits),
    .io_top_in_ready(cols_3_3_io_top_in_ready),
    .io_top_in_valid(cols_3_3_io_top_in_valid),
    .io_top_in_bits(cols_3_3_io_top_in_bits),
    .io_sum_ready(cols_3_3_io_sum_ready),
    .io_sum_valid(cols_3_3_io_sum_valid),
    .io_sum_bits(cols_3_3_io_sum_bits),
    .io_right_out_ready(cols_3_3_io_right_out_ready),
    .io_right_out_valid(cols_3_3_io_right_out_valid),
    .io_right_out_bits(cols_3_3_io_right_out_bits),
    .io_bottom_out_ready(cols_3_3_io_bottom_out_ready),
    .io_bottom_out_valid(cols_3_3_io_bottom_out_valid),
    .io_bottom_out_bits(cols_3_3_io_bottom_out_bits)
  );
  ProcessingElement cols_4_3 ( // @[Stab.scala 85:60]
    .clock(cols_4_3_clock),
    .reset(cols_4_3_reset),
    .io_left_in_ready(cols_4_3_io_left_in_ready),
    .io_left_in_valid(cols_4_3_io_left_in_valid),
    .io_left_in_bits(cols_4_3_io_left_in_bits),
    .io_top_in_ready(cols_4_3_io_top_in_ready),
    .io_top_in_valid(cols_4_3_io_top_in_valid),
    .io_top_in_bits(cols_4_3_io_top_in_bits),
    .io_sum_ready(cols_4_3_io_sum_ready),
    .io_sum_valid(cols_4_3_io_sum_valid),
    .io_sum_bits(cols_4_3_io_sum_bits),
    .io_right_out_ready(cols_4_3_io_right_out_ready),
    .io_right_out_valid(cols_4_3_io_right_out_valid),
    .io_right_out_bits(cols_4_3_io_right_out_bits),
    .io_bottom_out_ready(cols_4_3_io_bottom_out_ready),
    .io_bottom_out_valid(cols_4_3_io_bottom_out_valid),
    .io_bottom_out_bits(cols_4_3_io_bottom_out_bits)
  );
  ProcessingElement cols_5_3 ( // @[Stab.scala 85:60]
    .clock(cols_5_3_clock),
    .reset(cols_5_3_reset),
    .io_left_in_ready(cols_5_3_io_left_in_ready),
    .io_left_in_valid(cols_5_3_io_left_in_valid),
    .io_left_in_bits(cols_5_3_io_left_in_bits),
    .io_top_in_ready(cols_5_3_io_top_in_ready),
    .io_top_in_valid(cols_5_3_io_top_in_valid),
    .io_top_in_bits(cols_5_3_io_top_in_bits),
    .io_sum_ready(cols_5_3_io_sum_ready),
    .io_sum_valid(cols_5_3_io_sum_valid),
    .io_sum_bits(cols_5_3_io_sum_bits),
    .io_right_out_ready(cols_5_3_io_right_out_ready),
    .io_right_out_valid(cols_5_3_io_right_out_valid),
    .io_right_out_bits(cols_5_3_io_right_out_bits),
    .io_bottom_out_ready(cols_5_3_io_bottom_out_ready),
    .io_bottom_out_valid(cols_5_3_io_bottom_out_valid),
    .io_bottom_out_bits(cols_5_3_io_bottom_out_bits)
  );
  ProcessingElement cols_6_3 ( // @[Stab.scala 85:60]
    .clock(cols_6_3_clock),
    .reset(cols_6_3_reset),
    .io_left_in_ready(cols_6_3_io_left_in_ready),
    .io_left_in_valid(cols_6_3_io_left_in_valid),
    .io_left_in_bits(cols_6_3_io_left_in_bits),
    .io_top_in_ready(cols_6_3_io_top_in_ready),
    .io_top_in_valid(cols_6_3_io_top_in_valid),
    .io_top_in_bits(cols_6_3_io_top_in_bits),
    .io_sum_ready(cols_6_3_io_sum_ready),
    .io_sum_valid(cols_6_3_io_sum_valid),
    .io_sum_bits(cols_6_3_io_sum_bits),
    .io_right_out_ready(cols_6_3_io_right_out_ready),
    .io_right_out_valid(cols_6_3_io_right_out_valid),
    .io_right_out_bits(cols_6_3_io_right_out_bits),
    .io_bottom_out_ready(cols_6_3_io_bottom_out_ready),
    .io_bottom_out_valid(cols_6_3_io_bottom_out_valid),
    .io_bottom_out_bits(cols_6_3_io_bottom_out_bits)
  );
  ProcessingElement cols_7_3 ( // @[Stab.scala 85:60]
    .clock(cols_7_3_clock),
    .reset(cols_7_3_reset),
    .io_left_in_ready(cols_7_3_io_left_in_ready),
    .io_left_in_valid(cols_7_3_io_left_in_valid),
    .io_left_in_bits(cols_7_3_io_left_in_bits),
    .io_top_in_ready(cols_7_3_io_top_in_ready),
    .io_top_in_valid(cols_7_3_io_top_in_valid),
    .io_top_in_bits(cols_7_3_io_top_in_bits),
    .io_sum_ready(cols_7_3_io_sum_ready),
    .io_sum_valid(cols_7_3_io_sum_valid),
    .io_sum_bits(cols_7_3_io_sum_bits),
    .io_right_out_ready(cols_7_3_io_right_out_ready),
    .io_right_out_valid(cols_7_3_io_right_out_valid),
    .io_right_out_bits(cols_7_3_io_right_out_bits),
    .io_bottom_out_ready(cols_7_3_io_bottom_out_ready),
    .io_bottom_out_valid(cols_7_3_io_bottom_out_valid),
    .io_bottom_out_bits(cols_7_3_io_bottom_out_bits)
  );
  ProcessingElement cols_8_3 ( // @[Stab.scala 85:60]
    .clock(cols_8_3_clock),
    .reset(cols_8_3_reset),
    .io_left_in_ready(cols_8_3_io_left_in_ready),
    .io_left_in_valid(cols_8_3_io_left_in_valid),
    .io_left_in_bits(cols_8_3_io_left_in_bits),
    .io_top_in_ready(cols_8_3_io_top_in_ready),
    .io_top_in_valid(cols_8_3_io_top_in_valid),
    .io_top_in_bits(cols_8_3_io_top_in_bits),
    .io_sum_ready(cols_8_3_io_sum_ready),
    .io_sum_valid(cols_8_3_io_sum_valid),
    .io_sum_bits(cols_8_3_io_sum_bits),
    .io_right_out_ready(cols_8_3_io_right_out_ready),
    .io_right_out_valid(cols_8_3_io_right_out_valid),
    .io_right_out_bits(cols_8_3_io_right_out_bits),
    .io_bottom_out_ready(cols_8_3_io_bottom_out_ready),
    .io_bottom_out_valid(cols_8_3_io_bottom_out_valid),
    .io_bottom_out_bits(cols_8_3_io_bottom_out_bits)
  );
  ProcessingElement cols_9_3 ( // @[Stab.scala 85:60]
    .clock(cols_9_3_clock),
    .reset(cols_9_3_reset),
    .io_left_in_ready(cols_9_3_io_left_in_ready),
    .io_left_in_valid(cols_9_3_io_left_in_valid),
    .io_left_in_bits(cols_9_3_io_left_in_bits),
    .io_top_in_ready(cols_9_3_io_top_in_ready),
    .io_top_in_valid(cols_9_3_io_top_in_valid),
    .io_top_in_bits(cols_9_3_io_top_in_bits),
    .io_sum_ready(cols_9_3_io_sum_ready),
    .io_sum_valid(cols_9_3_io_sum_valid),
    .io_sum_bits(cols_9_3_io_sum_bits),
    .io_right_out_ready(cols_9_3_io_right_out_ready),
    .io_right_out_valid(cols_9_3_io_right_out_valid),
    .io_right_out_bits(cols_9_3_io_right_out_bits),
    .io_bottom_out_ready(cols_9_3_io_bottom_out_ready),
    .io_bottom_out_valid(cols_9_3_io_bottom_out_valid),
    .io_bottom_out_bits(cols_9_3_io_bottom_out_bits)
  );
  ProcessingElement cols_10_3 ( // @[Stab.scala 85:60]
    .clock(cols_10_3_clock),
    .reset(cols_10_3_reset),
    .io_left_in_ready(cols_10_3_io_left_in_ready),
    .io_left_in_valid(cols_10_3_io_left_in_valid),
    .io_left_in_bits(cols_10_3_io_left_in_bits),
    .io_top_in_ready(cols_10_3_io_top_in_ready),
    .io_top_in_valid(cols_10_3_io_top_in_valid),
    .io_top_in_bits(cols_10_3_io_top_in_bits),
    .io_sum_ready(cols_10_3_io_sum_ready),
    .io_sum_valid(cols_10_3_io_sum_valid),
    .io_sum_bits(cols_10_3_io_sum_bits),
    .io_right_out_ready(cols_10_3_io_right_out_ready),
    .io_right_out_valid(cols_10_3_io_right_out_valid),
    .io_right_out_bits(cols_10_3_io_right_out_bits),
    .io_bottom_out_ready(cols_10_3_io_bottom_out_ready),
    .io_bottom_out_valid(cols_10_3_io_bottom_out_valid),
    .io_bottom_out_bits(cols_10_3_io_bottom_out_bits)
  );
  ProcessingElement cols_11_3 ( // @[Stab.scala 85:60]
    .clock(cols_11_3_clock),
    .reset(cols_11_3_reset),
    .io_left_in_ready(cols_11_3_io_left_in_ready),
    .io_left_in_valid(cols_11_3_io_left_in_valid),
    .io_left_in_bits(cols_11_3_io_left_in_bits),
    .io_top_in_ready(cols_11_3_io_top_in_ready),
    .io_top_in_valid(cols_11_3_io_top_in_valid),
    .io_top_in_bits(cols_11_3_io_top_in_bits),
    .io_sum_ready(cols_11_3_io_sum_ready),
    .io_sum_valid(cols_11_3_io_sum_valid),
    .io_sum_bits(cols_11_3_io_sum_bits),
    .io_right_out_ready(cols_11_3_io_right_out_ready),
    .io_right_out_valid(cols_11_3_io_right_out_valid),
    .io_right_out_bits(cols_11_3_io_right_out_bits),
    .io_bottom_out_ready(cols_11_3_io_bottom_out_ready),
    .io_bottom_out_valid(cols_11_3_io_bottom_out_valid),
    .io_bottom_out_bits(cols_11_3_io_bottom_out_bits)
  );
  ProcessingElement cols_12_3 ( // @[Stab.scala 85:60]
    .clock(cols_12_3_clock),
    .reset(cols_12_3_reset),
    .io_left_in_ready(cols_12_3_io_left_in_ready),
    .io_left_in_valid(cols_12_3_io_left_in_valid),
    .io_left_in_bits(cols_12_3_io_left_in_bits),
    .io_top_in_ready(cols_12_3_io_top_in_ready),
    .io_top_in_valid(cols_12_3_io_top_in_valid),
    .io_top_in_bits(cols_12_3_io_top_in_bits),
    .io_sum_ready(cols_12_3_io_sum_ready),
    .io_sum_valid(cols_12_3_io_sum_valid),
    .io_sum_bits(cols_12_3_io_sum_bits),
    .io_right_out_ready(cols_12_3_io_right_out_ready),
    .io_right_out_valid(cols_12_3_io_right_out_valid),
    .io_right_out_bits(cols_12_3_io_right_out_bits),
    .io_bottom_out_ready(cols_12_3_io_bottom_out_ready),
    .io_bottom_out_valid(cols_12_3_io_bottom_out_valid),
    .io_bottom_out_bits(cols_12_3_io_bottom_out_bits)
  );
  ProcessingElement cols_13_3 ( // @[Stab.scala 85:60]
    .clock(cols_13_3_clock),
    .reset(cols_13_3_reset),
    .io_left_in_ready(cols_13_3_io_left_in_ready),
    .io_left_in_valid(cols_13_3_io_left_in_valid),
    .io_left_in_bits(cols_13_3_io_left_in_bits),
    .io_top_in_ready(cols_13_3_io_top_in_ready),
    .io_top_in_valid(cols_13_3_io_top_in_valid),
    .io_top_in_bits(cols_13_3_io_top_in_bits),
    .io_sum_ready(cols_13_3_io_sum_ready),
    .io_sum_valid(cols_13_3_io_sum_valid),
    .io_sum_bits(cols_13_3_io_sum_bits),
    .io_right_out_ready(cols_13_3_io_right_out_ready),
    .io_right_out_valid(cols_13_3_io_right_out_valid),
    .io_right_out_bits(cols_13_3_io_right_out_bits),
    .io_bottom_out_ready(cols_13_3_io_bottom_out_ready),
    .io_bottom_out_valid(cols_13_3_io_bottom_out_valid),
    .io_bottom_out_bits(cols_13_3_io_bottom_out_bits)
  );
  ProcessingElement cols_14_3 ( // @[Stab.scala 85:60]
    .clock(cols_14_3_clock),
    .reset(cols_14_3_reset),
    .io_left_in_ready(cols_14_3_io_left_in_ready),
    .io_left_in_valid(cols_14_3_io_left_in_valid),
    .io_left_in_bits(cols_14_3_io_left_in_bits),
    .io_top_in_ready(cols_14_3_io_top_in_ready),
    .io_top_in_valid(cols_14_3_io_top_in_valid),
    .io_top_in_bits(cols_14_3_io_top_in_bits),
    .io_sum_ready(cols_14_3_io_sum_ready),
    .io_sum_valid(cols_14_3_io_sum_valid),
    .io_sum_bits(cols_14_3_io_sum_bits),
    .io_right_out_ready(cols_14_3_io_right_out_ready),
    .io_right_out_valid(cols_14_3_io_right_out_valid),
    .io_right_out_bits(cols_14_3_io_right_out_bits),
    .io_bottom_out_ready(cols_14_3_io_bottom_out_ready),
    .io_bottom_out_valid(cols_14_3_io_bottom_out_valid),
    .io_bottom_out_bits(cols_14_3_io_bottom_out_bits)
  );
  ProcessingElement cols_15_3 ( // @[Stab.scala 85:60]
    .clock(cols_15_3_clock),
    .reset(cols_15_3_reset),
    .io_left_in_ready(cols_15_3_io_left_in_ready),
    .io_left_in_valid(cols_15_3_io_left_in_valid),
    .io_left_in_bits(cols_15_3_io_left_in_bits),
    .io_top_in_ready(cols_15_3_io_top_in_ready),
    .io_top_in_valid(cols_15_3_io_top_in_valid),
    .io_top_in_bits(cols_15_3_io_top_in_bits),
    .io_sum_ready(cols_15_3_io_sum_ready),
    .io_sum_valid(cols_15_3_io_sum_valid),
    .io_sum_bits(cols_15_3_io_sum_bits),
    .io_right_out_ready(cols_15_3_io_right_out_ready),
    .io_right_out_valid(cols_15_3_io_right_out_valid),
    .io_right_out_bits(cols_15_3_io_right_out_bits),
    .io_bottom_out_ready(cols_15_3_io_bottom_out_ready),
    .io_bottom_out_valid(cols_15_3_io_bottom_out_valid),
    .io_bottom_out_bits(cols_15_3_io_bottom_out_bits)
  );
  ProcessingElement cols_0_4 ( // @[Stab.scala 85:60]
    .clock(cols_0_4_clock),
    .reset(cols_0_4_reset),
    .io_left_in_ready(cols_0_4_io_left_in_ready),
    .io_left_in_valid(cols_0_4_io_left_in_valid),
    .io_left_in_bits(cols_0_4_io_left_in_bits),
    .io_top_in_ready(cols_0_4_io_top_in_ready),
    .io_top_in_valid(cols_0_4_io_top_in_valid),
    .io_top_in_bits(cols_0_4_io_top_in_bits),
    .io_sum_ready(cols_0_4_io_sum_ready),
    .io_sum_valid(cols_0_4_io_sum_valid),
    .io_sum_bits(cols_0_4_io_sum_bits),
    .io_right_out_ready(cols_0_4_io_right_out_ready),
    .io_right_out_valid(cols_0_4_io_right_out_valid),
    .io_right_out_bits(cols_0_4_io_right_out_bits),
    .io_bottom_out_ready(cols_0_4_io_bottom_out_ready),
    .io_bottom_out_valid(cols_0_4_io_bottom_out_valid),
    .io_bottom_out_bits(cols_0_4_io_bottom_out_bits)
  );
  ProcessingElement cols_1_4 ( // @[Stab.scala 85:60]
    .clock(cols_1_4_clock),
    .reset(cols_1_4_reset),
    .io_left_in_ready(cols_1_4_io_left_in_ready),
    .io_left_in_valid(cols_1_4_io_left_in_valid),
    .io_left_in_bits(cols_1_4_io_left_in_bits),
    .io_top_in_ready(cols_1_4_io_top_in_ready),
    .io_top_in_valid(cols_1_4_io_top_in_valid),
    .io_top_in_bits(cols_1_4_io_top_in_bits),
    .io_sum_ready(cols_1_4_io_sum_ready),
    .io_sum_valid(cols_1_4_io_sum_valid),
    .io_sum_bits(cols_1_4_io_sum_bits),
    .io_right_out_ready(cols_1_4_io_right_out_ready),
    .io_right_out_valid(cols_1_4_io_right_out_valid),
    .io_right_out_bits(cols_1_4_io_right_out_bits),
    .io_bottom_out_ready(cols_1_4_io_bottom_out_ready),
    .io_bottom_out_valid(cols_1_4_io_bottom_out_valid),
    .io_bottom_out_bits(cols_1_4_io_bottom_out_bits)
  );
  ProcessingElement cols_2_4 ( // @[Stab.scala 85:60]
    .clock(cols_2_4_clock),
    .reset(cols_2_4_reset),
    .io_left_in_ready(cols_2_4_io_left_in_ready),
    .io_left_in_valid(cols_2_4_io_left_in_valid),
    .io_left_in_bits(cols_2_4_io_left_in_bits),
    .io_top_in_ready(cols_2_4_io_top_in_ready),
    .io_top_in_valid(cols_2_4_io_top_in_valid),
    .io_top_in_bits(cols_2_4_io_top_in_bits),
    .io_sum_ready(cols_2_4_io_sum_ready),
    .io_sum_valid(cols_2_4_io_sum_valid),
    .io_sum_bits(cols_2_4_io_sum_bits),
    .io_right_out_ready(cols_2_4_io_right_out_ready),
    .io_right_out_valid(cols_2_4_io_right_out_valid),
    .io_right_out_bits(cols_2_4_io_right_out_bits),
    .io_bottom_out_ready(cols_2_4_io_bottom_out_ready),
    .io_bottom_out_valid(cols_2_4_io_bottom_out_valid),
    .io_bottom_out_bits(cols_2_4_io_bottom_out_bits)
  );
  ProcessingElement cols_3_4 ( // @[Stab.scala 85:60]
    .clock(cols_3_4_clock),
    .reset(cols_3_4_reset),
    .io_left_in_ready(cols_3_4_io_left_in_ready),
    .io_left_in_valid(cols_3_4_io_left_in_valid),
    .io_left_in_bits(cols_3_4_io_left_in_bits),
    .io_top_in_ready(cols_3_4_io_top_in_ready),
    .io_top_in_valid(cols_3_4_io_top_in_valid),
    .io_top_in_bits(cols_3_4_io_top_in_bits),
    .io_sum_ready(cols_3_4_io_sum_ready),
    .io_sum_valid(cols_3_4_io_sum_valid),
    .io_sum_bits(cols_3_4_io_sum_bits),
    .io_right_out_ready(cols_3_4_io_right_out_ready),
    .io_right_out_valid(cols_3_4_io_right_out_valid),
    .io_right_out_bits(cols_3_4_io_right_out_bits),
    .io_bottom_out_ready(cols_3_4_io_bottom_out_ready),
    .io_bottom_out_valid(cols_3_4_io_bottom_out_valid),
    .io_bottom_out_bits(cols_3_4_io_bottom_out_bits)
  );
  ProcessingElement cols_4_4 ( // @[Stab.scala 85:60]
    .clock(cols_4_4_clock),
    .reset(cols_4_4_reset),
    .io_left_in_ready(cols_4_4_io_left_in_ready),
    .io_left_in_valid(cols_4_4_io_left_in_valid),
    .io_left_in_bits(cols_4_4_io_left_in_bits),
    .io_top_in_ready(cols_4_4_io_top_in_ready),
    .io_top_in_valid(cols_4_4_io_top_in_valid),
    .io_top_in_bits(cols_4_4_io_top_in_bits),
    .io_sum_ready(cols_4_4_io_sum_ready),
    .io_sum_valid(cols_4_4_io_sum_valid),
    .io_sum_bits(cols_4_4_io_sum_bits),
    .io_right_out_ready(cols_4_4_io_right_out_ready),
    .io_right_out_valid(cols_4_4_io_right_out_valid),
    .io_right_out_bits(cols_4_4_io_right_out_bits),
    .io_bottom_out_ready(cols_4_4_io_bottom_out_ready),
    .io_bottom_out_valid(cols_4_4_io_bottom_out_valid),
    .io_bottom_out_bits(cols_4_4_io_bottom_out_bits)
  );
  ProcessingElement cols_5_4 ( // @[Stab.scala 85:60]
    .clock(cols_5_4_clock),
    .reset(cols_5_4_reset),
    .io_left_in_ready(cols_5_4_io_left_in_ready),
    .io_left_in_valid(cols_5_4_io_left_in_valid),
    .io_left_in_bits(cols_5_4_io_left_in_bits),
    .io_top_in_ready(cols_5_4_io_top_in_ready),
    .io_top_in_valid(cols_5_4_io_top_in_valid),
    .io_top_in_bits(cols_5_4_io_top_in_bits),
    .io_sum_ready(cols_5_4_io_sum_ready),
    .io_sum_valid(cols_5_4_io_sum_valid),
    .io_sum_bits(cols_5_4_io_sum_bits),
    .io_right_out_ready(cols_5_4_io_right_out_ready),
    .io_right_out_valid(cols_5_4_io_right_out_valid),
    .io_right_out_bits(cols_5_4_io_right_out_bits),
    .io_bottom_out_ready(cols_5_4_io_bottom_out_ready),
    .io_bottom_out_valid(cols_5_4_io_bottom_out_valid),
    .io_bottom_out_bits(cols_5_4_io_bottom_out_bits)
  );
  ProcessingElement cols_6_4 ( // @[Stab.scala 85:60]
    .clock(cols_6_4_clock),
    .reset(cols_6_4_reset),
    .io_left_in_ready(cols_6_4_io_left_in_ready),
    .io_left_in_valid(cols_6_4_io_left_in_valid),
    .io_left_in_bits(cols_6_4_io_left_in_bits),
    .io_top_in_ready(cols_6_4_io_top_in_ready),
    .io_top_in_valid(cols_6_4_io_top_in_valid),
    .io_top_in_bits(cols_6_4_io_top_in_bits),
    .io_sum_ready(cols_6_4_io_sum_ready),
    .io_sum_valid(cols_6_4_io_sum_valid),
    .io_sum_bits(cols_6_4_io_sum_bits),
    .io_right_out_ready(cols_6_4_io_right_out_ready),
    .io_right_out_valid(cols_6_4_io_right_out_valid),
    .io_right_out_bits(cols_6_4_io_right_out_bits),
    .io_bottom_out_ready(cols_6_4_io_bottom_out_ready),
    .io_bottom_out_valid(cols_6_4_io_bottom_out_valid),
    .io_bottom_out_bits(cols_6_4_io_bottom_out_bits)
  );
  ProcessingElement cols_7_4 ( // @[Stab.scala 85:60]
    .clock(cols_7_4_clock),
    .reset(cols_7_4_reset),
    .io_left_in_ready(cols_7_4_io_left_in_ready),
    .io_left_in_valid(cols_7_4_io_left_in_valid),
    .io_left_in_bits(cols_7_4_io_left_in_bits),
    .io_top_in_ready(cols_7_4_io_top_in_ready),
    .io_top_in_valid(cols_7_4_io_top_in_valid),
    .io_top_in_bits(cols_7_4_io_top_in_bits),
    .io_sum_ready(cols_7_4_io_sum_ready),
    .io_sum_valid(cols_7_4_io_sum_valid),
    .io_sum_bits(cols_7_4_io_sum_bits),
    .io_right_out_ready(cols_7_4_io_right_out_ready),
    .io_right_out_valid(cols_7_4_io_right_out_valid),
    .io_right_out_bits(cols_7_4_io_right_out_bits),
    .io_bottom_out_ready(cols_7_4_io_bottom_out_ready),
    .io_bottom_out_valid(cols_7_4_io_bottom_out_valid),
    .io_bottom_out_bits(cols_7_4_io_bottom_out_bits)
  );
  ProcessingElement cols_8_4 ( // @[Stab.scala 85:60]
    .clock(cols_8_4_clock),
    .reset(cols_8_4_reset),
    .io_left_in_ready(cols_8_4_io_left_in_ready),
    .io_left_in_valid(cols_8_4_io_left_in_valid),
    .io_left_in_bits(cols_8_4_io_left_in_bits),
    .io_top_in_ready(cols_8_4_io_top_in_ready),
    .io_top_in_valid(cols_8_4_io_top_in_valid),
    .io_top_in_bits(cols_8_4_io_top_in_bits),
    .io_sum_ready(cols_8_4_io_sum_ready),
    .io_sum_valid(cols_8_4_io_sum_valid),
    .io_sum_bits(cols_8_4_io_sum_bits),
    .io_right_out_ready(cols_8_4_io_right_out_ready),
    .io_right_out_valid(cols_8_4_io_right_out_valid),
    .io_right_out_bits(cols_8_4_io_right_out_bits),
    .io_bottom_out_ready(cols_8_4_io_bottom_out_ready),
    .io_bottom_out_valid(cols_8_4_io_bottom_out_valid),
    .io_bottom_out_bits(cols_8_4_io_bottom_out_bits)
  );
  ProcessingElement cols_9_4 ( // @[Stab.scala 85:60]
    .clock(cols_9_4_clock),
    .reset(cols_9_4_reset),
    .io_left_in_ready(cols_9_4_io_left_in_ready),
    .io_left_in_valid(cols_9_4_io_left_in_valid),
    .io_left_in_bits(cols_9_4_io_left_in_bits),
    .io_top_in_ready(cols_9_4_io_top_in_ready),
    .io_top_in_valid(cols_9_4_io_top_in_valid),
    .io_top_in_bits(cols_9_4_io_top_in_bits),
    .io_sum_ready(cols_9_4_io_sum_ready),
    .io_sum_valid(cols_9_4_io_sum_valid),
    .io_sum_bits(cols_9_4_io_sum_bits),
    .io_right_out_ready(cols_9_4_io_right_out_ready),
    .io_right_out_valid(cols_9_4_io_right_out_valid),
    .io_right_out_bits(cols_9_4_io_right_out_bits),
    .io_bottom_out_ready(cols_9_4_io_bottom_out_ready),
    .io_bottom_out_valid(cols_9_4_io_bottom_out_valid),
    .io_bottom_out_bits(cols_9_4_io_bottom_out_bits)
  );
  ProcessingElement cols_10_4 ( // @[Stab.scala 85:60]
    .clock(cols_10_4_clock),
    .reset(cols_10_4_reset),
    .io_left_in_ready(cols_10_4_io_left_in_ready),
    .io_left_in_valid(cols_10_4_io_left_in_valid),
    .io_left_in_bits(cols_10_4_io_left_in_bits),
    .io_top_in_ready(cols_10_4_io_top_in_ready),
    .io_top_in_valid(cols_10_4_io_top_in_valid),
    .io_top_in_bits(cols_10_4_io_top_in_bits),
    .io_sum_ready(cols_10_4_io_sum_ready),
    .io_sum_valid(cols_10_4_io_sum_valid),
    .io_sum_bits(cols_10_4_io_sum_bits),
    .io_right_out_ready(cols_10_4_io_right_out_ready),
    .io_right_out_valid(cols_10_4_io_right_out_valid),
    .io_right_out_bits(cols_10_4_io_right_out_bits),
    .io_bottom_out_ready(cols_10_4_io_bottom_out_ready),
    .io_bottom_out_valid(cols_10_4_io_bottom_out_valid),
    .io_bottom_out_bits(cols_10_4_io_bottom_out_bits)
  );
  ProcessingElement cols_11_4 ( // @[Stab.scala 85:60]
    .clock(cols_11_4_clock),
    .reset(cols_11_4_reset),
    .io_left_in_ready(cols_11_4_io_left_in_ready),
    .io_left_in_valid(cols_11_4_io_left_in_valid),
    .io_left_in_bits(cols_11_4_io_left_in_bits),
    .io_top_in_ready(cols_11_4_io_top_in_ready),
    .io_top_in_valid(cols_11_4_io_top_in_valid),
    .io_top_in_bits(cols_11_4_io_top_in_bits),
    .io_sum_ready(cols_11_4_io_sum_ready),
    .io_sum_valid(cols_11_4_io_sum_valid),
    .io_sum_bits(cols_11_4_io_sum_bits),
    .io_right_out_ready(cols_11_4_io_right_out_ready),
    .io_right_out_valid(cols_11_4_io_right_out_valid),
    .io_right_out_bits(cols_11_4_io_right_out_bits),
    .io_bottom_out_ready(cols_11_4_io_bottom_out_ready),
    .io_bottom_out_valid(cols_11_4_io_bottom_out_valid),
    .io_bottom_out_bits(cols_11_4_io_bottom_out_bits)
  );
  ProcessingElement cols_12_4 ( // @[Stab.scala 85:60]
    .clock(cols_12_4_clock),
    .reset(cols_12_4_reset),
    .io_left_in_ready(cols_12_4_io_left_in_ready),
    .io_left_in_valid(cols_12_4_io_left_in_valid),
    .io_left_in_bits(cols_12_4_io_left_in_bits),
    .io_top_in_ready(cols_12_4_io_top_in_ready),
    .io_top_in_valid(cols_12_4_io_top_in_valid),
    .io_top_in_bits(cols_12_4_io_top_in_bits),
    .io_sum_ready(cols_12_4_io_sum_ready),
    .io_sum_valid(cols_12_4_io_sum_valid),
    .io_sum_bits(cols_12_4_io_sum_bits),
    .io_right_out_ready(cols_12_4_io_right_out_ready),
    .io_right_out_valid(cols_12_4_io_right_out_valid),
    .io_right_out_bits(cols_12_4_io_right_out_bits),
    .io_bottom_out_ready(cols_12_4_io_bottom_out_ready),
    .io_bottom_out_valid(cols_12_4_io_bottom_out_valid),
    .io_bottom_out_bits(cols_12_4_io_bottom_out_bits)
  );
  ProcessingElement cols_13_4 ( // @[Stab.scala 85:60]
    .clock(cols_13_4_clock),
    .reset(cols_13_4_reset),
    .io_left_in_ready(cols_13_4_io_left_in_ready),
    .io_left_in_valid(cols_13_4_io_left_in_valid),
    .io_left_in_bits(cols_13_4_io_left_in_bits),
    .io_top_in_ready(cols_13_4_io_top_in_ready),
    .io_top_in_valid(cols_13_4_io_top_in_valid),
    .io_top_in_bits(cols_13_4_io_top_in_bits),
    .io_sum_ready(cols_13_4_io_sum_ready),
    .io_sum_valid(cols_13_4_io_sum_valid),
    .io_sum_bits(cols_13_4_io_sum_bits),
    .io_right_out_ready(cols_13_4_io_right_out_ready),
    .io_right_out_valid(cols_13_4_io_right_out_valid),
    .io_right_out_bits(cols_13_4_io_right_out_bits),
    .io_bottom_out_ready(cols_13_4_io_bottom_out_ready),
    .io_bottom_out_valid(cols_13_4_io_bottom_out_valid),
    .io_bottom_out_bits(cols_13_4_io_bottom_out_bits)
  );
  ProcessingElement cols_14_4 ( // @[Stab.scala 85:60]
    .clock(cols_14_4_clock),
    .reset(cols_14_4_reset),
    .io_left_in_ready(cols_14_4_io_left_in_ready),
    .io_left_in_valid(cols_14_4_io_left_in_valid),
    .io_left_in_bits(cols_14_4_io_left_in_bits),
    .io_top_in_ready(cols_14_4_io_top_in_ready),
    .io_top_in_valid(cols_14_4_io_top_in_valid),
    .io_top_in_bits(cols_14_4_io_top_in_bits),
    .io_sum_ready(cols_14_4_io_sum_ready),
    .io_sum_valid(cols_14_4_io_sum_valid),
    .io_sum_bits(cols_14_4_io_sum_bits),
    .io_right_out_ready(cols_14_4_io_right_out_ready),
    .io_right_out_valid(cols_14_4_io_right_out_valid),
    .io_right_out_bits(cols_14_4_io_right_out_bits),
    .io_bottom_out_ready(cols_14_4_io_bottom_out_ready),
    .io_bottom_out_valid(cols_14_4_io_bottom_out_valid),
    .io_bottom_out_bits(cols_14_4_io_bottom_out_bits)
  );
  ProcessingElement cols_15_4 ( // @[Stab.scala 85:60]
    .clock(cols_15_4_clock),
    .reset(cols_15_4_reset),
    .io_left_in_ready(cols_15_4_io_left_in_ready),
    .io_left_in_valid(cols_15_4_io_left_in_valid),
    .io_left_in_bits(cols_15_4_io_left_in_bits),
    .io_top_in_ready(cols_15_4_io_top_in_ready),
    .io_top_in_valid(cols_15_4_io_top_in_valid),
    .io_top_in_bits(cols_15_4_io_top_in_bits),
    .io_sum_ready(cols_15_4_io_sum_ready),
    .io_sum_valid(cols_15_4_io_sum_valid),
    .io_sum_bits(cols_15_4_io_sum_bits),
    .io_right_out_ready(cols_15_4_io_right_out_ready),
    .io_right_out_valid(cols_15_4_io_right_out_valid),
    .io_right_out_bits(cols_15_4_io_right_out_bits),
    .io_bottom_out_ready(cols_15_4_io_bottom_out_ready),
    .io_bottom_out_valid(cols_15_4_io_bottom_out_valid),
    .io_bottom_out_bits(cols_15_4_io_bottom_out_bits)
  );
  ProcessingElement cols_0_5 ( // @[Stab.scala 85:60]
    .clock(cols_0_5_clock),
    .reset(cols_0_5_reset),
    .io_left_in_ready(cols_0_5_io_left_in_ready),
    .io_left_in_valid(cols_0_5_io_left_in_valid),
    .io_left_in_bits(cols_0_5_io_left_in_bits),
    .io_top_in_ready(cols_0_5_io_top_in_ready),
    .io_top_in_valid(cols_0_5_io_top_in_valid),
    .io_top_in_bits(cols_0_5_io_top_in_bits),
    .io_sum_ready(cols_0_5_io_sum_ready),
    .io_sum_valid(cols_0_5_io_sum_valid),
    .io_sum_bits(cols_0_5_io_sum_bits),
    .io_right_out_ready(cols_0_5_io_right_out_ready),
    .io_right_out_valid(cols_0_5_io_right_out_valid),
    .io_right_out_bits(cols_0_5_io_right_out_bits),
    .io_bottom_out_ready(cols_0_5_io_bottom_out_ready),
    .io_bottom_out_valid(cols_0_5_io_bottom_out_valid),
    .io_bottom_out_bits(cols_0_5_io_bottom_out_bits)
  );
  ProcessingElement cols_1_5 ( // @[Stab.scala 85:60]
    .clock(cols_1_5_clock),
    .reset(cols_1_5_reset),
    .io_left_in_ready(cols_1_5_io_left_in_ready),
    .io_left_in_valid(cols_1_5_io_left_in_valid),
    .io_left_in_bits(cols_1_5_io_left_in_bits),
    .io_top_in_ready(cols_1_5_io_top_in_ready),
    .io_top_in_valid(cols_1_5_io_top_in_valid),
    .io_top_in_bits(cols_1_5_io_top_in_bits),
    .io_sum_ready(cols_1_5_io_sum_ready),
    .io_sum_valid(cols_1_5_io_sum_valid),
    .io_sum_bits(cols_1_5_io_sum_bits),
    .io_right_out_ready(cols_1_5_io_right_out_ready),
    .io_right_out_valid(cols_1_5_io_right_out_valid),
    .io_right_out_bits(cols_1_5_io_right_out_bits),
    .io_bottom_out_ready(cols_1_5_io_bottom_out_ready),
    .io_bottom_out_valid(cols_1_5_io_bottom_out_valid),
    .io_bottom_out_bits(cols_1_5_io_bottom_out_bits)
  );
  ProcessingElement cols_2_5 ( // @[Stab.scala 85:60]
    .clock(cols_2_5_clock),
    .reset(cols_2_5_reset),
    .io_left_in_ready(cols_2_5_io_left_in_ready),
    .io_left_in_valid(cols_2_5_io_left_in_valid),
    .io_left_in_bits(cols_2_5_io_left_in_bits),
    .io_top_in_ready(cols_2_5_io_top_in_ready),
    .io_top_in_valid(cols_2_5_io_top_in_valid),
    .io_top_in_bits(cols_2_5_io_top_in_bits),
    .io_sum_ready(cols_2_5_io_sum_ready),
    .io_sum_valid(cols_2_5_io_sum_valid),
    .io_sum_bits(cols_2_5_io_sum_bits),
    .io_right_out_ready(cols_2_5_io_right_out_ready),
    .io_right_out_valid(cols_2_5_io_right_out_valid),
    .io_right_out_bits(cols_2_5_io_right_out_bits),
    .io_bottom_out_ready(cols_2_5_io_bottom_out_ready),
    .io_bottom_out_valid(cols_2_5_io_bottom_out_valid),
    .io_bottom_out_bits(cols_2_5_io_bottom_out_bits)
  );
  ProcessingElement cols_3_5 ( // @[Stab.scala 85:60]
    .clock(cols_3_5_clock),
    .reset(cols_3_5_reset),
    .io_left_in_ready(cols_3_5_io_left_in_ready),
    .io_left_in_valid(cols_3_5_io_left_in_valid),
    .io_left_in_bits(cols_3_5_io_left_in_bits),
    .io_top_in_ready(cols_3_5_io_top_in_ready),
    .io_top_in_valid(cols_3_5_io_top_in_valid),
    .io_top_in_bits(cols_3_5_io_top_in_bits),
    .io_sum_ready(cols_3_5_io_sum_ready),
    .io_sum_valid(cols_3_5_io_sum_valid),
    .io_sum_bits(cols_3_5_io_sum_bits),
    .io_right_out_ready(cols_3_5_io_right_out_ready),
    .io_right_out_valid(cols_3_5_io_right_out_valid),
    .io_right_out_bits(cols_3_5_io_right_out_bits),
    .io_bottom_out_ready(cols_3_5_io_bottom_out_ready),
    .io_bottom_out_valid(cols_3_5_io_bottom_out_valid),
    .io_bottom_out_bits(cols_3_5_io_bottom_out_bits)
  );
  ProcessingElement cols_4_5 ( // @[Stab.scala 85:60]
    .clock(cols_4_5_clock),
    .reset(cols_4_5_reset),
    .io_left_in_ready(cols_4_5_io_left_in_ready),
    .io_left_in_valid(cols_4_5_io_left_in_valid),
    .io_left_in_bits(cols_4_5_io_left_in_bits),
    .io_top_in_ready(cols_4_5_io_top_in_ready),
    .io_top_in_valid(cols_4_5_io_top_in_valid),
    .io_top_in_bits(cols_4_5_io_top_in_bits),
    .io_sum_ready(cols_4_5_io_sum_ready),
    .io_sum_valid(cols_4_5_io_sum_valid),
    .io_sum_bits(cols_4_5_io_sum_bits),
    .io_right_out_ready(cols_4_5_io_right_out_ready),
    .io_right_out_valid(cols_4_5_io_right_out_valid),
    .io_right_out_bits(cols_4_5_io_right_out_bits),
    .io_bottom_out_ready(cols_4_5_io_bottom_out_ready),
    .io_bottom_out_valid(cols_4_5_io_bottom_out_valid),
    .io_bottom_out_bits(cols_4_5_io_bottom_out_bits)
  );
  ProcessingElement cols_5_5 ( // @[Stab.scala 85:60]
    .clock(cols_5_5_clock),
    .reset(cols_5_5_reset),
    .io_left_in_ready(cols_5_5_io_left_in_ready),
    .io_left_in_valid(cols_5_5_io_left_in_valid),
    .io_left_in_bits(cols_5_5_io_left_in_bits),
    .io_top_in_ready(cols_5_5_io_top_in_ready),
    .io_top_in_valid(cols_5_5_io_top_in_valid),
    .io_top_in_bits(cols_5_5_io_top_in_bits),
    .io_sum_ready(cols_5_5_io_sum_ready),
    .io_sum_valid(cols_5_5_io_sum_valid),
    .io_sum_bits(cols_5_5_io_sum_bits),
    .io_right_out_ready(cols_5_5_io_right_out_ready),
    .io_right_out_valid(cols_5_5_io_right_out_valid),
    .io_right_out_bits(cols_5_5_io_right_out_bits),
    .io_bottom_out_ready(cols_5_5_io_bottom_out_ready),
    .io_bottom_out_valid(cols_5_5_io_bottom_out_valid),
    .io_bottom_out_bits(cols_5_5_io_bottom_out_bits)
  );
  ProcessingElement cols_6_5 ( // @[Stab.scala 85:60]
    .clock(cols_6_5_clock),
    .reset(cols_6_5_reset),
    .io_left_in_ready(cols_6_5_io_left_in_ready),
    .io_left_in_valid(cols_6_5_io_left_in_valid),
    .io_left_in_bits(cols_6_5_io_left_in_bits),
    .io_top_in_ready(cols_6_5_io_top_in_ready),
    .io_top_in_valid(cols_6_5_io_top_in_valid),
    .io_top_in_bits(cols_6_5_io_top_in_bits),
    .io_sum_ready(cols_6_5_io_sum_ready),
    .io_sum_valid(cols_6_5_io_sum_valid),
    .io_sum_bits(cols_6_5_io_sum_bits),
    .io_right_out_ready(cols_6_5_io_right_out_ready),
    .io_right_out_valid(cols_6_5_io_right_out_valid),
    .io_right_out_bits(cols_6_5_io_right_out_bits),
    .io_bottom_out_ready(cols_6_5_io_bottom_out_ready),
    .io_bottom_out_valid(cols_6_5_io_bottom_out_valid),
    .io_bottom_out_bits(cols_6_5_io_bottom_out_bits)
  );
  ProcessingElement cols_7_5 ( // @[Stab.scala 85:60]
    .clock(cols_7_5_clock),
    .reset(cols_7_5_reset),
    .io_left_in_ready(cols_7_5_io_left_in_ready),
    .io_left_in_valid(cols_7_5_io_left_in_valid),
    .io_left_in_bits(cols_7_5_io_left_in_bits),
    .io_top_in_ready(cols_7_5_io_top_in_ready),
    .io_top_in_valid(cols_7_5_io_top_in_valid),
    .io_top_in_bits(cols_7_5_io_top_in_bits),
    .io_sum_ready(cols_7_5_io_sum_ready),
    .io_sum_valid(cols_7_5_io_sum_valid),
    .io_sum_bits(cols_7_5_io_sum_bits),
    .io_right_out_ready(cols_7_5_io_right_out_ready),
    .io_right_out_valid(cols_7_5_io_right_out_valid),
    .io_right_out_bits(cols_7_5_io_right_out_bits),
    .io_bottom_out_ready(cols_7_5_io_bottom_out_ready),
    .io_bottom_out_valid(cols_7_5_io_bottom_out_valid),
    .io_bottom_out_bits(cols_7_5_io_bottom_out_bits)
  );
  ProcessingElement cols_8_5 ( // @[Stab.scala 85:60]
    .clock(cols_8_5_clock),
    .reset(cols_8_5_reset),
    .io_left_in_ready(cols_8_5_io_left_in_ready),
    .io_left_in_valid(cols_8_5_io_left_in_valid),
    .io_left_in_bits(cols_8_5_io_left_in_bits),
    .io_top_in_ready(cols_8_5_io_top_in_ready),
    .io_top_in_valid(cols_8_5_io_top_in_valid),
    .io_top_in_bits(cols_8_5_io_top_in_bits),
    .io_sum_ready(cols_8_5_io_sum_ready),
    .io_sum_valid(cols_8_5_io_sum_valid),
    .io_sum_bits(cols_8_5_io_sum_bits),
    .io_right_out_ready(cols_8_5_io_right_out_ready),
    .io_right_out_valid(cols_8_5_io_right_out_valid),
    .io_right_out_bits(cols_8_5_io_right_out_bits),
    .io_bottom_out_ready(cols_8_5_io_bottom_out_ready),
    .io_bottom_out_valid(cols_8_5_io_bottom_out_valid),
    .io_bottom_out_bits(cols_8_5_io_bottom_out_bits)
  );
  ProcessingElement cols_9_5 ( // @[Stab.scala 85:60]
    .clock(cols_9_5_clock),
    .reset(cols_9_5_reset),
    .io_left_in_ready(cols_9_5_io_left_in_ready),
    .io_left_in_valid(cols_9_5_io_left_in_valid),
    .io_left_in_bits(cols_9_5_io_left_in_bits),
    .io_top_in_ready(cols_9_5_io_top_in_ready),
    .io_top_in_valid(cols_9_5_io_top_in_valid),
    .io_top_in_bits(cols_9_5_io_top_in_bits),
    .io_sum_ready(cols_9_5_io_sum_ready),
    .io_sum_valid(cols_9_5_io_sum_valid),
    .io_sum_bits(cols_9_5_io_sum_bits),
    .io_right_out_ready(cols_9_5_io_right_out_ready),
    .io_right_out_valid(cols_9_5_io_right_out_valid),
    .io_right_out_bits(cols_9_5_io_right_out_bits),
    .io_bottom_out_ready(cols_9_5_io_bottom_out_ready),
    .io_bottom_out_valid(cols_9_5_io_bottom_out_valid),
    .io_bottom_out_bits(cols_9_5_io_bottom_out_bits)
  );
  ProcessingElement cols_10_5 ( // @[Stab.scala 85:60]
    .clock(cols_10_5_clock),
    .reset(cols_10_5_reset),
    .io_left_in_ready(cols_10_5_io_left_in_ready),
    .io_left_in_valid(cols_10_5_io_left_in_valid),
    .io_left_in_bits(cols_10_5_io_left_in_bits),
    .io_top_in_ready(cols_10_5_io_top_in_ready),
    .io_top_in_valid(cols_10_5_io_top_in_valid),
    .io_top_in_bits(cols_10_5_io_top_in_bits),
    .io_sum_ready(cols_10_5_io_sum_ready),
    .io_sum_valid(cols_10_5_io_sum_valid),
    .io_sum_bits(cols_10_5_io_sum_bits),
    .io_right_out_ready(cols_10_5_io_right_out_ready),
    .io_right_out_valid(cols_10_5_io_right_out_valid),
    .io_right_out_bits(cols_10_5_io_right_out_bits),
    .io_bottom_out_ready(cols_10_5_io_bottom_out_ready),
    .io_bottom_out_valid(cols_10_5_io_bottom_out_valid),
    .io_bottom_out_bits(cols_10_5_io_bottom_out_bits)
  );
  ProcessingElement cols_11_5 ( // @[Stab.scala 85:60]
    .clock(cols_11_5_clock),
    .reset(cols_11_5_reset),
    .io_left_in_ready(cols_11_5_io_left_in_ready),
    .io_left_in_valid(cols_11_5_io_left_in_valid),
    .io_left_in_bits(cols_11_5_io_left_in_bits),
    .io_top_in_ready(cols_11_5_io_top_in_ready),
    .io_top_in_valid(cols_11_5_io_top_in_valid),
    .io_top_in_bits(cols_11_5_io_top_in_bits),
    .io_sum_ready(cols_11_5_io_sum_ready),
    .io_sum_valid(cols_11_5_io_sum_valid),
    .io_sum_bits(cols_11_5_io_sum_bits),
    .io_right_out_ready(cols_11_5_io_right_out_ready),
    .io_right_out_valid(cols_11_5_io_right_out_valid),
    .io_right_out_bits(cols_11_5_io_right_out_bits),
    .io_bottom_out_ready(cols_11_5_io_bottom_out_ready),
    .io_bottom_out_valid(cols_11_5_io_bottom_out_valid),
    .io_bottom_out_bits(cols_11_5_io_bottom_out_bits)
  );
  ProcessingElement cols_12_5 ( // @[Stab.scala 85:60]
    .clock(cols_12_5_clock),
    .reset(cols_12_5_reset),
    .io_left_in_ready(cols_12_5_io_left_in_ready),
    .io_left_in_valid(cols_12_5_io_left_in_valid),
    .io_left_in_bits(cols_12_5_io_left_in_bits),
    .io_top_in_ready(cols_12_5_io_top_in_ready),
    .io_top_in_valid(cols_12_5_io_top_in_valid),
    .io_top_in_bits(cols_12_5_io_top_in_bits),
    .io_sum_ready(cols_12_5_io_sum_ready),
    .io_sum_valid(cols_12_5_io_sum_valid),
    .io_sum_bits(cols_12_5_io_sum_bits),
    .io_right_out_ready(cols_12_5_io_right_out_ready),
    .io_right_out_valid(cols_12_5_io_right_out_valid),
    .io_right_out_bits(cols_12_5_io_right_out_bits),
    .io_bottom_out_ready(cols_12_5_io_bottom_out_ready),
    .io_bottom_out_valid(cols_12_5_io_bottom_out_valid),
    .io_bottom_out_bits(cols_12_5_io_bottom_out_bits)
  );
  ProcessingElement cols_13_5 ( // @[Stab.scala 85:60]
    .clock(cols_13_5_clock),
    .reset(cols_13_5_reset),
    .io_left_in_ready(cols_13_5_io_left_in_ready),
    .io_left_in_valid(cols_13_5_io_left_in_valid),
    .io_left_in_bits(cols_13_5_io_left_in_bits),
    .io_top_in_ready(cols_13_5_io_top_in_ready),
    .io_top_in_valid(cols_13_5_io_top_in_valid),
    .io_top_in_bits(cols_13_5_io_top_in_bits),
    .io_sum_ready(cols_13_5_io_sum_ready),
    .io_sum_valid(cols_13_5_io_sum_valid),
    .io_sum_bits(cols_13_5_io_sum_bits),
    .io_right_out_ready(cols_13_5_io_right_out_ready),
    .io_right_out_valid(cols_13_5_io_right_out_valid),
    .io_right_out_bits(cols_13_5_io_right_out_bits),
    .io_bottom_out_ready(cols_13_5_io_bottom_out_ready),
    .io_bottom_out_valid(cols_13_5_io_bottom_out_valid),
    .io_bottom_out_bits(cols_13_5_io_bottom_out_bits)
  );
  ProcessingElement cols_14_5 ( // @[Stab.scala 85:60]
    .clock(cols_14_5_clock),
    .reset(cols_14_5_reset),
    .io_left_in_ready(cols_14_5_io_left_in_ready),
    .io_left_in_valid(cols_14_5_io_left_in_valid),
    .io_left_in_bits(cols_14_5_io_left_in_bits),
    .io_top_in_ready(cols_14_5_io_top_in_ready),
    .io_top_in_valid(cols_14_5_io_top_in_valid),
    .io_top_in_bits(cols_14_5_io_top_in_bits),
    .io_sum_ready(cols_14_5_io_sum_ready),
    .io_sum_valid(cols_14_5_io_sum_valid),
    .io_sum_bits(cols_14_5_io_sum_bits),
    .io_right_out_ready(cols_14_5_io_right_out_ready),
    .io_right_out_valid(cols_14_5_io_right_out_valid),
    .io_right_out_bits(cols_14_5_io_right_out_bits),
    .io_bottom_out_ready(cols_14_5_io_bottom_out_ready),
    .io_bottom_out_valid(cols_14_5_io_bottom_out_valid),
    .io_bottom_out_bits(cols_14_5_io_bottom_out_bits)
  );
  ProcessingElement cols_15_5 ( // @[Stab.scala 85:60]
    .clock(cols_15_5_clock),
    .reset(cols_15_5_reset),
    .io_left_in_ready(cols_15_5_io_left_in_ready),
    .io_left_in_valid(cols_15_5_io_left_in_valid),
    .io_left_in_bits(cols_15_5_io_left_in_bits),
    .io_top_in_ready(cols_15_5_io_top_in_ready),
    .io_top_in_valid(cols_15_5_io_top_in_valid),
    .io_top_in_bits(cols_15_5_io_top_in_bits),
    .io_sum_ready(cols_15_5_io_sum_ready),
    .io_sum_valid(cols_15_5_io_sum_valid),
    .io_sum_bits(cols_15_5_io_sum_bits),
    .io_right_out_ready(cols_15_5_io_right_out_ready),
    .io_right_out_valid(cols_15_5_io_right_out_valid),
    .io_right_out_bits(cols_15_5_io_right_out_bits),
    .io_bottom_out_ready(cols_15_5_io_bottom_out_ready),
    .io_bottom_out_valid(cols_15_5_io_bottom_out_valid),
    .io_bottom_out_bits(cols_15_5_io_bottom_out_bits)
  );
  ProcessingElement cols_0_6 ( // @[Stab.scala 85:60]
    .clock(cols_0_6_clock),
    .reset(cols_0_6_reset),
    .io_left_in_ready(cols_0_6_io_left_in_ready),
    .io_left_in_valid(cols_0_6_io_left_in_valid),
    .io_left_in_bits(cols_0_6_io_left_in_bits),
    .io_top_in_ready(cols_0_6_io_top_in_ready),
    .io_top_in_valid(cols_0_6_io_top_in_valid),
    .io_top_in_bits(cols_0_6_io_top_in_bits),
    .io_sum_ready(cols_0_6_io_sum_ready),
    .io_sum_valid(cols_0_6_io_sum_valid),
    .io_sum_bits(cols_0_6_io_sum_bits),
    .io_right_out_ready(cols_0_6_io_right_out_ready),
    .io_right_out_valid(cols_0_6_io_right_out_valid),
    .io_right_out_bits(cols_0_6_io_right_out_bits),
    .io_bottom_out_ready(cols_0_6_io_bottom_out_ready),
    .io_bottom_out_valid(cols_0_6_io_bottom_out_valid),
    .io_bottom_out_bits(cols_0_6_io_bottom_out_bits)
  );
  ProcessingElement cols_1_6 ( // @[Stab.scala 85:60]
    .clock(cols_1_6_clock),
    .reset(cols_1_6_reset),
    .io_left_in_ready(cols_1_6_io_left_in_ready),
    .io_left_in_valid(cols_1_6_io_left_in_valid),
    .io_left_in_bits(cols_1_6_io_left_in_bits),
    .io_top_in_ready(cols_1_6_io_top_in_ready),
    .io_top_in_valid(cols_1_6_io_top_in_valid),
    .io_top_in_bits(cols_1_6_io_top_in_bits),
    .io_sum_ready(cols_1_6_io_sum_ready),
    .io_sum_valid(cols_1_6_io_sum_valid),
    .io_sum_bits(cols_1_6_io_sum_bits),
    .io_right_out_ready(cols_1_6_io_right_out_ready),
    .io_right_out_valid(cols_1_6_io_right_out_valid),
    .io_right_out_bits(cols_1_6_io_right_out_bits),
    .io_bottom_out_ready(cols_1_6_io_bottom_out_ready),
    .io_bottom_out_valid(cols_1_6_io_bottom_out_valid),
    .io_bottom_out_bits(cols_1_6_io_bottom_out_bits)
  );
  ProcessingElement cols_2_6 ( // @[Stab.scala 85:60]
    .clock(cols_2_6_clock),
    .reset(cols_2_6_reset),
    .io_left_in_ready(cols_2_6_io_left_in_ready),
    .io_left_in_valid(cols_2_6_io_left_in_valid),
    .io_left_in_bits(cols_2_6_io_left_in_bits),
    .io_top_in_ready(cols_2_6_io_top_in_ready),
    .io_top_in_valid(cols_2_6_io_top_in_valid),
    .io_top_in_bits(cols_2_6_io_top_in_bits),
    .io_sum_ready(cols_2_6_io_sum_ready),
    .io_sum_valid(cols_2_6_io_sum_valid),
    .io_sum_bits(cols_2_6_io_sum_bits),
    .io_right_out_ready(cols_2_6_io_right_out_ready),
    .io_right_out_valid(cols_2_6_io_right_out_valid),
    .io_right_out_bits(cols_2_6_io_right_out_bits),
    .io_bottom_out_ready(cols_2_6_io_bottom_out_ready),
    .io_bottom_out_valid(cols_2_6_io_bottom_out_valid),
    .io_bottom_out_bits(cols_2_6_io_bottom_out_bits)
  );
  ProcessingElement cols_3_6 ( // @[Stab.scala 85:60]
    .clock(cols_3_6_clock),
    .reset(cols_3_6_reset),
    .io_left_in_ready(cols_3_6_io_left_in_ready),
    .io_left_in_valid(cols_3_6_io_left_in_valid),
    .io_left_in_bits(cols_3_6_io_left_in_bits),
    .io_top_in_ready(cols_3_6_io_top_in_ready),
    .io_top_in_valid(cols_3_6_io_top_in_valid),
    .io_top_in_bits(cols_3_6_io_top_in_bits),
    .io_sum_ready(cols_3_6_io_sum_ready),
    .io_sum_valid(cols_3_6_io_sum_valid),
    .io_sum_bits(cols_3_6_io_sum_bits),
    .io_right_out_ready(cols_3_6_io_right_out_ready),
    .io_right_out_valid(cols_3_6_io_right_out_valid),
    .io_right_out_bits(cols_3_6_io_right_out_bits),
    .io_bottom_out_ready(cols_3_6_io_bottom_out_ready),
    .io_bottom_out_valid(cols_3_6_io_bottom_out_valid),
    .io_bottom_out_bits(cols_3_6_io_bottom_out_bits)
  );
  ProcessingElement cols_4_6 ( // @[Stab.scala 85:60]
    .clock(cols_4_6_clock),
    .reset(cols_4_6_reset),
    .io_left_in_ready(cols_4_6_io_left_in_ready),
    .io_left_in_valid(cols_4_6_io_left_in_valid),
    .io_left_in_bits(cols_4_6_io_left_in_bits),
    .io_top_in_ready(cols_4_6_io_top_in_ready),
    .io_top_in_valid(cols_4_6_io_top_in_valid),
    .io_top_in_bits(cols_4_6_io_top_in_bits),
    .io_sum_ready(cols_4_6_io_sum_ready),
    .io_sum_valid(cols_4_6_io_sum_valid),
    .io_sum_bits(cols_4_6_io_sum_bits),
    .io_right_out_ready(cols_4_6_io_right_out_ready),
    .io_right_out_valid(cols_4_6_io_right_out_valid),
    .io_right_out_bits(cols_4_6_io_right_out_bits),
    .io_bottom_out_ready(cols_4_6_io_bottom_out_ready),
    .io_bottom_out_valid(cols_4_6_io_bottom_out_valid),
    .io_bottom_out_bits(cols_4_6_io_bottom_out_bits)
  );
  ProcessingElement cols_5_6 ( // @[Stab.scala 85:60]
    .clock(cols_5_6_clock),
    .reset(cols_5_6_reset),
    .io_left_in_ready(cols_5_6_io_left_in_ready),
    .io_left_in_valid(cols_5_6_io_left_in_valid),
    .io_left_in_bits(cols_5_6_io_left_in_bits),
    .io_top_in_ready(cols_5_6_io_top_in_ready),
    .io_top_in_valid(cols_5_6_io_top_in_valid),
    .io_top_in_bits(cols_5_6_io_top_in_bits),
    .io_sum_ready(cols_5_6_io_sum_ready),
    .io_sum_valid(cols_5_6_io_sum_valid),
    .io_sum_bits(cols_5_6_io_sum_bits),
    .io_right_out_ready(cols_5_6_io_right_out_ready),
    .io_right_out_valid(cols_5_6_io_right_out_valid),
    .io_right_out_bits(cols_5_6_io_right_out_bits),
    .io_bottom_out_ready(cols_5_6_io_bottom_out_ready),
    .io_bottom_out_valid(cols_5_6_io_bottom_out_valid),
    .io_bottom_out_bits(cols_5_6_io_bottom_out_bits)
  );
  ProcessingElement cols_6_6 ( // @[Stab.scala 85:60]
    .clock(cols_6_6_clock),
    .reset(cols_6_6_reset),
    .io_left_in_ready(cols_6_6_io_left_in_ready),
    .io_left_in_valid(cols_6_6_io_left_in_valid),
    .io_left_in_bits(cols_6_6_io_left_in_bits),
    .io_top_in_ready(cols_6_6_io_top_in_ready),
    .io_top_in_valid(cols_6_6_io_top_in_valid),
    .io_top_in_bits(cols_6_6_io_top_in_bits),
    .io_sum_ready(cols_6_6_io_sum_ready),
    .io_sum_valid(cols_6_6_io_sum_valid),
    .io_sum_bits(cols_6_6_io_sum_bits),
    .io_right_out_ready(cols_6_6_io_right_out_ready),
    .io_right_out_valid(cols_6_6_io_right_out_valid),
    .io_right_out_bits(cols_6_6_io_right_out_bits),
    .io_bottom_out_ready(cols_6_6_io_bottom_out_ready),
    .io_bottom_out_valid(cols_6_6_io_bottom_out_valid),
    .io_bottom_out_bits(cols_6_6_io_bottom_out_bits)
  );
  ProcessingElement cols_7_6 ( // @[Stab.scala 85:60]
    .clock(cols_7_6_clock),
    .reset(cols_7_6_reset),
    .io_left_in_ready(cols_7_6_io_left_in_ready),
    .io_left_in_valid(cols_7_6_io_left_in_valid),
    .io_left_in_bits(cols_7_6_io_left_in_bits),
    .io_top_in_ready(cols_7_6_io_top_in_ready),
    .io_top_in_valid(cols_7_6_io_top_in_valid),
    .io_top_in_bits(cols_7_6_io_top_in_bits),
    .io_sum_ready(cols_7_6_io_sum_ready),
    .io_sum_valid(cols_7_6_io_sum_valid),
    .io_sum_bits(cols_7_6_io_sum_bits),
    .io_right_out_ready(cols_7_6_io_right_out_ready),
    .io_right_out_valid(cols_7_6_io_right_out_valid),
    .io_right_out_bits(cols_7_6_io_right_out_bits),
    .io_bottom_out_ready(cols_7_6_io_bottom_out_ready),
    .io_bottom_out_valid(cols_7_6_io_bottom_out_valid),
    .io_bottom_out_bits(cols_7_6_io_bottom_out_bits)
  );
  ProcessingElement cols_8_6 ( // @[Stab.scala 85:60]
    .clock(cols_8_6_clock),
    .reset(cols_8_6_reset),
    .io_left_in_ready(cols_8_6_io_left_in_ready),
    .io_left_in_valid(cols_8_6_io_left_in_valid),
    .io_left_in_bits(cols_8_6_io_left_in_bits),
    .io_top_in_ready(cols_8_6_io_top_in_ready),
    .io_top_in_valid(cols_8_6_io_top_in_valid),
    .io_top_in_bits(cols_8_6_io_top_in_bits),
    .io_sum_ready(cols_8_6_io_sum_ready),
    .io_sum_valid(cols_8_6_io_sum_valid),
    .io_sum_bits(cols_8_6_io_sum_bits),
    .io_right_out_ready(cols_8_6_io_right_out_ready),
    .io_right_out_valid(cols_8_6_io_right_out_valid),
    .io_right_out_bits(cols_8_6_io_right_out_bits),
    .io_bottom_out_ready(cols_8_6_io_bottom_out_ready),
    .io_bottom_out_valid(cols_8_6_io_bottom_out_valid),
    .io_bottom_out_bits(cols_8_6_io_bottom_out_bits)
  );
  ProcessingElement cols_9_6 ( // @[Stab.scala 85:60]
    .clock(cols_9_6_clock),
    .reset(cols_9_6_reset),
    .io_left_in_ready(cols_9_6_io_left_in_ready),
    .io_left_in_valid(cols_9_6_io_left_in_valid),
    .io_left_in_bits(cols_9_6_io_left_in_bits),
    .io_top_in_ready(cols_9_6_io_top_in_ready),
    .io_top_in_valid(cols_9_6_io_top_in_valid),
    .io_top_in_bits(cols_9_6_io_top_in_bits),
    .io_sum_ready(cols_9_6_io_sum_ready),
    .io_sum_valid(cols_9_6_io_sum_valid),
    .io_sum_bits(cols_9_6_io_sum_bits),
    .io_right_out_ready(cols_9_6_io_right_out_ready),
    .io_right_out_valid(cols_9_6_io_right_out_valid),
    .io_right_out_bits(cols_9_6_io_right_out_bits),
    .io_bottom_out_ready(cols_9_6_io_bottom_out_ready),
    .io_bottom_out_valid(cols_9_6_io_bottom_out_valid),
    .io_bottom_out_bits(cols_9_6_io_bottom_out_bits)
  );
  ProcessingElement cols_10_6 ( // @[Stab.scala 85:60]
    .clock(cols_10_6_clock),
    .reset(cols_10_6_reset),
    .io_left_in_ready(cols_10_6_io_left_in_ready),
    .io_left_in_valid(cols_10_6_io_left_in_valid),
    .io_left_in_bits(cols_10_6_io_left_in_bits),
    .io_top_in_ready(cols_10_6_io_top_in_ready),
    .io_top_in_valid(cols_10_6_io_top_in_valid),
    .io_top_in_bits(cols_10_6_io_top_in_bits),
    .io_sum_ready(cols_10_6_io_sum_ready),
    .io_sum_valid(cols_10_6_io_sum_valid),
    .io_sum_bits(cols_10_6_io_sum_bits),
    .io_right_out_ready(cols_10_6_io_right_out_ready),
    .io_right_out_valid(cols_10_6_io_right_out_valid),
    .io_right_out_bits(cols_10_6_io_right_out_bits),
    .io_bottom_out_ready(cols_10_6_io_bottom_out_ready),
    .io_bottom_out_valid(cols_10_6_io_bottom_out_valid),
    .io_bottom_out_bits(cols_10_6_io_bottom_out_bits)
  );
  ProcessingElement cols_11_6 ( // @[Stab.scala 85:60]
    .clock(cols_11_6_clock),
    .reset(cols_11_6_reset),
    .io_left_in_ready(cols_11_6_io_left_in_ready),
    .io_left_in_valid(cols_11_6_io_left_in_valid),
    .io_left_in_bits(cols_11_6_io_left_in_bits),
    .io_top_in_ready(cols_11_6_io_top_in_ready),
    .io_top_in_valid(cols_11_6_io_top_in_valid),
    .io_top_in_bits(cols_11_6_io_top_in_bits),
    .io_sum_ready(cols_11_6_io_sum_ready),
    .io_sum_valid(cols_11_6_io_sum_valid),
    .io_sum_bits(cols_11_6_io_sum_bits),
    .io_right_out_ready(cols_11_6_io_right_out_ready),
    .io_right_out_valid(cols_11_6_io_right_out_valid),
    .io_right_out_bits(cols_11_6_io_right_out_bits),
    .io_bottom_out_ready(cols_11_6_io_bottom_out_ready),
    .io_bottom_out_valid(cols_11_6_io_bottom_out_valid),
    .io_bottom_out_bits(cols_11_6_io_bottom_out_bits)
  );
  ProcessingElement cols_12_6 ( // @[Stab.scala 85:60]
    .clock(cols_12_6_clock),
    .reset(cols_12_6_reset),
    .io_left_in_ready(cols_12_6_io_left_in_ready),
    .io_left_in_valid(cols_12_6_io_left_in_valid),
    .io_left_in_bits(cols_12_6_io_left_in_bits),
    .io_top_in_ready(cols_12_6_io_top_in_ready),
    .io_top_in_valid(cols_12_6_io_top_in_valid),
    .io_top_in_bits(cols_12_6_io_top_in_bits),
    .io_sum_ready(cols_12_6_io_sum_ready),
    .io_sum_valid(cols_12_6_io_sum_valid),
    .io_sum_bits(cols_12_6_io_sum_bits),
    .io_right_out_ready(cols_12_6_io_right_out_ready),
    .io_right_out_valid(cols_12_6_io_right_out_valid),
    .io_right_out_bits(cols_12_6_io_right_out_bits),
    .io_bottom_out_ready(cols_12_6_io_bottom_out_ready),
    .io_bottom_out_valid(cols_12_6_io_bottom_out_valid),
    .io_bottom_out_bits(cols_12_6_io_bottom_out_bits)
  );
  ProcessingElement cols_13_6 ( // @[Stab.scala 85:60]
    .clock(cols_13_6_clock),
    .reset(cols_13_6_reset),
    .io_left_in_ready(cols_13_6_io_left_in_ready),
    .io_left_in_valid(cols_13_6_io_left_in_valid),
    .io_left_in_bits(cols_13_6_io_left_in_bits),
    .io_top_in_ready(cols_13_6_io_top_in_ready),
    .io_top_in_valid(cols_13_6_io_top_in_valid),
    .io_top_in_bits(cols_13_6_io_top_in_bits),
    .io_sum_ready(cols_13_6_io_sum_ready),
    .io_sum_valid(cols_13_6_io_sum_valid),
    .io_sum_bits(cols_13_6_io_sum_bits),
    .io_right_out_ready(cols_13_6_io_right_out_ready),
    .io_right_out_valid(cols_13_6_io_right_out_valid),
    .io_right_out_bits(cols_13_6_io_right_out_bits),
    .io_bottom_out_ready(cols_13_6_io_bottom_out_ready),
    .io_bottom_out_valid(cols_13_6_io_bottom_out_valid),
    .io_bottom_out_bits(cols_13_6_io_bottom_out_bits)
  );
  ProcessingElement cols_14_6 ( // @[Stab.scala 85:60]
    .clock(cols_14_6_clock),
    .reset(cols_14_6_reset),
    .io_left_in_ready(cols_14_6_io_left_in_ready),
    .io_left_in_valid(cols_14_6_io_left_in_valid),
    .io_left_in_bits(cols_14_6_io_left_in_bits),
    .io_top_in_ready(cols_14_6_io_top_in_ready),
    .io_top_in_valid(cols_14_6_io_top_in_valid),
    .io_top_in_bits(cols_14_6_io_top_in_bits),
    .io_sum_ready(cols_14_6_io_sum_ready),
    .io_sum_valid(cols_14_6_io_sum_valid),
    .io_sum_bits(cols_14_6_io_sum_bits),
    .io_right_out_ready(cols_14_6_io_right_out_ready),
    .io_right_out_valid(cols_14_6_io_right_out_valid),
    .io_right_out_bits(cols_14_6_io_right_out_bits),
    .io_bottom_out_ready(cols_14_6_io_bottom_out_ready),
    .io_bottom_out_valid(cols_14_6_io_bottom_out_valid),
    .io_bottom_out_bits(cols_14_6_io_bottom_out_bits)
  );
  ProcessingElement cols_15_6 ( // @[Stab.scala 85:60]
    .clock(cols_15_6_clock),
    .reset(cols_15_6_reset),
    .io_left_in_ready(cols_15_6_io_left_in_ready),
    .io_left_in_valid(cols_15_6_io_left_in_valid),
    .io_left_in_bits(cols_15_6_io_left_in_bits),
    .io_top_in_ready(cols_15_6_io_top_in_ready),
    .io_top_in_valid(cols_15_6_io_top_in_valid),
    .io_top_in_bits(cols_15_6_io_top_in_bits),
    .io_sum_ready(cols_15_6_io_sum_ready),
    .io_sum_valid(cols_15_6_io_sum_valid),
    .io_sum_bits(cols_15_6_io_sum_bits),
    .io_right_out_ready(cols_15_6_io_right_out_ready),
    .io_right_out_valid(cols_15_6_io_right_out_valid),
    .io_right_out_bits(cols_15_6_io_right_out_bits),
    .io_bottom_out_ready(cols_15_6_io_bottom_out_ready),
    .io_bottom_out_valid(cols_15_6_io_bottom_out_valid),
    .io_bottom_out_bits(cols_15_6_io_bottom_out_bits)
  );
  ProcessingElement cols_0_7 ( // @[Stab.scala 85:60]
    .clock(cols_0_7_clock),
    .reset(cols_0_7_reset),
    .io_left_in_ready(cols_0_7_io_left_in_ready),
    .io_left_in_valid(cols_0_7_io_left_in_valid),
    .io_left_in_bits(cols_0_7_io_left_in_bits),
    .io_top_in_ready(cols_0_7_io_top_in_ready),
    .io_top_in_valid(cols_0_7_io_top_in_valid),
    .io_top_in_bits(cols_0_7_io_top_in_bits),
    .io_sum_ready(cols_0_7_io_sum_ready),
    .io_sum_valid(cols_0_7_io_sum_valid),
    .io_sum_bits(cols_0_7_io_sum_bits),
    .io_right_out_ready(cols_0_7_io_right_out_ready),
    .io_right_out_valid(cols_0_7_io_right_out_valid),
    .io_right_out_bits(cols_0_7_io_right_out_bits),
    .io_bottom_out_ready(cols_0_7_io_bottom_out_ready),
    .io_bottom_out_valid(cols_0_7_io_bottom_out_valid),
    .io_bottom_out_bits(cols_0_7_io_bottom_out_bits)
  );
  ProcessingElement cols_1_7 ( // @[Stab.scala 85:60]
    .clock(cols_1_7_clock),
    .reset(cols_1_7_reset),
    .io_left_in_ready(cols_1_7_io_left_in_ready),
    .io_left_in_valid(cols_1_7_io_left_in_valid),
    .io_left_in_bits(cols_1_7_io_left_in_bits),
    .io_top_in_ready(cols_1_7_io_top_in_ready),
    .io_top_in_valid(cols_1_7_io_top_in_valid),
    .io_top_in_bits(cols_1_7_io_top_in_bits),
    .io_sum_ready(cols_1_7_io_sum_ready),
    .io_sum_valid(cols_1_7_io_sum_valid),
    .io_sum_bits(cols_1_7_io_sum_bits),
    .io_right_out_ready(cols_1_7_io_right_out_ready),
    .io_right_out_valid(cols_1_7_io_right_out_valid),
    .io_right_out_bits(cols_1_7_io_right_out_bits),
    .io_bottom_out_ready(cols_1_7_io_bottom_out_ready),
    .io_bottom_out_valid(cols_1_7_io_bottom_out_valid),
    .io_bottom_out_bits(cols_1_7_io_bottom_out_bits)
  );
  ProcessingElement cols_2_7 ( // @[Stab.scala 85:60]
    .clock(cols_2_7_clock),
    .reset(cols_2_7_reset),
    .io_left_in_ready(cols_2_7_io_left_in_ready),
    .io_left_in_valid(cols_2_7_io_left_in_valid),
    .io_left_in_bits(cols_2_7_io_left_in_bits),
    .io_top_in_ready(cols_2_7_io_top_in_ready),
    .io_top_in_valid(cols_2_7_io_top_in_valid),
    .io_top_in_bits(cols_2_7_io_top_in_bits),
    .io_sum_ready(cols_2_7_io_sum_ready),
    .io_sum_valid(cols_2_7_io_sum_valid),
    .io_sum_bits(cols_2_7_io_sum_bits),
    .io_right_out_ready(cols_2_7_io_right_out_ready),
    .io_right_out_valid(cols_2_7_io_right_out_valid),
    .io_right_out_bits(cols_2_7_io_right_out_bits),
    .io_bottom_out_ready(cols_2_7_io_bottom_out_ready),
    .io_bottom_out_valid(cols_2_7_io_bottom_out_valid),
    .io_bottom_out_bits(cols_2_7_io_bottom_out_bits)
  );
  ProcessingElement cols_3_7 ( // @[Stab.scala 85:60]
    .clock(cols_3_7_clock),
    .reset(cols_3_7_reset),
    .io_left_in_ready(cols_3_7_io_left_in_ready),
    .io_left_in_valid(cols_3_7_io_left_in_valid),
    .io_left_in_bits(cols_3_7_io_left_in_bits),
    .io_top_in_ready(cols_3_7_io_top_in_ready),
    .io_top_in_valid(cols_3_7_io_top_in_valid),
    .io_top_in_bits(cols_3_7_io_top_in_bits),
    .io_sum_ready(cols_3_7_io_sum_ready),
    .io_sum_valid(cols_3_7_io_sum_valid),
    .io_sum_bits(cols_3_7_io_sum_bits),
    .io_right_out_ready(cols_3_7_io_right_out_ready),
    .io_right_out_valid(cols_3_7_io_right_out_valid),
    .io_right_out_bits(cols_3_7_io_right_out_bits),
    .io_bottom_out_ready(cols_3_7_io_bottom_out_ready),
    .io_bottom_out_valid(cols_3_7_io_bottom_out_valid),
    .io_bottom_out_bits(cols_3_7_io_bottom_out_bits)
  );
  ProcessingElement cols_4_7 ( // @[Stab.scala 85:60]
    .clock(cols_4_7_clock),
    .reset(cols_4_7_reset),
    .io_left_in_ready(cols_4_7_io_left_in_ready),
    .io_left_in_valid(cols_4_7_io_left_in_valid),
    .io_left_in_bits(cols_4_7_io_left_in_bits),
    .io_top_in_ready(cols_4_7_io_top_in_ready),
    .io_top_in_valid(cols_4_7_io_top_in_valid),
    .io_top_in_bits(cols_4_7_io_top_in_bits),
    .io_sum_ready(cols_4_7_io_sum_ready),
    .io_sum_valid(cols_4_7_io_sum_valid),
    .io_sum_bits(cols_4_7_io_sum_bits),
    .io_right_out_ready(cols_4_7_io_right_out_ready),
    .io_right_out_valid(cols_4_7_io_right_out_valid),
    .io_right_out_bits(cols_4_7_io_right_out_bits),
    .io_bottom_out_ready(cols_4_7_io_bottom_out_ready),
    .io_bottom_out_valid(cols_4_7_io_bottom_out_valid),
    .io_bottom_out_bits(cols_4_7_io_bottom_out_bits)
  );
  ProcessingElement cols_5_7 ( // @[Stab.scala 85:60]
    .clock(cols_5_7_clock),
    .reset(cols_5_7_reset),
    .io_left_in_ready(cols_5_7_io_left_in_ready),
    .io_left_in_valid(cols_5_7_io_left_in_valid),
    .io_left_in_bits(cols_5_7_io_left_in_bits),
    .io_top_in_ready(cols_5_7_io_top_in_ready),
    .io_top_in_valid(cols_5_7_io_top_in_valid),
    .io_top_in_bits(cols_5_7_io_top_in_bits),
    .io_sum_ready(cols_5_7_io_sum_ready),
    .io_sum_valid(cols_5_7_io_sum_valid),
    .io_sum_bits(cols_5_7_io_sum_bits),
    .io_right_out_ready(cols_5_7_io_right_out_ready),
    .io_right_out_valid(cols_5_7_io_right_out_valid),
    .io_right_out_bits(cols_5_7_io_right_out_bits),
    .io_bottom_out_ready(cols_5_7_io_bottom_out_ready),
    .io_bottom_out_valid(cols_5_7_io_bottom_out_valid),
    .io_bottom_out_bits(cols_5_7_io_bottom_out_bits)
  );
  ProcessingElement cols_6_7 ( // @[Stab.scala 85:60]
    .clock(cols_6_7_clock),
    .reset(cols_6_7_reset),
    .io_left_in_ready(cols_6_7_io_left_in_ready),
    .io_left_in_valid(cols_6_7_io_left_in_valid),
    .io_left_in_bits(cols_6_7_io_left_in_bits),
    .io_top_in_ready(cols_6_7_io_top_in_ready),
    .io_top_in_valid(cols_6_7_io_top_in_valid),
    .io_top_in_bits(cols_6_7_io_top_in_bits),
    .io_sum_ready(cols_6_7_io_sum_ready),
    .io_sum_valid(cols_6_7_io_sum_valid),
    .io_sum_bits(cols_6_7_io_sum_bits),
    .io_right_out_ready(cols_6_7_io_right_out_ready),
    .io_right_out_valid(cols_6_7_io_right_out_valid),
    .io_right_out_bits(cols_6_7_io_right_out_bits),
    .io_bottom_out_ready(cols_6_7_io_bottom_out_ready),
    .io_bottom_out_valid(cols_6_7_io_bottom_out_valid),
    .io_bottom_out_bits(cols_6_7_io_bottom_out_bits)
  );
  ProcessingElement cols_7_7 ( // @[Stab.scala 85:60]
    .clock(cols_7_7_clock),
    .reset(cols_7_7_reset),
    .io_left_in_ready(cols_7_7_io_left_in_ready),
    .io_left_in_valid(cols_7_7_io_left_in_valid),
    .io_left_in_bits(cols_7_7_io_left_in_bits),
    .io_top_in_ready(cols_7_7_io_top_in_ready),
    .io_top_in_valid(cols_7_7_io_top_in_valid),
    .io_top_in_bits(cols_7_7_io_top_in_bits),
    .io_sum_ready(cols_7_7_io_sum_ready),
    .io_sum_valid(cols_7_7_io_sum_valid),
    .io_sum_bits(cols_7_7_io_sum_bits),
    .io_right_out_ready(cols_7_7_io_right_out_ready),
    .io_right_out_valid(cols_7_7_io_right_out_valid),
    .io_right_out_bits(cols_7_7_io_right_out_bits),
    .io_bottom_out_ready(cols_7_7_io_bottom_out_ready),
    .io_bottom_out_valid(cols_7_7_io_bottom_out_valid),
    .io_bottom_out_bits(cols_7_7_io_bottom_out_bits)
  );
  ProcessingElement cols_8_7 ( // @[Stab.scala 85:60]
    .clock(cols_8_7_clock),
    .reset(cols_8_7_reset),
    .io_left_in_ready(cols_8_7_io_left_in_ready),
    .io_left_in_valid(cols_8_7_io_left_in_valid),
    .io_left_in_bits(cols_8_7_io_left_in_bits),
    .io_top_in_ready(cols_8_7_io_top_in_ready),
    .io_top_in_valid(cols_8_7_io_top_in_valid),
    .io_top_in_bits(cols_8_7_io_top_in_bits),
    .io_sum_ready(cols_8_7_io_sum_ready),
    .io_sum_valid(cols_8_7_io_sum_valid),
    .io_sum_bits(cols_8_7_io_sum_bits),
    .io_right_out_ready(cols_8_7_io_right_out_ready),
    .io_right_out_valid(cols_8_7_io_right_out_valid),
    .io_right_out_bits(cols_8_7_io_right_out_bits),
    .io_bottom_out_ready(cols_8_7_io_bottom_out_ready),
    .io_bottom_out_valid(cols_8_7_io_bottom_out_valid),
    .io_bottom_out_bits(cols_8_7_io_bottom_out_bits)
  );
  ProcessingElement cols_9_7 ( // @[Stab.scala 85:60]
    .clock(cols_9_7_clock),
    .reset(cols_9_7_reset),
    .io_left_in_ready(cols_9_7_io_left_in_ready),
    .io_left_in_valid(cols_9_7_io_left_in_valid),
    .io_left_in_bits(cols_9_7_io_left_in_bits),
    .io_top_in_ready(cols_9_7_io_top_in_ready),
    .io_top_in_valid(cols_9_7_io_top_in_valid),
    .io_top_in_bits(cols_9_7_io_top_in_bits),
    .io_sum_ready(cols_9_7_io_sum_ready),
    .io_sum_valid(cols_9_7_io_sum_valid),
    .io_sum_bits(cols_9_7_io_sum_bits),
    .io_right_out_ready(cols_9_7_io_right_out_ready),
    .io_right_out_valid(cols_9_7_io_right_out_valid),
    .io_right_out_bits(cols_9_7_io_right_out_bits),
    .io_bottom_out_ready(cols_9_7_io_bottom_out_ready),
    .io_bottom_out_valid(cols_9_7_io_bottom_out_valid),
    .io_bottom_out_bits(cols_9_7_io_bottom_out_bits)
  );
  ProcessingElement cols_10_7 ( // @[Stab.scala 85:60]
    .clock(cols_10_7_clock),
    .reset(cols_10_7_reset),
    .io_left_in_ready(cols_10_7_io_left_in_ready),
    .io_left_in_valid(cols_10_7_io_left_in_valid),
    .io_left_in_bits(cols_10_7_io_left_in_bits),
    .io_top_in_ready(cols_10_7_io_top_in_ready),
    .io_top_in_valid(cols_10_7_io_top_in_valid),
    .io_top_in_bits(cols_10_7_io_top_in_bits),
    .io_sum_ready(cols_10_7_io_sum_ready),
    .io_sum_valid(cols_10_7_io_sum_valid),
    .io_sum_bits(cols_10_7_io_sum_bits),
    .io_right_out_ready(cols_10_7_io_right_out_ready),
    .io_right_out_valid(cols_10_7_io_right_out_valid),
    .io_right_out_bits(cols_10_7_io_right_out_bits),
    .io_bottom_out_ready(cols_10_7_io_bottom_out_ready),
    .io_bottom_out_valid(cols_10_7_io_bottom_out_valid),
    .io_bottom_out_bits(cols_10_7_io_bottom_out_bits)
  );
  ProcessingElement cols_11_7 ( // @[Stab.scala 85:60]
    .clock(cols_11_7_clock),
    .reset(cols_11_7_reset),
    .io_left_in_ready(cols_11_7_io_left_in_ready),
    .io_left_in_valid(cols_11_7_io_left_in_valid),
    .io_left_in_bits(cols_11_7_io_left_in_bits),
    .io_top_in_ready(cols_11_7_io_top_in_ready),
    .io_top_in_valid(cols_11_7_io_top_in_valid),
    .io_top_in_bits(cols_11_7_io_top_in_bits),
    .io_sum_ready(cols_11_7_io_sum_ready),
    .io_sum_valid(cols_11_7_io_sum_valid),
    .io_sum_bits(cols_11_7_io_sum_bits),
    .io_right_out_ready(cols_11_7_io_right_out_ready),
    .io_right_out_valid(cols_11_7_io_right_out_valid),
    .io_right_out_bits(cols_11_7_io_right_out_bits),
    .io_bottom_out_ready(cols_11_7_io_bottom_out_ready),
    .io_bottom_out_valid(cols_11_7_io_bottom_out_valid),
    .io_bottom_out_bits(cols_11_7_io_bottom_out_bits)
  );
  ProcessingElement cols_12_7 ( // @[Stab.scala 85:60]
    .clock(cols_12_7_clock),
    .reset(cols_12_7_reset),
    .io_left_in_ready(cols_12_7_io_left_in_ready),
    .io_left_in_valid(cols_12_7_io_left_in_valid),
    .io_left_in_bits(cols_12_7_io_left_in_bits),
    .io_top_in_ready(cols_12_7_io_top_in_ready),
    .io_top_in_valid(cols_12_7_io_top_in_valid),
    .io_top_in_bits(cols_12_7_io_top_in_bits),
    .io_sum_ready(cols_12_7_io_sum_ready),
    .io_sum_valid(cols_12_7_io_sum_valid),
    .io_sum_bits(cols_12_7_io_sum_bits),
    .io_right_out_ready(cols_12_7_io_right_out_ready),
    .io_right_out_valid(cols_12_7_io_right_out_valid),
    .io_right_out_bits(cols_12_7_io_right_out_bits),
    .io_bottom_out_ready(cols_12_7_io_bottom_out_ready),
    .io_bottom_out_valid(cols_12_7_io_bottom_out_valid),
    .io_bottom_out_bits(cols_12_7_io_bottom_out_bits)
  );
  ProcessingElement cols_13_7 ( // @[Stab.scala 85:60]
    .clock(cols_13_7_clock),
    .reset(cols_13_7_reset),
    .io_left_in_ready(cols_13_7_io_left_in_ready),
    .io_left_in_valid(cols_13_7_io_left_in_valid),
    .io_left_in_bits(cols_13_7_io_left_in_bits),
    .io_top_in_ready(cols_13_7_io_top_in_ready),
    .io_top_in_valid(cols_13_7_io_top_in_valid),
    .io_top_in_bits(cols_13_7_io_top_in_bits),
    .io_sum_ready(cols_13_7_io_sum_ready),
    .io_sum_valid(cols_13_7_io_sum_valid),
    .io_sum_bits(cols_13_7_io_sum_bits),
    .io_right_out_ready(cols_13_7_io_right_out_ready),
    .io_right_out_valid(cols_13_7_io_right_out_valid),
    .io_right_out_bits(cols_13_7_io_right_out_bits),
    .io_bottom_out_ready(cols_13_7_io_bottom_out_ready),
    .io_bottom_out_valid(cols_13_7_io_bottom_out_valid),
    .io_bottom_out_bits(cols_13_7_io_bottom_out_bits)
  );
  ProcessingElement cols_14_7 ( // @[Stab.scala 85:60]
    .clock(cols_14_7_clock),
    .reset(cols_14_7_reset),
    .io_left_in_ready(cols_14_7_io_left_in_ready),
    .io_left_in_valid(cols_14_7_io_left_in_valid),
    .io_left_in_bits(cols_14_7_io_left_in_bits),
    .io_top_in_ready(cols_14_7_io_top_in_ready),
    .io_top_in_valid(cols_14_7_io_top_in_valid),
    .io_top_in_bits(cols_14_7_io_top_in_bits),
    .io_sum_ready(cols_14_7_io_sum_ready),
    .io_sum_valid(cols_14_7_io_sum_valid),
    .io_sum_bits(cols_14_7_io_sum_bits),
    .io_right_out_ready(cols_14_7_io_right_out_ready),
    .io_right_out_valid(cols_14_7_io_right_out_valid),
    .io_right_out_bits(cols_14_7_io_right_out_bits),
    .io_bottom_out_ready(cols_14_7_io_bottom_out_ready),
    .io_bottom_out_valid(cols_14_7_io_bottom_out_valid),
    .io_bottom_out_bits(cols_14_7_io_bottom_out_bits)
  );
  ProcessingElement cols_15_7 ( // @[Stab.scala 85:60]
    .clock(cols_15_7_clock),
    .reset(cols_15_7_reset),
    .io_left_in_ready(cols_15_7_io_left_in_ready),
    .io_left_in_valid(cols_15_7_io_left_in_valid),
    .io_left_in_bits(cols_15_7_io_left_in_bits),
    .io_top_in_ready(cols_15_7_io_top_in_ready),
    .io_top_in_valid(cols_15_7_io_top_in_valid),
    .io_top_in_bits(cols_15_7_io_top_in_bits),
    .io_sum_ready(cols_15_7_io_sum_ready),
    .io_sum_valid(cols_15_7_io_sum_valid),
    .io_sum_bits(cols_15_7_io_sum_bits),
    .io_right_out_ready(cols_15_7_io_right_out_ready),
    .io_right_out_valid(cols_15_7_io_right_out_valid),
    .io_right_out_bits(cols_15_7_io_right_out_bits),
    .io_bottom_out_ready(cols_15_7_io_bottom_out_ready),
    .io_bottom_out_valid(cols_15_7_io_bottom_out_valid),
    .io_bottom_out_bits(cols_15_7_io_bottom_out_bits)
  );
  ProcessingElement cols_0_8 ( // @[Stab.scala 85:60]
    .clock(cols_0_8_clock),
    .reset(cols_0_8_reset),
    .io_left_in_ready(cols_0_8_io_left_in_ready),
    .io_left_in_valid(cols_0_8_io_left_in_valid),
    .io_left_in_bits(cols_0_8_io_left_in_bits),
    .io_top_in_ready(cols_0_8_io_top_in_ready),
    .io_top_in_valid(cols_0_8_io_top_in_valid),
    .io_top_in_bits(cols_0_8_io_top_in_bits),
    .io_sum_ready(cols_0_8_io_sum_ready),
    .io_sum_valid(cols_0_8_io_sum_valid),
    .io_sum_bits(cols_0_8_io_sum_bits),
    .io_right_out_ready(cols_0_8_io_right_out_ready),
    .io_right_out_valid(cols_0_8_io_right_out_valid),
    .io_right_out_bits(cols_0_8_io_right_out_bits),
    .io_bottom_out_ready(cols_0_8_io_bottom_out_ready),
    .io_bottom_out_valid(cols_0_8_io_bottom_out_valid),
    .io_bottom_out_bits(cols_0_8_io_bottom_out_bits)
  );
  ProcessingElement cols_1_8 ( // @[Stab.scala 85:60]
    .clock(cols_1_8_clock),
    .reset(cols_1_8_reset),
    .io_left_in_ready(cols_1_8_io_left_in_ready),
    .io_left_in_valid(cols_1_8_io_left_in_valid),
    .io_left_in_bits(cols_1_8_io_left_in_bits),
    .io_top_in_ready(cols_1_8_io_top_in_ready),
    .io_top_in_valid(cols_1_8_io_top_in_valid),
    .io_top_in_bits(cols_1_8_io_top_in_bits),
    .io_sum_ready(cols_1_8_io_sum_ready),
    .io_sum_valid(cols_1_8_io_sum_valid),
    .io_sum_bits(cols_1_8_io_sum_bits),
    .io_right_out_ready(cols_1_8_io_right_out_ready),
    .io_right_out_valid(cols_1_8_io_right_out_valid),
    .io_right_out_bits(cols_1_8_io_right_out_bits),
    .io_bottom_out_ready(cols_1_8_io_bottom_out_ready),
    .io_bottom_out_valid(cols_1_8_io_bottom_out_valid),
    .io_bottom_out_bits(cols_1_8_io_bottom_out_bits)
  );
  ProcessingElement cols_2_8 ( // @[Stab.scala 85:60]
    .clock(cols_2_8_clock),
    .reset(cols_2_8_reset),
    .io_left_in_ready(cols_2_8_io_left_in_ready),
    .io_left_in_valid(cols_2_8_io_left_in_valid),
    .io_left_in_bits(cols_2_8_io_left_in_bits),
    .io_top_in_ready(cols_2_8_io_top_in_ready),
    .io_top_in_valid(cols_2_8_io_top_in_valid),
    .io_top_in_bits(cols_2_8_io_top_in_bits),
    .io_sum_ready(cols_2_8_io_sum_ready),
    .io_sum_valid(cols_2_8_io_sum_valid),
    .io_sum_bits(cols_2_8_io_sum_bits),
    .io_right_out_ready(cols_2_8_io_right_out_ready),
    .io_right_out_valid(cols_2_8_io_right_out_valid),
    .io_right_out_bits(cols_2_8_io_right_out_bits),
    .io_bottom_out_ready(cols_2_8_io_bottom_out_ready),
    .io_bottom_out_valid(cols_2_8_io_bottom_out_valid),
    .io_bottom_out_bits(cols_2_8_io_bottom_out_bits)
  );
  ProcessingElement cols_3_8 ( // @[Stab.scala 85:60]
    .clock(cols_3_8_clock),
    .reset(cols_3_8_reset),
    .io_left_in_ready(cols_3_8_io_left_in_ready),
    .io_left_in_valid(cols_3_8_io_left_in_valid),
    .io_left_in_bits(cols_3_8_io_left_in_bits),
    .io_top_in_ready(cols_3_8_io_top_in_ready),
    .io_top_in_valid(cols_3_8_io_top_in_valid),
    .io_top_in_bits(cols_3_8_io_top_in_bits),
    .io_sum_ready(cols_3_8_io_sum_ready),
    .io_sum_valid(cols_3_8_io_sum_valid),
    .io_sum_bits(cols_3_8_io_sum_bits),
    .io_right_out_ready(cols_3_8_io_right_out_ready),
    .io_right_out_valid(cols_3_8_io_right_out_valid),
    .io_right_out_bits(cols_3_8_io_right_out_bits),
    .io_bottom_out_ready(cols_3_8_io_bottom_out_ready),
    .io_bottom_out_valid(cols_3_8_io_bottom_out_valid),
    .io_bottom_out_bits(cols_3_8_io_bottom_out_bits)
  );
  ProcessingElement cols_4_8 ( // @[Stab.scala 85:60]
    .clock(cols_4_8_clock),
    .reset(cols_4_8_reset),
    .io_left_in_ready(cols_4_8_io_left_in_ready),
    .io_left_in_valid(cols_4_8_io_left_in_valid),
    .io_left_in_bits(cols_4_8_io_left_in_bits),
    .io_top_in_ready(cols_4_8_io_top_in_ready),
    .io_top_in_valid(cols_4_8_io_top_in_valid),
    .io_top_in_bits(cols_4_8_io_top_in_bits),
    .io_sum_ready(cols_4_8_io_sum_ready),
    .io_sum_valid(cols_4_8_io_sum_valid),
    .io_sum_bits(cols_4_8_io_sum_bits),
    .io_right_out_ready(cols_4_8_io_right_out_ready),
    .io_right_out_valid(cols_4_8_io_right_out_valid),
    .io_right_out_bits(cols_4_8_io_right_out_bits),
    .io_bottom_out_ready(cols_4_8_io_bottom_out_ready),
    .io_bottom_out_valid(cols_4_8_io_bottom_out_valid),
    .io_bottom_out_bits(cols_4_8_io_bottom_out_bits)
  );
  ProcessingElement cols_5_8 ( // @[Stab.scala 85:60]
    .clock(cols_5_8_clock),
    .reset(cols_5_8_reset),
    .io_left_in_ready(cols_5_8_io_left_in_ready),
    .io_left_in_valid(cols_5_8_io_left_in_valid),
    .io_left_in_bits(cols_5_8_io_left_in_bits),
    .io_top_in_ready(cols_5_8_io_top_in_ready),
    .io_top_in_valid(cols_5_8_io_top_in_valid),
    .io_top_in_bits(cols_5_8_io_top_in_bits),
    .io_sum_ready(cols_5_8_io_sum_ready),
    .io_sum_valid(cols_5_8_io_sum_valid),
    .io_sum_bits(cols_5_8_io_sum_bits),
    .io_right_out_ready(cols_5_8_io_right_out_ready),
    .io_right_out_valid(cols_5_8_io_right_out_valid),
    .io_right_out_bits(cols_5_8_io_right_out_bits),
    .io_bottom_out_ready(cols_5_8_io_bottom_out_ready),
    .io_bottom_out_valid(cols_5_8_io_bottom_out_valid),
    .io_bottom_out_bits(cols_5_8_io_bottom_out_bits)
  );
  ProcessingElement cols_6_8 ( // @[Stab.scala 85:60]
    .clock(cols_6_8_clock),
    .reset(cols_6_8_reset),
    .io_left_in_ready(cols_6_8_io_left_in_ready),
    .io_left_in_valid(cols_6_8_io_left_in_valid),
    .io_left_in_bits(cols_6_8_io_left_in_bits),
    .io_top_in_ready(cols_6_8_io_top_in_ready),
    .io_top_in_valid(cols_6_8_io_top_in_valid),
    .io_top_in_bits(cols_6_8_io_top_in_bits),
    .io_sum_ready(cols_6_8_io_sum_ready),
    .io_sum_valid(cols_6_8_io_sum_valid),
    .io_sum_bits(cols_6_8_io_sum_bits),
    .io_right_out_ready(cols_6_8_io_right_out_ready),
    .io_right_out_valid(cols_6_8_io_right_out_valid),
    .io_right_out_bits(cols_6_8_io_right_out_bits),
    .io_bottom_out_ready(cols_6_8_io_bottom_out_ready),
    .io_bottom_out_valid(cols_6_8_io_bottom_out_valid),
    .io_bottom_out_bits(cols_6_8_io_bottom_out_bits)
  );
  ProcessingElement cols_7_8 ( // @[Stab.scala 85:60]
    .clock(cols_7_8_clock),
    .reset(cols_7_8_reset),
    .io_left_in_ready(cols_7_8_io_left_in_ready),
    .io_left_in_valid(cols_7_8_io_left_in_valid),
    .io_left_in_bits(cols_7_8_io_left_in_bits),
    .io_top_in_ready(cols_7_8_io_top_in_ready),
    .io_top_in_valid(cols_7_8_io_top_in_valid),
    .io_top_in_bits(cols_7_8_io_top_in_bits),
    .io_sum_ready(cols_7_8_io_sum_ready),
    .io_sum_valid(cols_7_8_io_sum_valid),
    .io_sum_bits(cols_7_8_io_sum_bits),
    .io_right_out_ready(cols_7_8_io_right_out_ready),
    .io_right_out_valid(cols_7_8_io_right_out_valid),
    .io_right_out_bits(cols_7_8_io_right_out_bits),
    .io_bottom_out_ready(cols_7_8_io_bottom_out_ready),
    .io_bottom_out_valid(cols_7_8_io_bottom_out_valid),
    .io_bottom_out_bits(cols_7_8_io_bottom_out_bits)
  );
  ProcessingElement cols_8_8 ( // @[Stab.scala 85:60]
    .clock(cols_8_8_clock),
    .reset(cols_8_8_reset),
    .io_left_in_ready(cols_8_8_io_left_in_ready),
    .io_left_in_valid(cols_8_8_io_left_in_valid),
    .io_left_in_bits(cols_8_8_io_left_in_bits),
    .io_top_in_ready(cols_8_8_io_top_in_ready),
    .io_top_in_valid(cols_8_8_io_top_in_valid),
    .io_top_in_bits(cols_8_8_io_top_in_bits),
    .io_sum_ready(cols_8_8_io_sum_ready),
    .io_sum_valid(cols_8_8_io_sum_valid),
    .io_sum_bits(cols_8_8_io_sum_bits),
    .io_right_out_ready(cols_8_8_io_right_out_ready),
    .io_right_out_valid(cols_8_8_io_right_out_valid),
    .io_right_out_bits(cols_8_8_io_right_out_bits),
    .io_bottom_out_ready(cols_8_8_io_bottom_out_ready),
    .io_bottom_out_valid(cols_8_8_io_bottom_out_valid),
    .io_bottom_out_bits(cols_8_8_io_bottom_out_bits)
  );
  ProcessingElement cols_9_8 ( // @[Stab.scala 85:60]
    .clock(cols_9_8_clock),
    .reset(cols_9_8_reset),
    .io_left_in_ready(cols_9_8_io_left_in_ready),
    .io_left_in_valid(cols_9_8_io_left_in_valid),
    .io_left_in_bits(cols_9_8_io_left_in_bits),
    .io_top_in_ready(cols_9_8_io_top_in_ready),
    .io_top_in_valid(cols_9_8_io_top_in_valid),
    .io_top_in_bits(cols_9_8_io_top_in_bits),
    .io_sum_ready(cols_9_8_io_sum_ready),
    .io_sum_valid(cols_9_8_io_sum_valid),
    .io_sum_bits(cols_9_8_io_sum_bits),
    .io_right_out_ready(cols_9_8_io_right_out_ready),
    .io_right_out_valid(cols_9_8_io_right_out_valid),
    .io_right_out_bits(cols_9_8_io_right_out_bits),
    .io_bottom_out_ready(cols_9_8_io_bottom_out_ready),
    .io_bottom_out_valid(cols_9_8_io_bottom_out_valid),
    .io_bottom_out_bits(cols_9_8_io_bottom_out_bits)
  );
  ProcessingElement cols_10_8 ( // @[Stab.scala 85:60]
    .clock(cols_10_8_clock),
    .reset(cols_10_8_reset),
    .io_left_in_ready(cols_10_8_io_left_in_ready),
    .io_left_in_valid(cols_10_8_io_left_in_valid),
    .io_left_in_bits(cols_10_8_io_left_in_bits),
    .io_top_in_ready(cols_10_8_io_top_in_ready),
    .io_top_in_valid(cols_10_8_io_top_in_valid),
    .io_top_in_bits(cols_10_8_io_top_in_bits),
    .io_sum_ready(cols_10_8_io_sum_ready),
    .io_sum_valid(cols_10_8_io_sum_valid),
    .io_sum_bits(cols_10_8_io_sum_bits),
    .io_right_out_ready(cols_10_8_io_right_out_ready),
    .io_right_out_valid(cols_10_8_io_right_out_valid),
    .io_right_out_bits(cols_10_8_io_right_out_bits),
    .io_bottom_out_ready(cols_10_8_io_bottom_out_ready),
    .io_bottom_out_valid(cols_10_8_io_bottom_out_valid),
    .io_bottom_out_bits(cols_10_8_io_bottom_out_bits)
  );
  ProcessingElement cols_11_8 ( // @[Stab.scala 85:60]
    .clock(cols_11_8_clock),
    .reset(cols_11_8_reset),
    .io_left_in_ready(cols_11_8_io_left_in_ready),
    .io_left_in_valid(cols_11_8_io_left_in_valid),
    .io_left_in_bits(cols_11_8_io_left_in_bits),
    .io_top_in_ready(cols_11_8_io_top_in_ready),
    .io_top_in_valid(cols_11_8_io_top_in_valid),
    .io_top_in_bits(cols_11_8_io_top_in_bits),
    .io_sum_ready(cols_11_8_io_sum_ready),
    .io_sum_valid(cols_11_8_io_sum_valid),
    .io_sum_bits(cols_11_8_io_sum_bits),
    .io_right_out_ready(cols_11_8_io_right_out_ready),
    .io_right_out_valid(cols_11_8_io_right_out_valid),
    .io_right_out_bits(cols_11_8_io_right_out_bits),
    .io_bottom_out_ready(cols_11_8_io_bottom_out_ready),
    .io_bottom_out_valid(cols_11_8_io_bottom_out_valid),
    .io_bottom_out_bits(cols_11_8_io_bottom_out_bits)
  );
  ProcessingElement cols_12_8 ( // @[Stab.scala 85:60]
    .clock(cols_12_8_clock),
    .reset(cols_12_8_reset),
    .io_left_in_ready(cols_12_8_io_left_in_ready),
    .io_left_in_valid(cols_12_8_io_left_in_valid),
    .io_left_in_bits(cols_12_8_io_left_in_bits),
    .io_top_in_ready(cols_12_8_io_top_in_ready),
    .io_top_in_valid(cols_12_8_io_top_in_valid),
    .io_top_in_bits(cols_12_8_io_top_in_bits),
    .io_sum_ready(cols_12_8_io_sum_ready),
    .io_sum_valid(cols_12_8_io_sum_valid),
    .io_sum_bits(cols_12_8_io_sum_bits),
    .io_right_out_ready(cols_12_8_io_right_out_ready),
    .io_right_out_valid(cols_12_8_io_right_out_valid),
    .io_right_out_bits(cols_12_8_io_right_out_bits),
    .io_bottom_out_ready(cols_12_8_io_bottom_out_ready),
    .io_bottom_out_valid(cols_12_8_io_bottom_out_valid),
    .io_bottom_out_bits(cols_12_8_io_bottom_out_bits)
  );
  ProcessingElement cols_13_8 ( // @[Stab.scala 85:60]
    .clock(cols_13_8_clock),
    .reset(cols_13_8_reset),
    .io_left_in_ready(cols_13_8_io_left_in_ready),
    .io_left_in_valid(cols_13_8_io_left_in_valid),
    .io_left_in_bits(cols_13_8_io_left_in_bits),
    .io_top_in_ready(cols_13_8_io_top_in_ready),
    .io_top_in_valid(cols_13_8_io_top_in_valid),
    .io_top_in_bits(cols_13_8_io_top_in_bits),
    .io_sum_ready(cols_13_8_io_sum_ready),
    .io_sum_valid(cols_13_8_io_sum_valid),
    .io_sum_bits(cols_13_8_io_sum_bits),
    .io_right_out_ready(cols_13_8_io_right_out_ready),
    .io_right_out_valid(cols_13_8_io_right_out_valid),
    .io_right_out_bits(cols_13_8_io_right_out_bits),
    .io_bottom_out_ready(cols_13_8_io_bottom_out_ready),
    .io_bottom_out_valid(cols_13_8_io_bottom_out_valid),
    .io_bottom_out_bits(cols_13_8_io_bottom_out_bits)
  );
  ProcessingElement cols_14_8 ( // @[Stab.scala 85:60]
    .clock(cols_14_8_clock),
    .reset(cols_14_8_reset),
    .io_left_in_ready(cols_14_8_io_left_in_ready),
    .io_left_in_valid(cols_14_8_io_left_in_valid),
    .io_left_in_bits(cols_14_8_io_left_in_bits),
    .io_top_in_ready(cols_14_8_io_top_in_ready),
    .io_top_in_valid(cols_14_8_io_top_in_valid),
    .io_top_in_bits(cols_14_8_io_top_in_bits),
    .io_sum_ready(cols_14_8_io_sum_ready),
    .io_sum_valid(cols_14_8_io_sum_valid),
    .io_sum_bits(cols_14_8_io_sum_bits),
    .io_right_out_ready(cols_14_8_io_right_out_ready),
    .io_right_out_valid(cols_14_8_io_right_out_valid),
    .io_right_out_bits(cols_14_8_io_right_out_bits),
    .io_bottom_out_ready(cols_14_8_io_bottom_out_ready),
    .io_bottom_out_valid(cols_14_8_io_bottom_out_valid),
    .io_bottom_out_bits(cols_14_8_io_bottom_out_bits)
  );
  ProcessingElement cols_15_8 ( // @[Stab.scala 85:60]
    .clock(cols_15_8_clock),
    .reset(cols_15_8_reset),
    .io_left_in_ready(cols_15_8_io_left_in_ready),
    .io_left_in_valid(cols_15_8_io_left_in_valid),
    .io_left_in_bits(cols_15_8_io_left_in_bits),
    .io_top_in_ready(cols_15_8_io_top_in_ready),
    .io_top_in_valid(cols_15_8_io_top_in_valid),
    .io_top_in_bits(cols_15_8_io_top_in_bits),
    .io_sum_ready(cols_15_8_io_sum_ready),
    .io_sum_valid(cols_15_8_io_sum_valid),
    .io_sum_bits(cols_15_8_io_sum_bits),
    .io_right_out_ready(cols_15_8_io_right_out_ready),
    .io_right_out_valid(cols_15_8_io_right_out_valid),
    .io_right_out_bits(cols_15_8_io_right_out_bits),
    .io_bottom_out_ready(cols_15_8_io_bottom_out_ready),
    .io_bottom_out_valid(cols_15_8_io_bottom_out_valid),
    .io_bottom_out_bits(cols_15_8_io_bottom_out_bits)
  );
  ProcessingElement cols_0_9 ( // @[Stab.scala 85:60]
    .clock(cols_0_9_clock),
    .reset(cols_0_9_reset),
    .io_left_in_ready(cols_0_9_io_left_in_ready),
    .io_left_in_valid(cols_0_9_io_left_in_valid),
    .io_left_in_bits(cols_0_9_io_left_in_bits),
    .io_top_in_ready(cols_0_9_io_top_in_ready),
    .io_top_in_valid(cols_0_9_io_top_in_valid),
    .io_top_in_bits(cols_0_9_io_top_in_bits),
    .io_sum_ready(cols_0_9_io_sum_ready),
    .io_sum_valid(cols_0_9_io_sum_valid),
    .io_sum_bits(cols_0_9_io_sum_bits),
    .io_right_out_ready(cols_0_9_io_right_out_ready),
    .io_right_out_valid(cols_0_9_io_right_out_valid),
    .io_right_out_bits(cols_0_9_io_right_out_bits),
    .io_bottom_out_ready(cols_0_9_io_bottom_out_ready),
    .io_bottom_out_valid(cols_0_9_io_bottom_out_valid),
    .io_bottom_out_bits(cols_0_9_io_bottom_out_bits)
  );
  ProcessingElement cols_1_9 ( // @[Stab.scala 85:60]
    .clock(cols_1_9_clock),
    .reset(cols_1_9_reset),
    .io_left_in_ready(cols_1_9_io_left_in_ready),
    .io_left_in_valid(cols_1_9_io_left_in_valid),
    .io_left_in_bits(cols_1_9_io_left_in_bits),
    .io_top_in_ready(cols_1_9_io_top_in_ready),
    .io_top_in_valid(cols_1_9_io_top_in_valid),
    .io_top_in_bits(cols_1_9_io_top_in_bits),
    .io_sum_ready(cols_1_9_io_sum_ready),
    .io_sum_valid(cols_1_9_io_sum_valid),
    .io_sum_bits(cols_1_9_io_sum_bits),
    .io_right_out_ready(cols_1_9_io_right_out_ready),
    .io_right_out_valid(cols_1_9_io_right_out_valid),
    .io_right_out_bits(cols_1_9_io_right_out_bits),
    .io_bottom_out_ready(cols_1_9_io_bottom_out_ready),
    .io_bottom_out_valid(cols_1_9_io_bottom_out_valid),
    .io_bottom_out_bits(cols_1_9_io_bottom_out_bits)
  );
  ProcessingElement cols_2_9 ( // @[Stab.scala 85:60]
    .clock(cols_2_9_clock),
    .reset(cols_2_9_reset),
    .io_left_in_ready(cols_2_9_io_left_in_ready),
    .io_left_in_valid(cols_2_9_io_left_in_valid),
    .io_left_in_bits(cols_2_9_io_left_in_bits),
    .io_top_in_ready(cols_2_9_io_top_in_ready),
    .io_top_in_valid(cols_2_9_io_top_in_valid),
    .io_top_in_bits(cols_2_9_io_top_in_bits),
    .io_sum_ready(cols_2_9_io_sum_ready),
    .io_sum_valid(cols_2_9_io_sum_valid),
    .io_sum_bits(cols_2_9_io_sum_bits),
    .io_right_out_ready(cols_2_9_io_right_out_ready),
    .io_right_out_valid(cols_2_9_io_right_out_valid),
    .io_right_out_bits(cols_2_9_io_right_out_bits),
    .io_bottom_out_ready(cols_2_9_io_bottom_out_ready),
    .io_bottom_out_valid(cols_2_9_io_bottom_out_valid),
    .io_bottom_out_bits(cols_2_9_io_bottom_out_bits)
  );
  ProcessingElement cols_3_9 ( // @[Stab.scala 85:60]
    .clock(cols_3_9_clock),
    .reset(cols_3_9_reset),
    .io_left_in_ready(cols_3_9_io_left_in_ready),
    .io_left_in_valid(cols_3_9_io_left_in_valid),
    .io_left_in_bits(cols_3_9_io_left_in_bits),
    .io_top_in_ready(cols_3_9_io_top_in_ready),
    .io_top_in_valid(cols_3_9_io_top_in_valid),
    .io_top_in_bits(cols_3_9_io_top_in_bits),
    .io_sum_ready(cols_3_9_io_sum_ready),
    .io_sum_valid(cols_3_9_io_sum_valid),
    .io_sum_bits(cols_3_9_io_sum_bits),
    .io_right_out_ready(cols_3_9_io_right_out_ready),
    .io_right_out_valid(cols_3_9_io_right_out_valid),
    .io_right_out_bits(cols_3_9_io_right_out_bits),
    .io_bottom_out_ready(cols_3_9_io_bottom_out_ready),
    .io_bottom_out_valid(cols_3_9_io_bottom_out_valid),
    .io_bottom_out_bits(cols_3_9_io_bottom_out_bits)
  );
  ProcessingElement cols_4_9 ( // @[Stab.scala 85:60]
    .clock(cols_4_9_clock),
    .reset(cols_4_9_reset),
    .io_left_in_ready(cols_4_9_io_left_in_ready),
    .io_left_in_valid(cols_4_9_io_left_in_valid),
    .io_left_in_bits(cols_4_9_io_left_in_bits),
    .io_top_in_ready(cols_4_9_io_top_in_ready),
    .io_top_in_valid(cols_4_9_io_top_in_valid),
    .io_top_in_bits(cols_4_9_io_top_in_bits),
    .io_sum_ready(cols_4_9_io_sum_ready),
    .io_sum_valid(cols_4_9_io_sum_valid),
    .io_sum_bits(cols_4_9_io_sum_bits),
    .io_right_out_ready(cols_4_9_io_right_out_ready),
    .io_right_out_valid(cols_4_9_io_right_out_valid),
    .io_right_out_bits(cols_4_9_io_right_out_bits),
    .io_bottom_out_ready(cols_4_9_io_bottom_out_ready),
    .io_bottom_out_valid(cols_4_9_io_bottom_out_valid),
    .io_bottom_out_bits(cols_4_9_io_bottom_out_bits)
  );
  ProcessingElement cols_5_9 ( // @[Stab.scala 85:60]
    .clock(cols_5_9_clock),
    .reset(cols_5_9_reset),
    .io_left_in_ready(cols_5_9_io_left_in_ready),
    .io_left_in_valid(cols_5_9_io_left_in_valid),
    .io_left_in_bits(cols_5_9_io_left_in_bits),
    .io_top_in_ready(cols_5_9_io_top_in_ready),
    .io_top_in_valid(cols_5_9_io_top_in_valid),
    .io_top_in_bits(cols_5_9_io_top_in_bits),
    .io_sum_ready(cols_5_9_io_sum_ready),
    .io_sum_valid(cols_5_9_io_sum_valid),
    .io_sum_bits(cols_5_9_io_sum_bits),
    .io_right_out_ready(cols_5_9_io_right_out_ready),
    .io_right_out_valid(cols_5_9_io_right_out_valid),
    .io_right_out_bits(cols_5_9_io_right_out_bits),
    .io_bottom_out_ready(cols_5_9_io_bottom_out_ready),
    .io_bottom_out_valid(cols_5_9_io_bottom_out_valid),
    .io_bottom_out_bits(cols_5_9_io_bottom_out_bits)
  );
  ProcessingElement cols_6_9 ( // @[Stab.scala 85:60]
    .clock(cols_6_9_clock),
    .reset(cols_6_9_reset),
    .io_left_in_ready(cols_6_9_io_left_in_ready),
    .io_left_in_valid(cols_6_9_io_left_in_valid),
    .io_left_in_bits(cols_6_9_io_left_in_bits),
    .io_top_in_ready(cols_6_9_io_top_in_ready),
    .io_top_in_valid(cols_6_9_io_top_in_valid),
    .io_top_in_bits(cols_6_9_io_top_in_bits),
    .io_sum_ready(cols_6_9_io_sum_ready),
    .io_sum_valid(cols_6_9_io_sum_valid),
    .io_sum_bits(cols_6_9_io_sum_bits),
    .io_right_out_ready(cols_6_9_io_right_out_ready),
    .io_right_out_valid(cols_6_9_io_right_out_valid),
    .io_right_out_bits(cols_6_9_io_right_out_bits),
    .io_bottom_out_ready(cols_6_9_io_bottom_out_ready),
    .io_bottom_out_valid(cols_6_9_io_bottom_out_valid),
    .io_bottom_out_bits(cols_6_9_io_bottom_out_bits)
  );
  ProcessingElement cols_7_9 ( // @[Stab.scala 85:60]
    .clock(cols_7_9_clock),
    .reset(cols_7_9_reset),
    .io_left_in_ready(cols_7_9_io_left_in_ready),
    .io_left_in_valid(cols_7_9_io_left_in_valid),
    .io_left_in_bits(cols_7_9_io_left_in_bits),
    .io_top_in_ready(cols_7_9_io_top_in_ready),
    .io_top_in_valid(cols_7_9_io_top_in_valid),
    .io_top_in_bits(cols_7_9_io_top_in_bits),
    .io_sum_ready(cols_7_9_io_sum_ready),
    .io_sum_valid(cols_7_9_io_sum_valid),
    .io_sum_bits(cols_7_9_io_sum_bits),
    .io_right_out_ready(cols_7_9_io_right_out_ready),
    .io_right_out_valid(cols_7_9_io_right_out_valid),
    .io_right_out_bits(cols_7_9_io_right_out_bits),
    .io_bottom_out_ready(cols_7_9_io_bottom_out_ready),
    .io_bottom_out_valid(cols_7_9_io_bottom_out_valid),
    .io_bottom_out_bits(cols_7_9_io_bottom_out_bits)
  );
  ProcessingElement cols_8_9 ( // @[Stab.scala 85:60]
    .clock(cols_8_9_clock),
    .reset(cols_8_9_reset),
    .io_left_in_ready(cols_8_9_io_left_in_ready),
    .io_left_in_valid(cols_8_9_io_left_in_valid),
    .io_left_in_bits(cols_8_9_io_left_in_bits),
    .io_top_in_ready(cols_8_9_io_top_in_ready),
    .io_top_in_valid(cols_8_9_io_top_in_valid),
    .io_top_in_bits(cols_8_9_io_top_in_bits),
    .io_sum_ready(cols_8_9_io_sum_ready),
    .io_sum_valid(cols_8_9_io_sum_valid),
    .io_sum_bits(cols_8_9_io_sum_bits),
    .io_right_out_ready(cols_8_9_io_right_out_ready),
    .io_right_out_valid(cols_8_9_io_right_out_valid),
    .io_right_out_bits(cols_8_9_io_right_out_bits),
    .io_bottom_out_ready(cols_8_9_io_bottom_out_ready),
    .io_bottom_out_valid(cols_8_9_io_bottom_out_valid),
    .io_bottom_out_bits(cols_8_9_io_bottom_out_bits)
  );
  ProcessingElement cols_9_9 ( // @[Stab.scala 85:60]
    .clock(cols_9_9_clock),
    .reset(cols_9_9_reset),
    .io_left_in_ready(cols_9_9_io_left_in_ready),
    .io_left_in_valid(cols_9_9_io_left_in_valid),
    .io_left_in_bits(cols_9_9_io_left_in_bits),
    .io_top_in_ready(cols_9_9_io_top_in_ready),
    .io_top_in_valid(cols_9_9_io_top_in_valid),
    .io_top_in_bits(cols_9_9_io_top_in_bits),
    .io_sum_ready(cols_9_9_io_sum_ready),
    .io_sum_valid(cols_9_9_io_sum_valid),
    .io_sum_bits(cols_9_9_io_sum_bits),
    .io_right_out_ready(cols_9_9_io_right_out_ready),
    .io_right_out_valid(cols_9_9_io_right_out_valid),
    .io_right_out_bits(cols_9_9_io_right_out_bits),
    .io_bottom_out_ready(cols_9_9_io_bottom_out_ready),
    .io_bottom_out_valid(cols_9_9_io_bottom_out_valid),
    .io_bottom_out_bits(cols_9_9_io_bottom_out_bits)
  );
  ProcessingElement cols_10_9 ( // @[Stab.scala 85:60]
    .clock(cols_10_9_clock),
    .reset(cols_10_9_reset),
    .io_left_in_ready(cols_10_9_io_left_in_ready),
    .io_left_in_valid(cols_10_9_io_left_in_valid),
    .io_left_in_bits(cols_10_9_io_left_in_bits),
    .io_top_in_ready(cols_10_9_io_top_in_ready),
    .io_top_in_valid(cols_10_9_io_top_in_valid),
    .io_top_in_bits(cols_10_9_io_top_in_bits),
    .io_sum_ready(cols_10_9_io_sum_ready),
    .io_sum_valid(cols_10_9_io_sum_valid),
    .io_sum_bits(cols_10_9_io_sum_bits),
    .io_right_out_ready(cols_10_9_io_right_out_ready),
    .io_right_out_valid(cols_10_9_io_right_out_valid),
    .io_right_out_bits(cols_10_9_io_right_out_bits),
    .io_bottom_out_ready(cols_10_9_io_bottom_out_ready),
    .io_bottom_out_valid(cols_10_9_io_bottom_out_valid),
    .io_bottom_out_bits(cols_10_9_io_bottom_out_bits)
  );
  ProcessingElement cols_11_9 ( // @[Stab.scala 85:60]
    .clock(cols_11_9_clock),
    .reset(cols_11_9_reset),
    .io_left_in_ready(cols_11_9_io_left_in_ready),
    .io_left_in_valid(cols_11_9_io_left_in_valid),
    .io_left_in_bits(cols_11_9_io_left_in_bits),
    .io_top_in_ready(cols_11_9_io_top_in_ready),
    .io_top_in_valid(cols_11_9_io_top_in_valid),
    .io_top_in_bits(cols_11_9_io_top_in_bits),
    .io_sum_ready(cols_11_9_io_sum_ready),
    .io_sum_valid(cols_11_9_io_sum_valid),
    .io_sum_bits(cols_11_9_io_sum_bits),
    .io_right_out_ready(cols_11_9_io_right_out_ready),
    .io_right_out_valid(cols_11_9_io_right_out_valid),
    .io_right_out_bits(cols_11_9_io_right_out_bits),
    .io_bottom_out_ready(cols_11_9_io_bottom_out_ready),
    .io_bottom_out_valid(cols_11_9_io_bottom_out_valid),
    .io_bottom_out_bits(cols_11_9_io_bottom_out_bits)
  );
  ProcessingElement cols_12_9 ( // @[Stab.scala 85:60]
    .clock(cols_12_9_clock),
    .reset(cols_12_9_reset),
    .io_left_in_ready(cols_12_9_io_left_in_ready),
    .io_left_in_valid(cols_12_9_io_left_in_valid),
    .io_left_in_bits(cols_12_9_io_left_in_bits),
    .io_top_in_ready(cols_12_9_io_top_in_ready),
    .io_top_in_valid(cols_12_9_io_top_in_valid),
    .io_top_in_bits(cols_12_9_io_top_in_bits),
    .io_sum_ready(cols_12_9_io_sum_ready),
    .io_sum_valid(cols_12_9_io_sum_valid),
    .io_sum_bits(cols_12_9_io_sum_bits),
    .io_right_out_ready(cols_12_9_io_right_out_ready),
    .io_right_out_valid(cols_12_9_io_right_out_valid),
    .io_right_out_bits(cols_12_9_io_right_out_bits),
    .io_bottom_out_ready(cols_12_9_io_bottom_out_ready),
    .io_bottom_out_valid(cols_12_9_io_bottom_out_valid),
    .io_bottom_out_bits(cols_12_9_io_bottom_out_bits)
  );
  ProcessingElement cols_13_9 ( // @[Stab.scala 85:60]
    .clock(cols_13_9_clock),
    .reset(cols_13_9_reset),
    .io_left_in_ready(cols_13_9_io_left_in_ready),
    .io_left_in_valid(cols_13_9_io_left_in_valid),
    .io_left_in_bits(cols_13_9_io_left_in_bits),
    .io_top_in_ready(cols_13_9_io_top_in_ready),
    .io_top_in_valid(cols_13_9_io_top_in_valid),
    .io_top_in_bits(cols_13_9_io_top_in_bits),
    .io_sum_ready(cols_13_9_io_sum_ready),
    .io_sum_valid(cols_13_9_io_sum_valid),
    .io_sum_bits(cols_13_9_io_sum_bits),
    .io_right_out_ready(cols_13_9_io_right_out_ready),
    .io_right_out_valid(cols_13_9_io_right_out_valid),
    .io_right_out_bits(cols_13_9_io_right_out_bits),
    .io_bottom_out_ready(cols_13_9_io_bottom_out_ready),
    .io_bottom_out_valid(cols_13_9_io_bottom_out_valid),
    .io_bottom_out_bits(cols_13_9_io_bottom_out_bits)
  );
  ProcessingElement cols_14_9 ( // @[Stab.scala 85:60]
    .clock(cols_14_9_clock),
    .reset(cols_14_9_reset),
    .io_left_in_ready(cols_14_9_io_left_in_ready),
    .io_left_in_valid(cols_14_9_io_left_in_valid),
    .io_left_in_bits(cols_14_9_io_left_in_bits),
    .io_top_in_ready(cols_14_9_io_top_in_ready),
    .io_top_in_valid(cols_14_9_io_top_in_valid),
    .io_top_in_bits(cols_14_9_io_top_in_bits),
    .io_sum_ready(cols_14_9_io_sum_ready),
    .io_sum_valid(cols_14_9_io_sum_valid),
    .io_sum_bits(cols_14_9_io_sum_bits),
    .io_right_out_ready(cols_14_9_io_right_out_ready),
    .io_right_out_valid(cols_14_9_io_right_out_valid),
    .io_right_out_bits(cols_14_9_io_right_out_bits),
    .io_bottom_out_ready(cols_14_9_io_bottom_out_ready),
    .io_bottom_out_valid(cols_14_9_io_bottom_out_valid),
    .io_bottom_out_bits(cols_14_9_io_bottom_out_bits)
  );
  ProcessingElement cols_15_9 ( // @[Stab.scala 85:60]
    .clock(cols_15_9_clock),
    .reset(cols_15_9_reset),
    .io_left_in_ready(cols_15_9_io_left_in_ready),
    .io_left_in_valid(cols_15_9_io_left_in_valid),
    .io_left_in_bits(cols_15_9_io_left_in_bits),
    .io_top_in_ready(cols_15_9_io_top_in_ready),
    .io_top_in_valid(cols_15_9_io_top_in_valid),
    .io_top_in_bits(cols_15_9_io_top_in_bits),
    .io_sum_ready(cols_15_9_io_sum_ready),
    .io_sum_valid(cols_15_9_io_sum_valid),
    .io_sum_bits(cols_15_9_io_sum_bits),
    .io_right_out_ready(cols_15_9_io_right_out_ready),
    .io_right_out_valid(cols_15_9_io_right_out_valid),
    .io_right_out_bits(cols_15_9_io_right_out_bits),
    .io_bottom_out_ready(cols_15_9_io_bottom_out_ready),
    .io_bottom_out_valid(cols_15_9_io_bottom_out_valid),
    .io_bottom_out_bits(cols_15_9_io_bottom_out_bits)
  );
  ProcessingElement cols_0_10 ( // @[Stab.scala 85:60]
    .clock(cols_0_10_clock),
    .reset(cols_0_10_reset),
    .io_left_in_ready(cols_0_10_io_left_in_ready),
    .io_left_in_valid(cols_0_10_io_left_in_valid),
    .io_left_in_bits(cols_0_10_io_left_in_bits),
    .io_top_in_ready(cols_0_10_io_top_in_ready),
    .io_top_in_valid(cols_0_10_io_top_in_valid),
    .io_top_in_bits(cols_0_10_io_top_in_bits),
    .io_sum_ready(cols_0_10_io_sum_ready),
    .io_sum_valid(cols_0_10_io_sum_valid),
    .io_sum_bits(cols_0_10_io_sum_bits),
    .io_right_out_ready(cols_0_10_io_right_out_ready),
    .io_right_out_valid(cols_0_10_io_right_out_valid),
    .io_right_out_bits(cols_0_10_io_right_out_bits),
    .io_bottom_out_ready(cols_0_10_io_bottom_out_ready),
    .io_bottom_out_valid(cols_0_10_io_bottom_out_valid),
    .io_bottom_out_bits(cols_0_10_io_bottom_out_bits)
  );
  ProcessingElement cols_1_10 ( // @[Stab.scala 85:60]
    .clock(cols_1_10_clock),
    .reset(cols_1_10_reset),
    .io_left_in_ready(cols_1_10_io_left_in_ready),
    .io_left_in_valid(cols_1_10_io_left_in_valid),
    .io_left_in_bits(cols_1_10_io_left_in_bits),
    .io_top_in_ready(cols_1_10_io_top_in_ready),
    .io_top_in_valid(cols_1_10_io_top_in_valid),
    .io_top_in_bits(cols_1_10_io_top_in_bits),
    .io_sum_ready(cols_1_10_io_sum_ready),
    .io_sum_valid(cols_1_10_io_sum_valid),
    .io_sum_bits(cols_1_10_io_sum_bits),
    .io_right_out_ready(cols_1_10_io_right_out_ready),
    .io_right_out_valid(cols_1_10_io_right_out_valid),
    .io_right_out_bits(cols_1_10_io_right_out_bits),
    .io_bottom_out_ready(cols_1_10_io_bottom_out_ready),
    .io_bottom_out_valid(cols_1_10_io_bottom_out_valid),
    .io_bottom_out_bits(cols_1_10_io_bottom_out_bits)
  );
  ProcessingElement cols_2_10 ( // @[Stab.scala 85:60]
    .clock(cols_2_10_clock),
    .reset(cols_2_10_reset),
    .io_left_in_ready(cols_2_10_io_left_in_ready),
    .io_left_in_valid(cols_2_10_io_left_in_valid),
    .io_left_in_bits(cols_2_10_io_left_in_bits),
    .io_top_in_ready(cols_2_10_io_top_in_ready),
    .io_top_in_valid(cols_2_10_io_top_in_valid),
    .io_top_in_bits(cols_2_10_io_top_in_bits),
    .io_sum_ready(cols_2_10_io_sum_ready),
    .io_sum_valid(cols_2_10_io_sum_valid),
    .io_sum_bits(cols_2_10_io_sum_bits),
    .io_right_out_ready(cols_2_10_io_right_out_ready),
    .io_right_out_valid(cols_2_10_io_right_out_valid),
    .io_right_out_bits(cols_2_10_io_right_out_bits),
    .io_bottom_out_ready(cols_2_10_io_bottom_out_ready),
    .io_bottom_out_valid(cols_2_10_io_bottom_out_valid),
    .io_bottom_out_bits(cols_2_10_io_bottom_out_bits)
  );
  ProcessingElement cols_3_10 ( // @[Stab.scala 85:60]
    .clock(cols_3_10_clock),
    .reset(cols_3_10_reset),
    .io_left_in_ready(cols_3_10_io_left_in_ready),
    .io_left_in_valid(cols_3_10_io_left_in_valid),
    .io_left_in_bits(cols_3_10_io_left_in_bits),
    .io_top_in_ready(cols_3_10_io_top_in_ready),
    .io_top_in_valid(cols_3_10_io_top_in_valid),
    .io_top_in_bits(cols_3_10_io_top_in_bits),
    .io_sum_ready(cols_3_10_io_sum_ready),
    .io_sum_valid(cols_3_10_io_sum_valid),
    .io_sum_bits(cols_3_10_io_sum_bits),
    .io_right_out_ready(cols_3_10_io_right_out_ready),
    .io_right_out_valid(cols_3_10_io_right_out_valid),
    .io_right_out_bits(cols_3_10_io_right_out_bits),
    .io_bottom_out_ready(cols_3_10_io_bottom_out_ready),
    .io_bottom_out_valid(cols_3_10_io_bottom_out_valid),
    .io_bottom_out_bits(cols_3_10_io_bottom_out_bits)
  );
  ProcessingElement cols_4_10 ( // @[Stab.scala 85:60]
    .clock(cols_4_10_clock),
    .reset(cols_4_10_reset),
    .io_left_in_ready(cols_4_10_io_left_in_ready),
    .io_left_in_valid(cols_4_10_io_left_in_valid),
    .io_left_in_bits(cols_4_10_io_left_in_bits),
    .io_top_in_ready(cols_4_10_io_top_in_ready),
    .io_top_in_valid(cols_4_10_io_top_in_valid),
    .io_top_in_bits(cols_4_10_io_top_in_bits),
    .io_sum_ready(cols_4_10_io_sum_ready),
    .io_sum_valid(cols_4_10_io_sum_valid),
    .io_sum_bits(cols_4_10_io_sum_bits),
    .io_right_out_ready(cols_4_10_io_right_out_ready),
    .io_right_out_valid(cols_4_10_io_right_out_valid),
    .io_right_out_bits(cols_4_10_io_right_out_bits),
    .io_bottom_out_ready(cols_4_10_io_bottom_out_ready),
    .io_bottom_out_valid(cols_4_10_io_bottom_out_valid),
    .io_bottom_out_bits(cols_4_10_io_bottom_out_bits)
  );
  ProcessingElement cols_5_10 ( // @[Stab.scala 85:60]
    .clock(cols_5_10_clock),
    .reset(cols_5_10_reset),
    .io_left_in_ready(cols_5_10_io_left_in_ready),
    .io_left_in_valid(cols_5_10_io_left_in_valid),
    .io_left_in_bits(cols_5_10_io_left_in_bits),
    .io_top_in_ready(cols_5_10_io_top_in_ready),
    .io_top_in_valid(cols_5_10_io_top_in_valid),
    .io_top_in_bits(cols_5_10_io_top_in_bits),
    .io_sum_ready(cols_5_10_io_sum_ready),
    .io_sum_valid(cols_5_10_io_sum_valid),
    .io_sum_bits(cols_5_10_io_sum_bits),
    .io_right_out_ready(cols_5_10_io_right_out_ready),
    .io_right_out_valid(cols_5_10_io_right_out_valid),
    .io_right_out_bits(cols_5_10_io_right_out_bits),
    .io_bottom_out_ready(cols_5_10_io_bottom_out_ready),
    .io_bottom_out_valid(cols_5_10_io_bottom_out_valid),
    .io_bottom_out_bits(cols_5_10_io_bottom_out_bits)
  );
  ProcessingElement cols_6_10 ( // @[Stab.scala 85:60]
    .clock(cols_6_10_clock),
    .reset(cols_6_10_reset),
    .io_left_in_ready(cols_6_10_io_left_in_ready),
    .io_left_in_valid(cols_6_10_io_left_in_valid),
    .io_left_in_bits(cols_6_10_io_left_in_bits),
    .io_top_in_ready(cols_6_10_io_top_in_ready),
    .io_top_in_valid(cols_6_10_io_top_in_valid),
    .io_top_in_bits(cols_6_10_io_top_in_bits),
    .io_sum_ready(cols_6_10_io_sum_ready),
    .io_sum_valid(cols_6_10_io_sum_valid),
    .io_sum_bits(cols_6_10_io_sum_bits),
    .io_right_out_ready(cols_6_10_io_right_out_ready),
    .io_right_out_valid(cols_6_10_io_right_out_valid),
    .io_right_out_bits(cols_6_10_io_right_out_bits),
    .io_bottom_out_ready(cols_6_10_io_bottom_out_ready),
    .io_bottom_out_valid(cols_6_10_io_bottom_out_valid),
    .io_bottom_out_bits(cols_6_10_io_bottom_out_bits)
  );
  ProcessingElement cols_7_10 ( // @[Stab.scala 85:60]
    .clock(cols_7_10_clock),
    .reset(cols_7_10_reset),
    .io_left_in_ready(cols_7_10_io_left_in_ready),
    .io_left_in_valid(cols_7_10_io_left_in_valid),
    .io_left_in_bits(cols_7_10_io_left_in_bits),
    .io_top_in_ready(cols_7_10_io_top_in_ready),
    .io_top_in_valid(cols_7_10_io_top_in_valid),
    .io_top_in_bits(cols_7_10_io_top_in_bits),
    .io_sum_ready(cols_7_10_io_sum_ready),
    .io_sum_valid(cols_7_10_io_sum_valid),
    .io_sum_bits(cols_7_10_io_sum_bits),
    .io_right_out_ready(cols_7_10_io_right_out_ready),
    .io_right_out_valid(cols_7_10_io_right_out_valid),
    .io_right_out_bits(cols_7_10_io_right_out_bits),
    .io_bottom_out_ready(cols_7_10_io_bottom_out_ready),
    .io_bottom_out_valid(cols_7_10_io_bottom_out_valid),
    .io_bottom_out_bits(cols_7_10_io_bottom_out_bits)
  );
  ProcessingElement cols_8_10 ( // @[Stab.scala 85:60]
    .clock(cols_8_10_clock),
    .reset(cols_8_10_reset),
    .io_left_in_ready(cols_8_10_io_left_in_ready),
    .io_left_in_valid(cols_8_10_io_left_in_valid),
    .io_left_in_bits(cols_8_10_io_left_in_bits),
    .io_top_in_ready(cols_8_10_io_top_in_ready),
    .io_top_in_valid(cols_8_10_io_top_in_valid),
    .io_top_in_bits(cols_8_10_io_top_in_bits),
    .io_sum_ready(cols_8_10_io_sum_ready),
    .io_sum_valid(cols_8_10_io_sum_valid),
    .io_sum_bits(cols_8_10_io_sum_bits),
    .io_right_out_ready(cols_8_10_io_right_out_ready),
    .io_right_out_valid(cols_8_10_io_right_out_valid),
    .io_right_out_bits(cols_8_10_io_right_out_bits),
    .io_bottom_out_ready(cols_8_10_io_bottom_out_ready),
    .io_bottom_out_valid(cols_8_10_io_bottom_out_valid),
    .io_bottom_out_bits(cols_8_10_io_bottom_out_bits)
  );
  ProcessingElement cols_9_10 ( // @[Stab.scala 85:60]
    .clock(cols_9_10_clock),
    .reset(cols_9_10_reset),
    .io_left_in_ready(cols_9_10_io_left_in_ready),
    .io_left_in_valid(cols_9_10_io_left_in_valid),
    .io_left_in_bits(cols_9_10_io_left_in_bits),
    .io_top_in_ready(cols_9_10_io_top_in_ready),
    .io_top_in_valid(cols_9_10_io_top_in_valid),
    .io_top_in_bits(cols_9_10_io_top_in_bits),
    .io_sum_ready(cols_9_10_io_sum_ready),
    .io_sum_valid(cols_9_10_io_sum_valid),
    .io_sum_bits(cols_9_10_io_sum_bits),
    .io_right_out_ready(cols_9_10_io_right_out_ready),
    .io_right_out_valid(cols_9_10_io_right_out_valid),
    .io_right_out_bits(cols_9_10_io_right_out_bits),
    .io_bottom_out_ready(cols_9_10_io_bottom_out_ready),
    .io_bottom_out_valid(cols_9_10_io_bottom_out_valid),
    .io_bottom_out_bits(cols_9_10_io_bottom_out_bits)
  );
  ProcessingElement cols_10_10 ( // @[Stab.scala 85:60]
    .clock(cols_10_10_clock),
    .reset(cols_10_10_reset),
    .io_left_in_ready(cols_10_10_io_left_in_ready),
    .io_left_in_valid(cols_10_10_io_left_in_valid),
    .io_left_in_bits(cols_10_10_io_left_in_bits),
    .io_top_in_ready(cols_10_10_io_top_in_ready),
    .io_top_in_valid(cols_10_10_io_top_in_valid),
    .io_top_in_bits(cols_10_10_io_top_in_bits),
    .io_sum_ready(cols_10_10_io_sum_ready),
    .io_sum_valid(cols_10_10_io_sum_valid),
    .io_sum_bits(cols_10_10_io_sum_bits),
    .io_right_out_ready(cols_10_10_io_right_out_ready),
    .io_right_out_valid(cols_10_10_io_right_out_valid),
    .io_right_out_bits(cols_10_10_io_right_out_bits),
    .io_bottom_out_ready(cols_10_10_io_bottom_out_ready),
    .io_bottom_out_valid(cols_10_10_io_bottom_out_valid),
    .io_bottom_out_bits(cols_10_10_io_bottom_out_bits)
  );
  ProcessingElement cols_11_10 ( // @[Stab.scala 85:60]
    .clock(cols_11_10_clock),
    .reset(cols_11_10_reset),
    .io_left_in_ready(cols_11_10_io_left_in_ready),
    .io_left_in_valid(cols_11_10_io_left_in_valid),
    .io_left_in_bits(cols_11_10_io_left_in_bits),
    .io_top_in_ready(cols_11_10_io_top_in_ready),
    .io_top_in_valid(cols_11_10_io_top_in_valid),
    .io_top_in_bits(cols_11_10_io_top_in_bits),
    .io_sum_ready(cols_11_10_io_sum_ready),
    .io_sum_valid(cols_11_10_io_sum_valid),
    .io_sum_bits(cols_11_10_io_sum_bits),
    .io_right_out_ready(cols_11_10_io_right_out_ready),
    .io_right_out_valid(cols_11_10_io_right_out_valid),
    .io_right_out_bits(cols_11_10_io_right_out_bits),
    .io_bottom_out_ready(cols_11_10_io_bottom_out_ready),
    .io_bottom_out_valid(cols_11_10_io_bottom_out_valid),
    .io_bottom_out_bits(cols_11_10_io_bottom_out_bits)
  );
  ProcessingElement cols_12_10 ( // @[Stab.scala 85:60]
    .clock(cols_12_10_clock),
    .reset(cols_12_10_reset),
    .io_left_in_ready(cols_12_10_io_left_in_ready),
    .io_left_in_valid(cols_12_10_io_left_in_valid),
    .io_left_in_bits(cols_12_10_io_left_in_bits),
    .io_top_in_ready(cols_12_10_io_top_in_ready),
    .io_top_in_valid(cols_12_10_io_top_in_valid),
    .io_top_in_bits(cols_12_10_io_top_in_bits),
    .io_sum_ready(cols_12_10_io_sum_ready),
    .io_sum_valid(cols_12_10_io_sum_valid),
    .io_sum_bits(cols_12_10_io_sum_bits),
    .io_right_out_ready(cols_12_10_io_right_out_ready),
    .io_right_out_valid(cols_12_10_io_right_out_valid),
    .io_right_out_bits(cols_12_10_io_right_out_bits),
    .io_bottom_out_ready(cols_12_10_io_bottom_out_ready),
    .io_bottom_out_valid(cols_12_10_io_bottom_out_valid),
    .io_bottom_out_bits(cols_12_10_io_bottom_out_bits)
  );
  ProcessingElement cols_13_10 ( // @[Stab.scala 85:60]
    .clock(cols_13_10_clock),
    .reset(cols_13_10_reset),
    .io_left_in_ready(cols_13_10_io_left_in_ready),
    .io_left_in_valid(cols_13_10_io_left_in_valid),
    .io_left_in_bits(cols_13_10_io_left_in_bits),
    .io_top_in_ready(cols_13_10_io_top_in_ready),
    .io_top_in_valid(cols_13_10_io_top_in_valid),
    .io_top_in_bits(cols_13_10_io_top_in_bits),
    .io_sum_ready(cols_13_10_io_sum_ready),
    .io_sum_valid(cols_13_10_io_sum_valid),
    .io_sum_bits(cols_13_10_io_sum_bits),
    .io_right_out_ready(cols_13_10_io_right_out_ready),
    .io_right_out_valid(cols_13_10_io_right_out_valid),
    .io_right_out_bits(cols_13_10_io_right_out_bits),
    .io_bottom_out_ready(cols_13_10_io_bottom_out_ready),
    .io_bottom_out_valid(cols_13_10_io_bottom_out_valid),
    .io_bottom_out_bits(cols_13_10_io_bottom_out_bits)
  );
  ProcessingElement cols_14_10 ( // @[Stab.scala 85:60]
    .clock(cols_14_10_clock),
    .reset(cols_14_10_reset),
    .io_left_in_ready(cols_14_10_io_left_in_ready),
    .io_left_in_valid(cols_14_10_io_left_in_valid),
    .io_left_in_bits(cols_14_10_io_left_in_bits),
    .io_top_in_ready(cols_14_10_io_top_in_ready),
    .io_top_in_valid(cols_14_10_io_top_in_valid),
    .io_top_in_bits(cols_14_10_io_top_in_bits),
    .io_sum_ready(cols_14_10_io_sum_ready),
    .io_sum_valid(cols_14_10_io_sum_valid),
    .io_sum_bits(cols_14_10_io_sum_bits),
    .io_right_out_ready(cols_14_10_io_right_out_ready),
    .io_right_out_valid(cols_14_10_io_right_out_valid),
    .io_right_out_bits(cols_14_10_io_right_out_bits),
    .io_bottom_out_ready(cols_14_10_io_bottom_out_ready),
    .io_bottom_out_valid(cols_14_10_io_bottom_out_valid),
    .io_bottom_out_bits(cols_14_10_io_bottom_out_bits)
  );
  ProcessingElement cols_15_10 ( // @[Stab.scala 85:60]
    .clock(cols_15_10_clock),
    .reset(cols_15_10_reset),
    .io_left_in_ready(cols_15_10_io_left_in_ready),
    .io_left_in_valid(cols_15_10_io_left_in_valid),
    .io_left_in_bits(cols_15_10_io_left_in_bits),
    .io_top_in_ready(cols_15_10_io_top_in_ready),
    .io_top_in_valid(cols_15_10_io_top_in_valid),
    .io_top_in_bits(cols_15_10_io_top_in_bits),
    .io_sum_ready(cols_15_10_io_sum_ready),
    .io_sum_valid(cols_15_10_io_sum_valid),
    .io_sum_bits(cols_15_10_io_sum_bits),
    .io_right_out_ready(cols_15_10_io_right_out_ready),
    .io_right_out_valid(cols_15_10_io_right_out_valid),
    .io_right_out_bits(cols_15_10_io_right_out_bits),
    .io_bottom_out_ready(cols_15_10_io_bottom_out_ready),
    .io_bottom_out_valid(cols_15_10_io_bottom_out_valid),
    .io_bottom_out_bits(cols_15_10_io_bottom_out_bits)
  );
  ProcessingElement cols_0_11 ( // @[Stab.scala 85:60]
    .clock(cols_0_11_clock),
    .reset(cols_0_11_reset),
    .io_left_in_ready(cols_0_11_io_left_in_ready),
    .io_left_in_valid(cols_0_11_io_left_in_valid),
    .io_left_in_bits(cols_0_11_io_left_in_bits),
    .io_top_in_ready(cols_0_11_io_top_in_ready),
    .io_top_in_valid(cols_0_11_io_top_in_valid),
    .io_top_in_bits(cols_0_11_io_top_in_bits),
    .io_sum_ready(cols_0_11_io_sum_ready),
    .io_sum_valid(cols_0_11_io_sum_valid),
    .io_sum_bits(cols_0_11_io_sum_bits),
    .io_right_out_ready(cols_0_11_io_right_out_ready),
    .io_right_out_valid(cols_0_11_io_right_out_valid),
    .io_right_out_bits(cols_0_11_io_right_out_bits),
    .io_bottom_out_ready(cols_0_11_io_bottom_out_ready),
    .io_bottom_out_valid(cols_0_11_io_bottom_out_valid),
    .io_bottom_out_bits(cols_0_11_io_bottom_out_bits)
  );
  ProcessingElement cols_1_11 ( // @[Stab.scala 85:60]
    .clock(cols_1_11_clock),
    .reset(cols_1_11_reset),
    .io_left_in_ready(cols_1_11_io_left_in_ready),
    .io_left_in_valid(cols_1_11_io_left_in_valid),
    .io_left_in_bits(cols_1_11_io_left_in_bits),
    .io_top_in_ready(cols_1_11_io_top_in_ready),
    .io_top_in_valid(cols_1_11_io_top_in_valid),
    .io_top_in_bits(cols_1_11_io_top_in_bits),
    .io_sum_ready(cols_1_11_io_sum_ready),
    .io_sum_valid(cols_1_11_io_sum_valid),
    .io_sum_bits(cols_1_11_io_sum_bits),
    .io_right_out_ready(cols_1_11_io_right_out_ready),
    .io_right_out_valid(cols_1_11_io_right_out_valid),
    .io_right_out_bits(cols_1_11_io_right_out_bits),
    .io_bottom_out_ready(cols_1_11_io_bottom_out_ready),
    .io_bottom_out_valid(cols_1_11_io_bottom_out_valid),
    .io_bottom_out_bits(cols_1_11_io_bottom_out_bits)
  );
  ProcessingElement cols_2_11 ( // @[Stab.scala 85:60]
    .clock(cols_2_11_clock),
    .reset(cols_2_11_reset),
    .io_left_in_ready(cols_2_11_io_left_in_ready),
    .io_left_in_valid(cols_2_11_io_left_in_valid),
    .io_left_in_bits(cols_2_11_io_left_in_bits),
    .io_top_in_ready(cols_2_11_io_top_in_ready),
    .io_top_in_valid(cols_2_11_io_top_in_valid),
    .io_top_in_bits(cols_2_11_io_top_in_bits),
    .io_sum_ready(cols_2_11_io_sum_ready),
    .io_sum_valid(cols_2_11_io_sum_valid),
    .io_sum_bits(cols_2_11_io_sum_bits),
    .io_right_out_ready(cols_2_11_io_right_out_ready),
    .io_right_out_valid(cols_2_11_io_right_out_valid),
    .io_right_out_bits(cols_2_11_io_right_out_bits),
    .io_bottom_out_ready(cols_2_11_io_bottom_out_ready),
    .io_bottom_out_valid(cols_2_11_io_bottom_out_valid),
    .io_bottom_out_bits(cols_2_11_io_bottom_out_bits)
  );
  ProcessingElement cols_3_11 ( // @[Stab.scala 85:60]
    .clock(cols_3_11_clock),
    .reset(cols_3_11_reset),
    .io_left_in_ready(cols_3_11_io_left_in_ready),
    .io_left_in_valid(cols_3_11_io_left_in_valid),
    .io_left_in_bits(cols_3_11_io_left_in_bits),
    .io_top_in_ready(cols_3_11_io_top_in_ready),
    .io_top_in_valid(cols_3_11_io_top_in_valid),
    .io_top_in_bits(cols_3_11_io_top_in_bits),
    .io_sum_ready(cols_3_11_io_sum_ready),
    .io_sum_valid(cols_3_11_io_sum_valid),
    .io_sum_bits(cols_3_11_io_sum_bits),
    .io_right_out_ready(cols_3_11_io_right_out_ready),
    .io_right_out_valid(cols_3_11_io_right_out_valid),
    .io_right_out_bits(cols_3_11_io_right_out_bits),
    .io_bottom_out_ready(cols_3_11_io_bottom_out_ready),
    .io_bottom_out_valid(cols_3_11_io_bottom_out_valid),
    .io_bottom_out_bits(cols_3_11_io_bottom_out_bits)
  );
  ProcessingElement cols_4_11 ( // @[Stab.scala 85:60]
    .clock(cols_4_11_clock),
    .reset(cols_4_11_reset),
    .io_left_in_ready(cols_4_11_io_left_in_ready),
    .io_left_in_valid(cols_4_11_io_left_in_valid),
    .io_left_in_bits(cols_4_11_io_left_in_bits),
    .io_top_in_ready(cols_4_11_io_top_in_ready),
    .io_top_in_valid(cols_4_11_io_top_in_valid),
    .io_top_in_bits(cols_4_11_io_top_in_bits),
    .io_sum_ready(cols_4_11_io_sum_ready),
    .io_sum_valid(cols_4_11_io_sum_valid),
    .io_sum_bits(cols_4_11_io_sum_bits),
    .io_right_out_ready(cols_4_11_io_right_out_ready),
    .io_right_out_valid(cols_4_11_io_right_out_valid),
    .io_right_out_bits(cols_4_11_io_right_out_bits),
    .io_bottom_out_ready(cols_4_11_io_bottom_out_ready),
    .io_bottom_out_valid(cols_4_11_io_bottom_out_valid),
    .io_bottom_out_bits(cols_4_11_io_bottom_out_bits)
  );
  ProcessingElement cols_5_11 ( // @[Stab.scala 85:60]
    .clock(cols_5_11_clock),
    .reset(cols_5_11_reset),
    .io_left_in_ready(cols_5_11_io_left_in_ready),
    .io_left_in_valid(cols_5_11_io_left_in_valid),
    .io_left_in_bits(cols_5_11_io_left_in_bits),
    .io_top_in_ready(cols_5_11_io_top_in_ready),
    .io_top_in_valid(cols_5_11_io_top_in_valid),
    .io_top_in_bits(cols_5_11_io_top_in_bits),
    .io_sum_ready(cols_5_11_io_sum_ready),
    .io_sum_valid(cols_5_11_io_sum_valid),
    .io_sum_bits(cols_5_11_io_sum_bits),
    .io_right_out_ready(cols_5_11_io_right_out_ready),
    .io_right_out_valid(cols_5_11_io_right_out_valid),
    .io_right_out_bits(cols_5_11_io_right_out_bits),
    .io_bottom_out_ready(cols_5_11_io_bottom_out_ready),
    .io_bottom_out_valid(cols_5_11_io_bottom_out_valid),
    .io_bottom_out_bits(cols_5_11_io_bottom_out_bits)
  );
  ProcessingElement cols_6_11 ( // @[Stab.scala 85:60]
    .clock(cols_6_11_clock),
    .reset(cols_6_11_reset),
    .io_left_in_ready(cols_6_11_io_left_in_ready),
    .io_left_in_valid(cols_6_11_io_left_in_valid),
    .io_left_in_bits(cols_6_11_io_left_in_bits),
    .io_top_in_ready(cols_6_11_io_top_in_ready),
    .io_top_in_valid(cols_6_11_io_top_in_valid),
    .io_top_in_bits(cols_6_11_io_top_in_bits),
    .io_sum_ready(cols_6_11_io_sum_ready),
    .io_sum_valid(cols_6_11_io_sum_valid),
    .io_sum_bits(cols_6_11_io_sum_bits),
    .io_right_out_ready(cols_6_11_io_right_out_ready),
    .io_right_out_valid(cols_6_11_io_right_out_valid),
    .io_right_out_bits(cols_6_11_io_right_out_bits),
    .io_bottom_out_ready(cols_6_11_io_bottom_out_ready),
    .io_bottom_out_valid(cols_6_11_io_bottom_out_valid),
    .io_bottom_out_bits(cols_6_11_io_bottom_out_bits)
  );
  ProcessingElement cols_7_11 ( // @[Stab.scala 85:60]
    .clock(cols_7_11_clock),
    .reset(cols_7_11_reset),
    .io_left_in_ready(cols_7_11_io_left_in_ready),
    .io_left_in_valid(cols_7_11_io_left_in_valid),
    .io_left_in_bits(cols_7_11_io_left_in_bits),
    .io_top_in_ready(cols_7_11_io_top_in_ready),
    .io_top_in_valid(cols_7_11_io_top_in_valid),
    .io_top_in_bits(cols_7_11_io_top_in_bits),
    .io_sum_ready(cols_7_11_io_sum_ready),
    .io_sum_valid(cols_7_11_io_sum_valid),
    .io_sum_bits(cols_7_11_io_sum_bits),
    .io_right_out_ready(cols_7_11_io_right_out_ready),
    .io_right_out_valid(cols_7_11_io_right_out_valid),
    .io_right_out_bits(cols_7_11_io_right_out_bits),
    .io_bottom_out_ready(cols_7_11_io_bottom_out_ready),
    .io_bottom_out_valid(cols_7_11_io_bottom_out_valid),
    .io_bottom_out_bits(cols_7_11_io_bottom_out_bits)
  );
  ProcessingElement cols_8_11 ( // @[Stab.scala 85:60]
    .clock(cols_8_11_clock),
    .reset(cols_8_11_reset),
    .io_left_in_ready(cols_8_11_io_left_in_ready),
    .io_left_in_valid(cols_8_11_io_left_in_valid),
    .io_left_in_bits(cols_8_11_io_left_in_bits),
    .io_top_in_ready(cols_8_11_io_top_in_ready),
    .io_top_in_valid(cols_8_11_io_top_in_valid),
    .io_top_in_bits(cols_8_11_io_top_in_bits),
    .io_sum_ready(cols_8_11_io_sum_ready),
    .io_sum_valid(cols_8_11_io_sum_valid),
    .io_sum_bits(cols_8_11_io_sum_bits),
    .io_right_out_ready(cols_8_11_io_right_out_ready),
    .io_right_out_valid(cols_8_11_io_right_out_valid),
    .io_right_out_bits(cols_8_11_io_right_out_bits),
    .io_bottom_out_ready(cols_8_11_io_bottom_out_ready),
    .io_bottom_out_valid(cols_8_11_io_bottom_out_valid),
    .io_bottom_out_bits(cols_8_11_io_bottom_out_bits)
  );
  ProcessingElement cols_9_11 ( // @[Stab.scala 85:60]
    .clock(cols_9_11_clock),
    .reset(cols_9_11_reset),
    .io_left_in_ready(cols_9_11_io_left_in_ready),
    .io_left_in_valid(cols_9_11_io_left_in_valid),
    .io_left_in_bits(cols_9_11_io_left_in_bits),
    .io_top_in_ready(cols_9_11_io_top_in_ready),
    .io_top_in_valid(cols_9_11_io_top_in_valid),
    .io_top_in_bits(cols_9_11_io_top_in_bits),
    .io_sum_ready(cols_9_11_io_sum_ready),
    .io_sum_valid(cols_9_11_io_sum_valid),
    .io_sum_bits(cols_9_11_io_sum_bits),
    .io_right_out_ready(cols_9_11_io_right_out_ready),
    .io_right_out_valid(cols_9_11_io_right_out_valid),
    .io_right_out_bits(cols_9_11_io_right_out_bits),
    .io_bottom_out_ready(cols_9_11_io_bottom_out_ready),
    .io_bottom_out_valid(cols_9_11_io_bottom_out_valid),
    .io_bottom_out_bits(cols_9_11_io_bottom_out_bits)
  );
  ProcessingElement cols_10_11 ( // @[Stab.scala 85:60]
    .clock(cols_10_11_clock),
    .reset(cols_10_11_reset),
    .io_left_in_ready(cols_10_11_io_left_in_ready),
    .io_left_in_valid(cols_10_11_io_left_in_valid),
    .io_left_in_bits(cols_10_11_io_left_in_bits),
    .io_top_in_ready(cols_10_11_io_top_in_ready),
    .io_top_in_valid(cols_10_11_io_top_in_valid),
    .io_top_in_bits(cols_10_11_io_top_in_bits),
    .io_sum_ready(cols_10_11_io_sum_ready),
    .io_sum_valid(cols_10_11_io_sum_valid),
    .io_sum_bits(cols_10_11_io_sum_bits),
    .io_right_out_ready(cols_10_11_io_right_out_ready),
    .io_right_out_valid(cols_10_11_io_right_out_valid),
    .io_right_out_bits(cols_10_11_io_right_out_bits),
    .io_bottom_out_ready(cols_10_11_io_bottom_out_ready),
    .io_bottom_out_valid(cols_10_11_io_bottom_out_valid),
    .io_bottom_out_bits(cols_10_11_io_bottom_out_bits)
  );
  ProcessingElement cols_11_11 ( // @[Stab.scala 85:60]
    .clock(cols_11_11_clock),
    .reset(cols_11_11_reset),
    .io_left_in_ready(cols_11_11_io_left_in_ready),
    .io_left_in_valid(cols_11_11_io_left_in_valid),
    .io_left_in_bits(cols_11_11_io_left_in_bits),
    .io_top_in_ready(cols_11_11_io_top_in_ready),
    .io_top_in_valid(cols_11_11_io_top_in_valid),
    .io_top_in_bits(cols_11_11_io_top_in_bits),
    .io_sum_ready(cols_11_11_io_sum_ready),
    .io_sum_valid(cols_11_11_io_sum_valid),
    .io_sum_bits(cols_11_11_io_sum_bits),
    .io_right_out_ready(cols_11_11_io_right_out_ready),
    .io_right_out_valid(cols_11_11_io_right_out_valid),
    .io_right_out_bits(cols_11_11_io_right_out_bits),
    .io_bottom_out_ready(cols_11_11_io_bottom_out_ready),
    .io_bottom_out_valid(cols_11_11_io_bottom_out_valid),
    .io_bottom_out_bits(cols_11_11_io_bottom_out_bits)
  );
  ProcessingElement cols_12_11 ( // @[Stab.scala 85:60]
    .clock(cols_12_11_clock),
    .reset(cols_12_11_reset),
    .io_left_in_ready(cols_12_11_io_left_in_ready),
    .io_left_in_valid(cols_12_11_io_left_in_valid),
    .io_left_in_bits(cols_12_11_io_left_in_bits),
    .io_top_in_ready(cols_12_11_io_top_in_ready),
    .io_top_in_valid(cols_12_11_io_top_in_valid),
    .io_top_in_bits(cols_12_11_io_top_in_bits),
    .io_sum_ready(cols_12_11_io_sum_ready),
    .io_sum_valid(cols_12_11_io_sum_valid),
    .io_sum_bits(cols_12_11_io_sum_bits),
    .io_right_out_ready(cols_12_11_io_right_out_ready),
    .io_right_out_valid(cols_12_11_io_right_out_valid),
    .io_right_out_bits(cols_12_11_io_right_out_bits),
    .io_bottom_out_ready(cols_12_11_io_bottom_out_ready),
    .io_bottom_out_valid(cols_12_11_io_bottom_out_valid),
    .io_bottom_out_bits(cols_12_11_io_bottom_out_bits)
  );
  ProcessingElement cols_13_11 ( // @[Stab.scala 85:60]
    .clock(cols_13_11_clock),
    .reset(cols_13_11_reset),
    .io_left_in_ready(cols_13_11_io_left_in_ready),
    .io_left_in_valid(cols_13_11_io_left_in_valid),
    .io_left_in_bits(cols_13_11_io_left_in_bits),
    .io_top_in_ready(cols_13_11_io_top_in_ready),
    .io_top_in_valid(cols_13_11_io_top_in_valid),
    .io_top_in_bits(cols_13_11_io_top_in_bits),
    .io_sum_ready(cols_13_11_io_sum_ready),
    .io_sum_valid(cols_13_11_io_sum_valid),
    .io_sum_bits(cols_13_11_io_sum_bits),
    .io_right_out_ready(cols_13_11_io_right_out_ready),
    .io_right_out_valid(cols_13_11_io_right_out_valid),
    .io_right_out_bits(cols_13_11_io_right_out_bits),
    .io_bottom_out_ready(cols_13_11_io_bottom_out_ready),
    .io_bottom_out_valid(cols_13_11_io_bottom_out_valid),
    .io_bottom_out_bits(cols_13_11_io_bottom_out_bits)
  );
  ProcessingElement cols_14_11 ( // @[Stab.scala 85:60]
    .clock(cols_14_11_clock),
    .reset(cols_14_11_reset),
    .io_left_in_ready(cols_14_11_io_left_in_ready),
    .io_left_in_valid(cols_14_11_io_left_in_valid),
    .io_left_in_bits(cols_14_11_io_left_in_bits),
    .io_top_in_ready(cols_14_11_io_top_in_ready),
    .io_top_in_valid(cols_14_11_io_top_in_valid),
    .io_top_in_bits(cols_14_11_io_top_in_bits),
    .io_sum_ready(cols_14_11_io_sum_ready),
    .io_sum_valid(cols_14_11_io_sum_valid),
    .io_sum_bits(cols_14_11_io_sum_bits),
    .io_right_out_ready(cols_14_11_io_right_out_ready),
    .io_right_out_valid(cols_14_11_io_right_out_valid),
    .io_right_out_bits(cols_14_11_io_right_out_bits),
    .io_bottom_out_ready(cols_14_11_io_bottom_out_ready),
    .io_bottom_out_valid(cols_14_11_io_bottom_out_valid),
    .io_bottom_out_bits(cols_14_11_io_bottom_out_bits)
  );
  ProcessingElement cols_15_11 ( // @[Stab.scala 85:60]
    .clock(cols_15_11_clock),
    .reset(cols_15_11_reset),
    .io_left_in_ready(cols_15_11_io_left_in_ready),
    .io_left_in_valid(cols_15_11_io_left_in_valid),
    .io_left_in_bits(cols_15_11_io_left_in_bits),
    .io_top_in_ready(cols_15_11_io_top_in_ready),
    .io_top_in_valid(cols_15_11_io_top_in_valid),
    .io_top_in_bits(cols_15_11_io_top_in_bits),
    .io_sum_ready(cols_15_11_io_sum_ready),
    .io_sum_valid(cols_15_11_io_sum_valid),
    .io_sum_bits(cols_15_11_io_sum_bits),
    .io_right_out_ready(cols_15_11_io_right_out_ready),
    .io_right_out_valid(cols_15_11_io_right_out_valid),
    .io_right_out_bits(cols_15_11_io_right_out_bits),
    .io_bottom_out_ready(cols_15_11_io_bottom_out_ready),
    .io_bottom_out_valid(cols_15_11_io_bottom_out_valid),
    .io_bottom_out_bits(cols_15_11_io_bottom_out_bits)
  );
  ProcessingElement cols_0_12 ( // @[Stab.scala 85:60]
    .clock(cols_0_12_clock),
    .reset(cols_0_12_reset),
    .io_left_in_ready(cols_0_12_io_left_in_ready),
    .io_left_in_valid(cols_0_12_io_left_in_valid),
    .io_left_in_bits(cols_0_12_io_left_in_bits),
    .io_top_in_ready(cols_0_12_io_top_in_ready),
    .io_top_in_valid(cols_0_12_io_top_in_valid),
    .io_top_in_bits(cols_0_12_io_top_in_bits),
    .io_sum_ready(cols_0_12_io_sum_ready),
    .io_sum_valid(cols_0_12_io_sum_valid),
    .io_sum_bits(cols_0_12_io_sum_bits),
    .io_right_out_ready(cols_0_12_io_right_out_ready),
    .io_right_out_valid(cols_0_12_io_right_out_valid),
    .io_right_out_bits(cols_0_12_io_right_out_bits),
    .io_bottom_out_ready(cols_0_12_io_bottom_out_ready),
    .io_bottom_out_valid(cols_0_12_io_bottom_out_valid),
    .io_bottom_out_bits(cols_0_12_io_bottom_out_bits)
  );
  ProcessingElement cols_1_12 ( // @[Stab.scala 85:60]
    .clock(cols_1_12_clock),
    .reset(cols_1_12_reset),
    .io_left_in_ready(cols_1_12_io_left_in_ready),
    .io_left_in_valid(cols_1_12_io_left_in_valid),
    .io_left_in_bits(cols_1_12_io_left_in_bits),
    .io_top_in_ready(cols_1_12_io_top_in_ready),
    .io_top_in_valid(cols_1_12_io_top_in_valid),
    .io_top_in_bits(cols_1_12_io_top_in_bits),
    .io_sum_ready(cols_1_12_io_sum_ready),
    .io_sum_valid(cols_1_12_io_sum_valid),
    .io_sum_bits(cols_1_12_io_sum_bits),
    .io_right_out_ready(cols_1_12_io_right_out_ready),
    .io_right_out_valid(cols_1_12_io_right_out_valid),
    .io_right_out_bits(cols_1_12_io_right_out_bits),
    .io_bottom_out_ready(cols_1_12_io_bottom_out_ready),
    .io_bottom_out_valid(cols_1_12_io_bottom_out_valid),
    .io_bottom_out_bits(cols_1_12_io_bottom_out_bits)
  );
  ProcessingElement cols_2_12 ( // @[Stab.scala 85:60]
    .clock(cols_2_12_clock),
    .reset(cols_2_12_reset),
    .io_left_in_ready(cols_2_12_io_left_in_ready),
    .io_left_in_valid(cols_2_12_io_left_in_valid),
    .io_left_in_bits(cols_2_12_io_left_in_bits),
    .io_top_in_ready(cols_2_12_io_top_in_ready),
    .io_top_in_valid(cols_2_12_io_top_in_valid),
    .io_top_in_bits(cols_2_12_io_top_in_bits),
    .io_sum_ready(cols_2_12_io_sum_ready),
    .io_sum_valid(cols_2_12_io_sum_valid),
    .io_sum_bits(cols_2_12_io_sum_bits),
    .io_right_out_ready(cols_2_12_io_right_out_ready),
    .io_right_out_valid(cols_2_12_io_right_out_valid),
    .io_right_out_bits(cols_2_12_io_right_out_bits),
    .io_bottom_out_ready(cols_2_12_io_bottom_out_ready),
    .io_bottom_out_valid(cols_2_12_io_bottom_out_valid),
    .io_bottom_out_bits(cols_2_12_io_bottom_out_bits)
  );
  ProcessingElement cols_3_12 ( // @[Stab.scala 85:60]
    .clock(cols_3_12_clock),
    .reset(cols_3_12_reset),
    .io_left_in_ready(cols_3_12_io_left_in_ready),
    .io_left_in_valid(cols_3_12_io_left_in_valid),
    .io_left_in_bits(cols_3_12_io_left_in_bits),
    .io_top_in_ready(cols_3_12_io_top_in_ready),
    .io_top_in_valid(cols_3_12_io_top_in_valid),
    .io_top_in_bits(cols_3_12_io_top_in_bits),
    .io_sum_ready(cols_3_12_io_sum_ready),
    .io_sum_valid(cols_3_12_io_sum_valid),
    .io_sum_bits(cols_3_12_io_sum_bits),
    .io_right_out_ready(cols_3_12_io_right_out_ready),
    .io_right_out_valid(cols_3_12_io_right_out_valid),
    .io_right_out_bits(cols_3_12_io_right_out_bits),
    .io_bottom_out_ready(cols_3_12_io_bottom_out_ready),
    .io_bottom_out_valid(cols_3_12_io_bottom_out_valid),
    .io_bottom_out_bits(cols_3_12_io_bottom_out_bits)
  );
  ProcessingElement cols_4_12 ( // @[Stab.scala 85:60]
    .clock(cols_4_12_clock),
    .reset(cols_4_12_reset),
    .io_left_in_ready(cols_4_12_io_left_in_ready),
    .io_left_in_valid(cols_4_12_io_left_in_valid),
    .io_left_in_bits(cols_4_12_io_left_in_bits),
    .io_top_in_ready(cols_4_12_io_top_in_ready),
    .io_top_in_valid(cols_4_12_io_top_in_valid),
    .io_top_in_bits(cols_4_12_io_top_in_bits),
    .io_sum_ready(cols_4_12_io_sum_ready),
    .io_sum_valid(cols_4_12_io_sum_valid),
    .io_sum_bits(cols_4_12_io_sum_bits),
    .io_right_out_ready(cols_4_12_io_right_out_ready),
    .io_right_out_valid(cols_4_12_io_right_out_valid),
    .io_right_out_bits(cols_4_12_io_right_out_bits),
    .io_bottom_out_ready(cols_4_12_io_bottom_out_ready),
    .io_bottom_out_valid(cols_4_12_io_bottom_out_valid),
    .io_bottom_out_bits(cols_4_12_io_bottom_out_bits)
  );
  ProcessingElement cols_5_12 ( // @[Stab.scala 85:60]
    .clock(cols_5_12_clock),
    .reset(cols_5_12_reset),
    .io_left_in_ready(cols_5_12_io_left_in_ready),
    .io_left_in_valid(cols_5_12_io_left_in_valid),
    .io_left_in_bits(cols_5_12_io_left_in_bits),
    .io_top_in_ready(cols_5_12_io_top_in_ready),
    .io_top_in_valid(cols_5_12_io_top_in_valid),
    .io_top_in_bits(cols_5_12_io_top_in_bits),
    .io_sum_ready(cols_5_12_io_sum_ready),
    .io_sum_valid(cols_5_12_io_sum_valid),
    .io_sum_bits(cols_5_12_io_sum_bits),
    .io_right_out_ready(cols_5_12_io_right_out_ready),
    .io_right_out_valid(cols_5_12_io_right_out_valid),
    .io_right_out_bits(cols_5_12_io_right_out_bits),
    .io_bottom_out_ready(cols_5_12_io_bottom_out_ready),
    .io_bottom_out_valid(cols_5_12_io_bottom_out_valid),
    .io_bottom_out_bits(cols_5_12_io_bottom_out_bits)
  );
  ProcessingElement cols_6_12 ( // @[Stab.scala 85:60]
    .clock(cols_6_12_clock),
    .reset(cols_6_12_reset),
    .io_left_in_ready(cols_6_12_io_left_in_ready),
    .io_left_in_valid(cols_6_12_io_left_in_valid),
    .io_left_in_bits(cols_6_12_io_left_in_bits),
    .io_top_in_ready(cols_6_12_io_top_in_ready),
    .io_top_in_valid(cols_6_12_io_top_in_valid),
    .io_top_in_bits(cols_6_12_io_top_in_bits),
    .io_sum_ready(cols_6_12_io_sum_ready),
    .io_sum_valid(cols_6_12_io_sum_valid),
    .io_sum_bits(cols_6_12_io_sum_bits),
    .io_right_out_ready(cols_6_12_io_right_out_ready),
    .io_right_out_valid(cols_6_12_io_right_out_valid),
    .io_right_out_bits(cols_6_12_io_right_out_bits),
    .io_bottom_out_ready(cols_6_12_io_bottom_out_ready),
    .io_bottom_out_valid(cols_6_12_io_bottom_out_valid),
    .io_bottom_out_bits(cols_6_12_io_bottom_out_bits)
  );
  ProcessingElement cols_7_12 ( // @[Stab.scala 85:60]
    .clock(cols_7_12_clock),
    .reset(cols_7_12_reset),
    .io_left_in_ready(cols_7_12_io_left_in_ready),
    .io_left_in_valid(cols_7_12_io_left_in_valid),
    .io_left_in_bits(cols_7_12_io_left_in_bits),
    .io_top_in_ready(cols_7_12_io_top_in_ready),
    .io_top_in_valid(cols_7_12_io_top_in_valid),
    .io_top_in_bits(cols_7_12_io_top_in_bits),
    .io_sum_ready(cols_7_12_io_sum_ready),
    .io_sum_valid(cols_7_12_io_sum_valid),
    .io_sum_bits(cols_7_12_io_sum_bits),
    .io_right_out_ready(cols_7_12_io_right_out_ready),
    .io_right_out_valid(cols_7_12_io_right_out_valid),
    .io_right_out_bits(cols_7_12_io_right_out_bits),
    .io_bottom_out_ready(cols_7_12_io_bottom_out_ready),
    .io_bottom_out_valid(cols_7_12_io_bottom_out_valid),
    .io_bottom_out_bits(cols_7_12_io_bottom_out_bits)
  );
  ProcessingElement cols_8_12 ( // @[Stab.scala 85:60]
    .clock(cols_8_12_clock),
    .reset(cols_8_12_reset),
    .io_left_in_ready(cols_8_12_io_left_in_ready),
    .io_left_in_valid(cols_8_12_io_left_in_valid),
    .io_left_in_bits(cols_8_12_io_left_in_bits),
    .io_top_in_ready(cols_8_12_io_top_in_ready),
    .io_top_in_valid(cols_8_12_io_top_in_valid),
    .io_top_in_bits(cols_8_12_io_top_in_bits),
    .io_sum_ready(cols_8_12_io_sum_ready),
    .io_sum_valid(cols_8_12_io_sum_valid),
    .io_sum_bits(cols_8_12_io_sum_bits),
    .io_right_out_ready(cols_8_12_io_right_out_ready),
    .io_right_out_valid(cols_8_12_io_right_out_valid),
    .io_right_out_bits(cols_8_12_io_right_out_bits),
    .io_bottom_out_ready(cols_8_12_io_bottom_out_ready),
    .io_bottom_out_valid(cols_8_12_io_bottom_out_valid),
    .io_bottom_out_bits(cols_8_12_io_bottom_out_bits)
  );
  ProcessingElement cols_9_12 ( // @[Stab.scala 85:60]
    .clock(cols_9_12_clock),
    .reset(cols_9_12_reset),
    .io_left_in_ready(cols_9_12_io_left_in_ready),
    .io_left_in_valid(cols_9_12_io_left_in_valid),
    .io_left_in_bits(cols_9_12_io_left_in_bits),
    .io_top_in_ready(cols_9_12_io_top_in_ready),
    .io_top_in_valid(cols_9_12_io_top_in_valid),
    .io_top_in_bits(cols_9_12_io_top_in_bits),
    .io_sum_ready(cols_9_12_io_sum_ready),
    .io_sum_valid(cols_9_12_io_sum_valid),
    .io_sum_bits(cols_9_12_io_sum_bits),
    .io_right_out_ready(cols_9_12_io_right_out_ready),
    .io_right_out_valid(cols_9_12_io_right_out_valid),
    .io_right_out_bits(cols_9_12_io_right_out_bits),
    .io_bottom_out_ready(cols_9_12_io_bottom_out_ready),
    .io_bottom_out_valid(cols_9_12_io_bottom_out_valid),
    .io_bottom_out_bits(cols_9_12_io_bottom_out_bits)
  );
  ProcessingElement cols_10_12 ( // @[Stab.scala 85:60]
    .clock(cols_10_12_clock),
    .reset(cols_10_12_reset),
    .io_left_in_ready(cols_10_12_io_left_in_ready),
    .io_left_in_valid(cols_10_12_io_left_in_valid),
    .io_left_in_bits(cols_10_12_io_left_in_bits),
    .io_top_in_ready(cols_10_12_io_top_in_ready),
    .io_top_in_valid(cols_10_12_io_top_in_valid),
    .io_top_in_bits(cols_10_12_io_top_in_bits),
    .io_sum_ready(cols_10_12_io_sum_ready),
    .io_sum_valid(cols_10_12_io_sum_valid),
    .io_sum_bits(cols_10_12_io_sum_bits),
    .io_right_out_ready(cols_10_12_io_right_out_ready),
    .io_right_out_valid(cols_10_12_io_right_out_valid),
    .io_right_out_bits(cols_10_12_io_right_out_bits),
    .io_bottom_out_ready(cols_10_12_io_bottom_out_ready),
    .io_bottom_out_valid(cols_10_12_io_bottom_out_valid),
    .io_bottom_out_bits(cols_10_12_io_bottom_out_bits)
  );
  ProcessingElement cols_11_12 ( // @[Stab.scala 85:60]
    .clock(cols_11_12_clock),
    .reset(cols_11_12_reset),
    .io_left_in_ready(cols_11_12_io_left_in_ready),
    .io_left_in_valid(cols_11_12_io_left_in_valid),
    .io_left_in_bits(cols_11_12_io_left_in_bits),
    .io_top_in_ready(cols_11_12_io_top_in_ready),
    .io_top_in_valid(cols_11_12_io_top_in_valid),
    .io_top_in_bits(cols_11_12_io_top_in_bits),
    .io_sum_ready(cols_11_12_io_sum_ready),
    .io_sum_valid(cols_11_12_io_sum_valid),
    .io_sum_bits(cols_11_12_io_sum_bits),
    .io_right_out_ready(cols_11_12_io_right_out_ready),
    .io_right_out_valid(cols_11_12_io_right_out_valid),
    .io_right_out_bits(cols_11_12_io_right_out_bits),
    .io_bottom_out_ready(cols_11_12_io_bottom_out_ready),
    .io_bottom_out_valid(cols_11_12_io_bottom_out_valid),
    .io_bottom_out_bits(cols_11_12_io_bottom_out_bits)
  );
  ProcessingElement cols_12_12 ( // @[Stab.scala 85:60]
    .clock(cols_12_12_clock),
    .reset(cols_12_12_reset),
    .io_left_in_ready(cols_12_12_io_left_in_ready),
    .io_left_in_valid(cols_12_12_io_left_in_valid),
    .io_left_in_bits(cols_12_12_io_left_in_bits),
    .io_top_in_ready(cols_12_12_io_top_in_ready),
    .io_top_in_valid(cols_12_12_io_top_in_valid),
    .io_top_in_bits(cols_12_12_io_top_in_bits),
    .io_sum_ready(cols_12_12_io_sum_ready),
    .io_sum_valid(cols_12_12_io_sum_valid),
    .io_sum_bits(cols_12_12_io_sum_bits),
    .io_right_out_ready(cols_12_12_io_right_out_ready),
    .io_right_out_valid(cols_12_12_io_right_out_valid),
    .io_right_out_bits(cols_12_12_io_right_out_bits),
    .io_bottom_out_ready(cols_12_12_io_bottom_out_ready),
    .io_bottom_out_valid(cols_12_12_io_bottom_out_valid),
    .io_bottom_out_bits(cols_12_12_io_bottom_out_bits)
  );
  ProcessingElement cols_13_12 ( // @[Stab.scala 85:60]
    .clock(cols_13_12_clock),
    .reset(cols_13_12_reset),
    .io_left_in_ready(cols_13_12_io_left_in_ready),
    .io_left_in_valid(cols_13_12_io_left_in_valid),
    .io_left_in_bits(cols_13_12_io_left_in_bits),
    .io_top_in_ready(cols_13_12_io_top_in_ready),
    .io_top_in_valid(cols_13_12_io_top_in_valid),
    .io_top_in_bits(cols_13_12_io_top_in_bits),
    .io_sum_ready(cols_13_12_io_sum_ready),
    .io_sum_valid(cols_13_12_io_sum_valid),
    .io_sum_bits(cols_13_12_io_sum_bits),
    .io_right_out_ready(cols_13_12_io_right_out_ready),
    .io_right_out_valid(cols_13_12_io_right_out_valid),
    .io_right_out_bits(cols_13_12_io_right_out_bits),
    .io_bottom_out_ready(cols_13_12_io_bottom_out_ready),
    .io_bottom_out_valid(cols_13_12_io_bottom_out_valid),
    .io_bottom_out_bits(cols_13_12_io_bottom_out_bits)
  );
  ProcessingElement cols_14_12 ( // @[Stab.scala 85:60]
    .clock(cols_14_12_clock),
    .reset(cols_14_12_reset),
    .io_left_in_ready(cols_14_12_io_left_in_ready),
    .io_left_in_valid(cols_14_12_io_left_in_valid),
    .io_left_in_bits(cols_14_12_io_left_in_bits),
    .io_top_in_ready(cols_14_12_io_top_in_ready),
    .io_top_in_valid(cols_14_12_io_top_in_valid),
    .io_top_in_bits(cols_14_12_io_top_in_bits),
    .io_sum_ready(cols_14_12_io_sum_ready),
    .io_sum_valid(cols_14_12_io_sum_valid),
    .io_sum_bits(cols_14_12_io_sum_bits),
    .io_right_out_ready(cols_14_12_io_right_out_ready),
    .io_right_out_valid(cols_14_12_io_right_out_valid),
    .io_right_out_bits(cols_14_12_io_right_out_bits),
    .io_bottom_out_ready(cols_14_12_io_bottom_out_ready),
    .io_bottom_out_valid(cols_14_12_io_bottom_out_valid),
    .io_bottom_out_bits(cols_14_12_io_bottom_out_bits)
  );
  ProcessingElement cols_15_12 ( // @[Stab.scala 85:60]
    .clock(cols_15_12_clock),
    .reset(cols_15_12_reset),
    .io_left_in_ready(cols_15_12_io_left_in_ready),
    .io_left_in_valid(cols_15_12_io_left_in_valid),
    .io_left_in_bits(cols_15_12_io_left_in_bits),
    .io_top_in_ready(cols_15_12_io_top_in_ready),
    .io_top_in_valid(cols_15_12_io_top_in_valid),
    .io_top_in_bits(cols_15_12_io_top_in_bits),
    .io_sum_ready(cols_15_12_io_sum_ready),
    .io_sum_valid(cols_15_12_io_sum_valid),
    .io_sum_bits(cols_15_12_io_sum_bits),
    .io_right_out_ready(cols_15_12_io_right_out_ready),
    .io_right_out_valid(cols_15_12_io_right_out_valid),
    .io_right_out_bits(cols_15_12_io_right_out_bits),
    .io_bottom_out_ready(cols_15_12_io_bottom_out_ready),
    .io_bottom_out_valid(cols_15_12_io_bottom_out_valid),
    .io_bottom_out_bits(cols_15_12_io_bottom_out_bits)
  );
  ProcessingElement cols_0_13 ( // @[Stab.scala 85:60]
    .clock(cols_0_13_clock),
    .reset(cols_0_13_reset),
    .io_left_in_ready(cols_0_13_io_left_in_ready),
    .io_left_in_valid(cols_0_13_io_left_in_valid),
    .io_left_in_bits(cols_0_13_io_left_in_bits),
    .io_top_in_ready(cols_0_13_io_top_in_ready),
    .io_top_in_valid(cols_0_13_io_top_in_valid),
    .io_top_in_bits(cols_0_13_io_top_in_bits),
    .io_sum_ready(cols_0_13_io_sum_ready),
    .io_sum_valid(cols_0_13_io_sum_valid),
    .io_sum_bits(cols_0_13_io_sum_bits),
    .io_right_out_ready(cols_0_13_io_right_out_ready),
    .io_right_out_valid(cols_0_13_io_right_out_valid),
    .io_right_out_bits(cols_0_13_io_right_out_bits),
    .io_bottom_out_ready(cols_0_13_io_bottom_out_ready),
    .io_bottom_out_valid(cols_0_13_io_bottom_out_valid),
    .io_bottom_out_bits(cols_0_13_io_bottom_out_bits)
  );
  ProcessingElement cols_1_13 ( // @[Stab.scala 85:60]
    .clock(cols_1_13_clock),
    .reset(cols_1_13_reset),
    .io_left_in_ready(cols_1_13_io_left_in_ready),
    .io_left_in_valid(cols_1_13_io_left_in_valid),
    .io_left_in_bits(cols_1_13_io_left_in_bits),
    .io_top_in_ready(cols_1_13_io_top_in_ready),
    .io_top_in_valid(cols_1_13_io_top_in_valid),
    .io_top_in_bits(cols_1_13_io_top_in_bits),
    .io_sum_ready(cols_1_13_io_sum_ready),
    .io_sum_valid(cols_1_13_io_sum_valid),
    .io_sum_bits(cols_1_13_io_sum_bits),
    .io_right_out_ready(cols_1_13_io_right_out_ready),
    .io_right_out_valid(cols_1_13_io_right_out_valid),
    .io_right_out_bits(cols_1_13_io_right_out_bits),
    .io_bottom_out_ready(cols_1_13_io_bottom_out_ready),
    .io_bottom_out_valid(cols_1_13_io_bottom_out_valid),
    .io_bottom_out_bits(cols_1_13_io_bottom_out_bits)
  );
  ProcessingElement cols_2_13 ( // @[Stab.scala 85:60]
    .clock(cols_2_13_clock),
    .reset(cols_2_13_reset),
    .io_left_in_ready(cols_2_13_io_left_in_ready),
    .io_left_in_valid(cols_2_13_io_left_in_valid),
    .io_left_in_bits(cols_2_13_io_left_in_bits),
    .io_top_in_ready(cols_2_13_io_top_in_ready),
    .io_top_in_valid(cols_2_13_io_top_in_valid),
    .io_top_in_bits(cols_2_13_io_top_in_bits),
    .io_sum_ready(cols_2_13_io_sum_ready),
    .io_sum_valid(cols_2_13_io_sum_valid),
    .io_sum_bits(cols_2_13_io_sum_bits),
    .io_right_out_ready(cols_2_13_io_right_out_ready),
    .io_right_out_valid(cols_2_13_io_right_out_valid),
    .io_right_out_bits(cols_2_13_io_right_out_bits),
    .io_bottom_out_ready(cols_2_13_io_bottom_out_ready),
    .io_bottom_out_valid(cols_2_13_io_bottom_out_valid),
    .io_bottom_out_bits(cols_2_13_io_bottom_out_bits)
  );
  ProcessingElement cols_3_13 ( // @[Stab.scala 85:60]
    .clock(cols_3_13_clock),
    .reset(cols_3_13_reset),
    .io_left_in_ready(cols_3_13_io_left_in_ready),
    .io_left_in_valid(cols_3_13_io_left_in_valid),
    .io_left_in_bits(cols_3_13_io_left_in_bits),
    .io_top_in_ready(cols_3_13_io_top_in_ready),
    .io_top_in_valid(cols_3_13_io_top_in_valid),
    .io_top_in_bits(cols_3_13_io_top_in_bits),
    .io_sum_ready(cols_3_13_io_sum_ready),
    .io_sum_valid(cols_3_13_io_sum_valid),
    .io_sum_bits(cols_3_13_io_sum_bits),
    .io_right_out_ready(cols_3_13_io_right_out_ready),
    .io_right_out_valid(cols_3_13_io_right_out_valid),
    .io_right_out_bits(cols_3_13_io_right_out_bits),
    .io_bottom_out_ready(cols_3_13_io_bottom_out_ready),
    .io_bottom_out_valid(cols_3_13_io_bottom_out_valid),
    .io_bottom_out_bits(cols_3_13_io_bottom_out_bits)
  );
  ProcessingElement cols_4_13 ( // @[Stab.scala 85:60]
    .clock(cols_4_13_clock),
    .reset(cols_4_13_reset),
    .io_left_in_ready(cols_4_13_io_left_in_ready),
    .io_left_in_valid(cols_4_13_io_left_in_valid),
    .io_left_in_bits(cols_4_13_io_left_in_bits),
    .io_top_in_ready(cols_4_13_io_top_in_ready),
    .io_top_in_valid(cols_4_13_io_top_in_valid),
    .io_top_in_bits(cols_4_13_io_top_in_bits),
    .io_sum_ready(cols_4_13_io_sum_ready),
    .io_sum_valid(cols_4_13_io_sum_valid),
    .io_sum_bits(cols_4_13_io_sum_bits),
    .io_right_out_ready(cols_4_13_io_right_out_ready),
    .io_right_out_valid(cols_4_13_io_right_out_valid),
    .io_right_out_bits(cols_4_13_io_right_out_bits),
    .io_bottom_out_ready(cols_4_13_io_bottom_out_ready),
    .io_bottom_out_valid(cols_4_13_io_bottom_out_valid),
    .io_bottom_out_bits(cols_4_13_io_bottom_out_bits)
  );
  ProcessingElement cols_5_13 ( // @[Stab.scala 85:60]
    .clock(cols_5_13_clock),
    .reset(cols_5_13_reset),
    .io_left_in_ready(cols_5_13_io_left_in_ready),
    .io_left_in_valid(cols_5_13_io_left_in_valid),
    .io_left_in_bits(cols_5_13_io_left_in_bits),
    .io_top_in_ready(cols_5_13_io_top_in_ready),
    .io_top_in_valid(cols_5_13_io_top_in_valid),
    .io_top_in_bits(cols_5_13_io_top_in_bits),
    .io_sum_ready(cols_5_13_io_sum_ready),
    .io_sum_valid(cols_5_13_io_sum_valid),
    .io_sum_bits(cols_5_13_io_sum_bits),
    .io_right_out_ready(cols_5_13_io_right_out_ready),
    .io_right_out_valid(cols_5_13_io_right_out_valid),
    .io_right_out_bits(cols_5_13_io_right_out_bits),
    .io_bottom_out_ready(cols_5_13_io_bottom_out_ready),
    .io_bottom_out_valid(cols_5_13_io_bottom_out_valid),
    .io_bottom_out_bits(cols_5_13_io_bottom_out_bits)
  );
  ProcessingElement cols_6_13 ( // @[Stab.scala 85:60]
    .clock(cols_6_13_clock),
    .reset(cols_6_13_reset),
    .io_left_in_ready(cols_6_13_io_left_in_ready),
    .io_left_in_valid(cols_6_13_io_left_in_valid),
    .io_left_in_bits(cols_6_13_io_left_in_bits),
    .io_top_in_ready(cols_6_13_io_top_in_ready),
    .io_top_in_valid(cols_6_13_io_top_in_valid),
    .io_top_in_bits(cols_6_13_io_top_in_bits),
    .io_sum_ready(cols_6_13_io_sum_ready),
    .io_sum_valid(cols_6_13_io_sum_valid),
    .io_sum_bits(cols_6_13_io_sum_bits),
    .io_right_out_ready(cols_6_13_io_right_out_ready),
    .io_right_out_valid(cols_6_13_io_right_out_valid),
    .io_right_out_bits(cols_6_13_io_right_out_bits),
    .io_bottom_out_ready(cols_6_13_io_bottom_out_ready),
    .io_bottom_out_valid(cols_6_13_io_bottom_out_valid),
    .io_bottom_out_bits(cols_6_13_io_bottom_out_bits)
  );
  ProcessingElement cols_7_13 ( // @[Stab.scala 85:60]
    .clock(cols_7_13_clock),
    .reset(cols_7_13_reset),
    .io_left_in_ready(cols_7_13_io_left_in_ready),
    .io_left_in_valid(cols_7_13_io_left_in_valid),
    .io_left_in_bits(cols_7_13_io_left_in_bits),
    .io_top_in_ready(cols_7_13_io_top_in_ready),
    .io_top_in_valid(cols_7_13_io_top_in_valid),
    .io_top_in_bits(cols_7_13_io_top_in_bits),
    .io_sum_ready(cols_7_13_io_sum_ready),
    .io_sum_valid(cols_7_13_io_sum_valid),
    .io_sum_bits(cols_7_13_io_sum_bits),
    .io_right_out_ready(cols_7_13_io_right_out_ready),
    .io_right_out_valid(cols_7_13_io_right_out_valid),
    .io_right_out_bits(cols_7_13_io_right_out_bits),
    .io_bottom_out_ready(cols_7_13_io_bottom_out_ready),
    .io_bottom_out_valid(cols_7_13_io_bottom_out_valid),
    .io_bottom_out_bits(cols_7_13_io_bottom_out_bits)
  );
  ProcessingElement cols_8_13 ( // @[Stab.scala 85:60]
    .clock(cols_8_13_clock),
    .reset(cols_8_13_reset),
    .io_left_in_ready(cols_8_13_io_left_in_ready),
    .io_left_in_valid(cols_8_13_io_left_in_valid),
    .io_left_in_bits(cols_8_13_io_left_in_bits),
    .io_top_in_ready(cols_8_13_io_top_in_ready),
    .io_top_in_valid(cols_8_13_io_top_in_valid),
    .io_top_in_bits(cols_8_13_io_top_in_bits),
    .io_sum_ready(cols_8_13_io_sum_ready),
    .io_sum_valid(cols_8_13_io_sum_valid),
    .io_sum_bits(cols_8_13_io_sum_bits),
    .io_right_out_ready(cols_8_13_io_right_out_ready),
    .io_right_out_valid(cols_8_13_io_right_out_valid),
    .io_right_out_bits(cols_8_13_io_right_out_bits),
    .io_bottom_out_ready(cols_8_13_io_bottom_out_ready),
    .io_bottom_out_valid(cols_8_13_io_bottom_out_valid),
    .io_bottom_out_bits(cols_8_13_io_bottom_out_bits)
  );
  ProcessingElement cols_9_13 ( // @[Stab.scala 85:60]
    .clock(cols_9_13_clock),
    .reset(cols_9_13_reset),
    .io_left_in_ready(cols_9_13_io_left_in_ready),
    .io_left_in_valid(cols_9_13_io_left_in_valid),
    .io_left_in_bits(cols_9_13_io_left_in_bits),
    .io_top_in_ready(cols_9_13_io_top_in_ready),
    .io_top_in_valid(cols_9_13_io_top_in_valid),
    .io_top_in_bits(cols_9_13_io_top_in_bits),
    .io_sum_ready(cols_9_13_io_sum_ready),
    .io_sum_valid(cols_9_13_io_sum_valid),
    .io_sum_bits(cols_9_13_io_sum_bits),
    .io_right_out_ready(cols_9_13_io_right_out_ready),
    .io_right_out_valid(cols_9_13_io_right_out_valid),
    .io_right_out_bits(cols_9_13_io_right_out_bits),
    .io_bottom_out_ready(cols_9_13_io_bottom_out_ready),
    .io_bottom_out_valid(cols_9_13_io_bottom_out_valid),
    .io_bottom_out_bits(cols_9_13_io_bottom_out_bits)
  );
  ProcessingElement cols_10_13 ( // @[Stab.scala 85:60]
    .clock(cols_10_13_clock),
    .reset(cols_10_13_reset),
    .io_left_in_ready(cols_10_13_io_left_in_ready),
    .io_left_in_valid(cols_10_13_io_left_in_valid),
    .io_left_in_bits(cols_10_13_io_left_in_bits),
    .io_top_in_ready(cols_10_13_io_top_in_ready),
    .io_top_in_valid(cols_10_13_io_top_in_valid),
    .io_top_in_bits(cols_10_13_io_top_in_bits),
    .io_sum_ready(cols_10_13_io_sum_ready),
    .io_sum_valid(cols_10_13_io_sum_valid),
    .io_sum_bits(cols_10_13_io_sum_bits),
    .io_right_out_ready(cols_10_13_io_right_out_ready),
    .io_right_out_valid(cols_10_13_io_right_out_valid),
    .io_right_out_bits(cols_10_13_io_right_out_bits),
    .io_bottom_out_ready(cols_10_13_io_bottom_out_ready),
    .io_bottom_out_valid(cols_10_13_io_bottom_out_valid),
    .io_bottom_out_bits(cols_10_13_io_bottom_out_bits)
  );
  ProcessingElement cols_11_13 ( // @[Stab.scala 85:60]
    .clock(cols_11_13_clock),
    .reset(cols_11_13_reset),
    .io_left_in_ready(cols_11_13_io_left_in_ready),
    .io_left_in_valid(cols_11_13_io_left_in_valid),
    .io_left_in_bits(cols_11_13_io_left_in_bits),
    .io_top_in_ready(cols_11_13_io_top_in_ready),
    .io_top_in_valid(cols_11_13_io_top_in_valid),
    .io_top_in_bits(cols_11_13_io_top_in_bits),
    .io_sum_ready(cols_11_13_io_sum_ready),
    .io_sum_valid(cols_11_13_io_sum_valid),
    .io_sum_bits(cols_11_13_io_sum_bits),
    .io_right_out_ready(cols_11_13_io_right_out_ready),
    .io_right_out_valid(cols_11_13_io_right_out_valid),
    .io_right_out_bits(cols_11_13_io_right_out_bits),
    .io_bottom_out_ready(cols_11_13_io_bottom_out_ready),
    .io_bottom_out_valid(cols_11_13_io_bottom_out_valid),
    .io_bottom_out_bits(cols_11_13_io_bottom_out_bits)
  );
  ProcessingElement cols_12_13 ( // @[Stab.scala 85:60]
    .clock(cols_12_13_clock),
    .reset(cols_12_13_reset),
    .io_left_in_ready(cols_12_13_io_left_in_ready),
    .io_left_in_valid(cols_12_13_io_left_in_valid),
    .io_left_in_bits(cols_12_13_io_left_in_bits),
    .io_top_in_ready(cols_12_13_io_top_in_ready),
    .io_top_in_valid(cols_12_13_io_top_in_valid),
    .io_top_in_bits(cols_12_13_io_top_in_bits),
    .io_sum_ready(cols_12_13_io_sum_ready),
    .io_sum_valid(cols_12_13_io_sum_valid),
    .io_sum_bits(cols_12_13_io_sum_bits),
    .io_right_out_ready(cols_12_13_io_right_out_ready),
    .io_right_out_valid(cols_12_13_io_right_out_valid),
    .io_right_out_bits(cols_12_13_io_right_out_bits),
    .io_bottom_out_ready(cols_12_13_io_bottom_out_ready),
    .io_bottom_out_valid(cols_12_13_io_bottom_out_valid),
    .io_bottom_out_bits(cols_12_13_io_bottom_out_bits)
  );
  ProcessingElement cols_13_13 ( // @[Stab.scala 85:60]
    .clock(cols_13_13_clock),
    .reset(cols_13_13_reset),
    .io_left_in_ready(cols_13_13_io_left_in_ready),
    .io_left_in_valid(cols_13_13_io_left_in_valid),
    .io_left_in_bits(cols_13_13_io_left_in_bits),
    .io_top_in_ready(cols_13_13_io_top_in_ready),
    .io_top_in_valid(cols_13_13_io_top_in_valid),
    .io_top_in_bits(cols_13_13_io_top_in_bits),
    .io_sum_ready(cols_13_13_io_sum_ready),
    .io_sum_valid(cols_13_13_io_sum_valid),
    .io_sum_bits(cols_13_13_io_sum_bits),
    .io_right_out_ready(cols_13_13_io_right_out_ready),
    .io_right_out_valid(cols_13_13_io_right_out_valid),
    .io_right_out_bits(cols_13_13_io_right_out_bits),
    .io_bottom_out_ready(cols_13_13_io_bottom_out_ready),
    .io_bottom_out_valid(cols_13_13_io_bottom_out_valid),
    .io_bottom_out_bits(cols_13_13_io_bottom_out_bits)
  );
  ProcessingElement cols_14_13 ( // @[Stab.scala 85:60]
    .clock(cols_14_13_clock),
    .reset(cols_14_13_reset),
    .io_left_in_ready(cols_14_13_io_left_in_ready),
    .io_left_in_valid(cols_14_13_io_left_in_valid),
    .io_left_in_bits(cols_14_13_io_left_in_bits),
    .io_top_in_ready(cols_14_13_io_top_in_ready),
    .io_top_in_valid(cols_14_13_io_top_in_valid),
    .io_top_in_bits(cols_14_13_io_top_in_bits),
    .io_sum_ready(cols_14_13_io_sum_ready),
    .io_sum_valid(cols_14_13_io_sum_valid),
    .io_sum_bits(cols_14_13_io_sum_bits),
    .io_right_out_ready(cols_14_13_io_right_out_ready),
    .io_right_out_valid(cols_14_13_io_right_out_valid),
    .io_right_out_bits(cols_14_13_io_right_out_bits),
    .io_bottom_out_ready(cols_14_13_io_bottom_out_ready),
    .io_bottom_out_valid(cols_14_13_io_bottom_out_valid),
    .io_bottom_out_bits(cols_14_13_io_bottom_out_bits)
  );
  ProcessingElement cols_15_13 ( // @[Stab.scala 85:60]
    .clock(cols_15_13_clock),
    .reset(cols_15_13_reset),
    .io_left_in_ready(cols_15_13_io_left_in_ready),
    .io_left_in_valid(cols_15_13_io_left_in_valid),
    .io_left_in_bits(cols_15_13_io_left_in_bits),
    .io_top_in_ready(cols_15_13_io_top_in_ready),
    .io_top_in_valid(cols_15_13_io_top_in_valid),
    .io_top_in_bits(cols_15_13_io_top_in_bits),
    .io_sum_ready(cols_15_13_io_sum_ready),
    .io_sum_valid(cols_15_13_io_sum_valid),
    .io_sum_bits(cols_15_13_io_sum_bits),
    .io_right_out_ready(cols_15_13_io_right_out_ready),
    .io_right_out_valid(cols_15_13_io_right_out_valid),
    .io_right_out_bits(cols_15_13_io_right_out_bits),
    .io_bottom_out_ready(cols_15_13_io_bottom_out_ready),
    .io_bottom_out_valid(cols_15_13_io_bottom_out_valid),
    .io_bottom_out_bits(cols_15_13_io_bottom_out_bits)
  );
  ProcessingElement cols_0_14 ( // @[Stab.scala 85:60]
    .clock(cols_0_14_clock),
    .reset(cols_0_14_reset),
    .io_left_in_ready(cols_0_14_io_left_in_ready),
    .io_left_in_valid(cols_0_14_io_left_in_valid),
    .io_left_in_bits(cols_0_14_io_left_in_bits),
    .io_top_in_ready(cols_0_14_io_top_in_ready),
    .io_top_in_valid(cols_0_14_io_top_in_valid),
    .io_top_in_bits(cols_0_14_io_top_in_bits),
    .io_sum_ready(cols_0_14_io_sum_ready),
    .io_sum_valid(cols_0_14_io_sum_valid),
    .io_sum_bits(cols_0_14_io_sum_bits),
    .io_right_out_ready(cols_0_14_io_right_out_ready),
    .io_right_out_valid(cols_0_14_io_right_out_valid),
    .io_right_out_bits(cols_0_14_io_right_out_bits),
    .io_bottom_out_ready(cols_0_14_io_bottom_out_ready),
    .io_bottom_out_valid(cols_0_14_io_bottom_out_valid),
    .io_bottom_out_bits(cols_0_14_io_bottom_out_bits)
  );
  ProcessingElement cols_1_14 ( // @[Stab.scala 85:60]
    .clock(cols_1_14_clock),
    .reset(cols_1_14_reset),
    .io_left_in_ready(cols_1_14_io_left_in_ready),
    .io_left_in_valid(cols_1_14_io_left_in_valid),
    .io_left_in_bits(cols_1_14_io_left_in_bits),
    .io_top_in_ready(cols_1_14_io_top_in_ready),
    .io_top_in_valid(cols_1_14_io_top_in_valid),
    .io_top_in_bits(cols_1_14_io_top_in_bits),
    .io_sum_ready(cols_1_14_io_sum_ready),
    .io_sum_valid(cols_1_14_io_sum_valid),
    .io_sum_bits(cols_1_14_io_sum_bits),
    .io_right_out_ready(cols_1_14_io_right_out_ready),
    .io_right_out_valid(cols_1_14_io_right_out_valid),
    .io_right_out_bits(cols_1_14_io_right_out_bits),
    .io_bottom_out_ready(cols_1_14_io_bottom_out_ready),
    .io_bottom_out_valid(cols_1_14_io_bottom_out_valid),
    .io_bottom_out_bits(cols_1_14_io_bottom_out_bits)
  );
  ProcessingElement cols_2_14 ( // @[Stab.scala 85:60]
    .clock(cols_2_14_clock),
    .reset(cols_2_14_reset),
    .io_left_in_ready(cols_2_14_io_left_in_ready),
    .io_left_in_valid(cols_2_14_io_left_in_valid),
    .io_left_in_bits(cols_2_14_io_left_in_bits),
    .io_top_in_ready(cols_2_14_io_top_in_ready),
    .io_top_in_valid(cols_2_14_io_top_in_valid),
    .io_top_in_bits(cols_2_14_io_top_in_bits),
    .io_sum_ready(cols_2_14_io_sum_ready),
    .io_sum_valid(cols_2_14_io_sum_valid),
    .io_sum_bits(cols_2_14_io_sum_bits),
    .io_right_out_ready(cols_2_14_io_right_out_ready),
    .io_right_out_valid(cols_2_14_io_right_out_valid),
    .io_right_out_bits(cols_2_14_io_right_out_bits),
    .io_bottom_out_ready(cols_2_14_io_bottom_out_ready),
    .io_bottom_out_valid(cols_2_14_io_bottom_out_valid),
    .io_bottom_out_bits(cols_2_14_io_bottom_out_bits)
  );
  ProcessingElement cols_3_14 ( // @[Stab.scala 85:60]
    .clock(cols_3_14_clock),
    .reset(cols_3_14_reset),
    .io_left_in_ready(cols_3_14_io_left_in_ready),
    .io_left_in_valid(cols_3_14_io_left_in_valid),
    .io_left_in_bits(cols_3_14_io_left_in_bits),
    .io_top_in_ready(cols_3_14_io_top_in_ready),
    .io_top_in_valid(cols_3_14_io_top_in_valid),
    .io_top_in_bits(cols_3_14_io_top_in_bits),
    .io_sum_ready(cols_3_14_io_sum_ready),
    .io_sum_valid(cols_3_14_io_sum_valid),
    .io_sum_bits(cols_3_14_io_sum_bits),
    .io_right_out_ready(cols_3_14_io_right_out_ready),
    .io_right_out_valid(cols_3_14_io_right_out_valid),
    .io_right_out_bits(cols_3_14_io_right_out_bits),
    .io_bottom_out_ready(cols_3_14_io_bottom_out_ready),
    .io_bottom_out_valid(cols_3_14_io_bottom_out_valid),
    .io_bottom_out_bits(cols_3_14_io_bottom_out_bits)
  );
  ProcessingElement cols_4_14 ( // @[Stab.scala 85:60]
    .clock(cols_4_14_clock),
    .reset(cols_4_14_reset),
    .io_left_in_ready(cols_4_14_io_left_in_ready),
    .io_left_in_valid(cols_4_14_io_left_in_valid),
    .io_left_in_bits(cols_4_14_io_left_in_bits),
    .io_top_in_ready(cols_4_14_io_top_in_ready),
    .io_top_in_valid(cols_4_14_io_top_in_valid),
    .io_top_in_bits(cols_4_14_io_top_in_bits),
    .io_sum_ready(cols_4_14_io_sum_ready),
    .io_sum_valid(cols_4_14_io_sum_valid),
    .io_sum_bits(cols_4_14_io_sum_bits),
    .io_right_out_ready(cols_4_14_io_right_out_ready),
    .io_right_out_valid(cols_4_14_io_right_out_valid),
    .io_right_out_bits(cols_4_14_io_right_out_bits),
    .io_bottom_out_ready(cols_4_14_io_bottom_out_ready),
    .io_bottom_out_valid(cols_4_14_io_bottom_out_valid),
    .io_bottom_out_bits(cols_4_14_io_bottom_out_bits)
  );
  ProcessingElement cols_5_14 ( // @[Stab.scala 85:60]
    .clock(cols_5_14_clock),
    .reset(cols_5_14_reset),
    .io_left_in_ready(cols_5_14_io_left_in_ready),
    .io_left_in_valid(cols_5_14_io_left_in_valid),
    .io_left_in_bits(cols_5_14_io_left_in_bits),
    .io_top_in_ready(cols_5_14_io_top_in_ready),
    .io_top_in_valid(cols_5_14_io_top_in_valid),
    .io_top_in_bits(cols_5_14_io_top_in_bits),
    .io_sum_ready(cols_5_14_io_sum_ready),
    .io_sum_valid(cols_5_14_io_sum_valid),
    .io_sum_bits(cols_5_14_io_sum_bits),
    .io_right_out_ready(cols_5_14_io_right_out_ready),
    .io_right_out_valid(cols_5_14_io_right_out_valid),
    .io_right_out_bits(cols_5_14_io_right_out_bits),
    .io_bottom_out_ready(cols_5_14_io_bottom_out_ready),
    .io_bottom_out_valid(cols_5_14_io_bottom_out_valid),
    .io_bottom_out_bits(cols_5_14_io_bottom_out_bits)
  );
  ProcessingElement cols_6_14 ( // @[Stab.scala 85:60]
    .clock(cols_6_14_clock),
    .reset(cols_6_14_reset),
    .io_left_in_ready(cols_6_14_io_left_in_ready),
    .io_left_in_valid(cols_6_14_io_left_in_valid),
    .io_left_in_bits(cols_6_14_io_left_in_bits),
    .io_top_in_ready(cols_6_14_io_top_in_ready),
    .io_top_in_valid(cols_6_14_io_top_in_valid),
    .io_top_in_bits(cols_6_14_io_top_in_bits),
    .io_sum_ready(cols_6_14_io_sum_ready),
    .io_sum_valid(cols_6_14_io_sum_valid),
    .io_sum_bits(cols_6_14_io_sum_bits),
    .io_right_out_ready(cols_6_14_io_right_out_ready),
    .io_right_out_valid(cols_6_14_io_right_out_valid),
    .io_right_out_bits(cols_6_14_io_right_out_bits),
    .io_bottom_out_ready(cols_6_14_io_bottom_out_ready),
    .io_bottom_out_valid(cols_6_14_io_bottom_out_valid),
    .io_bottom_out_bits(cols_6_14_io_bottom_out_bits)
  );
  ProcessingElement cols_7_14 ( // @[Stab.scala 85:60]
    .clock(cols_7_14_clock),
    .reset(cols_7_14_reset),
    .io_left_in_ready(cols_7_14_io_left_in_ready),
    .io_left_in_valid(cols_7_14_io_left_in_valid),
    .io_left_in_bits(cols_7_14_io_left_in_bits),
    .io_top_in_ready(cols_7_14_io_top_in_ready),
    .io_top_in_valid(cols_7_14_io_top_in_valid),
    .io_top_in_bits(cols_7_14_io_top_in_bits),
    .io_sum_ready(cols_7_14_io_sum_ready),
    .io_sum_valid(cols_7_14_io_sum_valid),
    .io_sum_bits(cols_7_14_io_sum_bits),
    .io_right_out_ready(cols_7_14_io_right_out_ready),
    .io_right_out_valid(cols_7_14_io_right_out_valid),
    .io_right_out_bits(cols_7_14_io_right_out_bits),
    .io_bottom_out_ready(cols_7_14_io_bottom_out_ready),
    .io_bottom_out_valid(cols_7_14_io_bottom_out_valid),
    .io_bottom_out_bits(cols_7_14_io_bottom_out_bits)
  );
  ProcessingElement cols_8_14 ( // @[Stab.scala 85:60]
    .clock(cols_8_14_clock),
    .reset(cols_8_14_reset),
    .io_left_in_ready(cols_8_14_io_left_in_ready),
    .io_left_in_valid(cols_8_14_io_left_in_valid),
    .io_left_in_bits(cols_8_14_io_left_in_bits),
    .io_top_in_ready(cols_8_14_io_top_in_ready),
    .io_top_in_valid(cols_8_14_io_top_in_valid),
    .io_top_in_bits(cols_8_14_io_top_in_bits),
    .io_sum_ready(cols_8_14_io_sum_ready),
    .io_sum_valid(cols_8_14_io_sum_valid),
    .io_sum_bits(cols_8_14_io_sum_bits),
    .io_right_out_ready(cols_8_14_io_right_out_ready),
    .io_right_out_valid(cols_8_14_io_right_out_valid),
    .io_right_out_bits(cols_8_14_io_right_out_bits),
    .io_bottom_out_ready(cols_8_14_io_bottom_out_ready),
    .io_bottom_out_valid(cols_8_14_io_bottom_out_valid),
    .io_bottom_out_bits(cols_8_14_io_bottom_out_bits)
  );
  ProcessingElement cols_9_14 ( // @[Stab.scala 85:60]
    .clock(cols_9_14_clock),
    .reset(cols_9_14_reset),
    .io_left_in_ready(cols_9_14_io_left_in_ready),
    .io_left_in_valid(cols_9_14_io_left_in_valid),
    .io_left_in_bits(cols_9_14_io_left_in_bits),
    .io_top_in_ready(cols_9_14_io_top_in_ready),
    .io_top_in_valid(cols_9_14_io_top_in_valid),
    .io_top_in_bits(cols_9_14_io_top_in_bits),
    .io_sum_ready(cols_9_14_io_sum_ready),
    .io_sum_valid(cols_9_14_io_sum_valid),
    .io_sum_bits(cols_9_14_io_sum_bits),
    .io_right_out_ready(cols_9_14_io_right_out_ready),
    .io_right_out_valid(cols_9_14_io_right_out_valid),
    .io_right_out_bits(cols_9_14_io_right_out_bits),
    .io_bottom_out_ready(cols_9_14_io_bottom_out_ready),
    .io_bottom_out_valid(cols_9_14_io_bottom_out_valid),
    .io_bottom_out_bits(cols_9_14_io_bottom_out_bits)
  );
  ProcessingElement cols_10_14 ( // @[Stab.scala 85:60]
    .clock(cols_10_14_clock),
    .reset(cols_10_14_reset),
    .io_left_in_ready(cols_10_14_io_left_in_ready),
    .io_left_in_valid(cols_10_14_io_left_in_valid),
    .io_left_in_bits(cols_10_14_io_left_in_bits),
    .io_top_in_ready(cols_10_14_io_top_in_ready),
    .io_top_in_valid(cols_10_14_io_top_in_valid),
    .io_top_in_bits(cols_10_14_io_top_in_bits),
    .io_sum_ready(cols_10_14_io_sum_ready),
    .io_sum_valid(cols_10_14_io_sum_valid),
    .io_sum_bits(cols_10_14_io_sum_bits),
    .io_right_out_ready(cols_10_14_io_right_out_ready),
    .io_right_out_valid(cols_10_14_io_right_out_valid),
    .io_right_out_bits(cols_10_14_io_right_out_bits),
    .io_bottom_out_ready(cols_10_14_io_bottom_out_ready),
    .io_bottom_out_valid(cols_10_14_io_bottom_out_valid),
    .io_bottom_out_bits(cols_10_14_io_bottom_out_bits)
  );
  ProcessingElement cols_11_14 ( // @[Stab.scala 85:60]
    .clock(cols_11_14_clock),
    .reset(cols_11_14_reset),
    .io_left_in_ready(cols_11_14_io_left_in_ready),
    .io_left_in_valid(cols_11_14_io_left_in_valid),
    .io_left_in_bits(cols_11_14_io_left_in_bits),
    .io_top_in_ready(cols_11_14_io_top_in_ready),
    .io_top_in_valid(cols_11_14_io_top_in_valid),
    .io_top_in_bits(cols_11_14_io_top_in_bits),
    .io_sum_ready(cols_11_14_io_sum_ready),
    .io_sum_valid(cols_11_14_io_sum_valid),
    .io_sum_bits(cols_11_14_io_sum_bits),
    .io_right_out_ready(cols_11_14_io_right_out_ready),
    .io_right_out_valid(cols_11_14_io_right_out_valid),
    .io_right_out_bits(cols_11_14_io_right_out_bits),
    .io_bottom_out_ready(cols_11_14_io_bottom_out_ready),
    .io_bottom_out_valid(cols_11_14_io_bottom_out_valid),
    .io_bottom_out_bits(cols_11_14_io_bottom_out_bits)
  );
  ProcessingElement cols_12_14 ( // @[Stab.scala 85:60]
    .clock(cols_12_14_clock),
    .reset(cols_12_14_reset),
    .io_left_in_ready(cols_12_14_io_left_in_ready),
    .io_left_in_valid(cols_12_14_io_left_in_valid),
    .io_left_in_bits(cols_12_14_io_left_in_bits),
    .io_top_in_ready(cols_12_14_io_top_in_ready),
    .io_top_in_valid(cols_12_14_io_top_in_valid),
    .io_top_in_bits(cols_12_14_io_top_in_bits),
    .io_sum_ready(cols_12_14_io_sum_ready),
    .io_sum_valid(cols_12_14_io_sum_valid),
    .io_sum_bits(cols_12_14_io_sum_bits),
    .io_right_out_ready(cols_12_14_io_right_out_ready),
    .io_right_out_valid(cols_12_14_io_right_out_valid),
    .io_right_out_bits(cols_12_14_io_right_out_bits),
    .io_bottom_out_ready(cols_12_14_io_bottom_out_ready),
    .io_bottom_out_valid(cols_12_14_io_bottom_out_valid),
    .io_bottom_out_bits(cols_12_14_io_bottom_out_bits)
  );
  ProcessingElement cols_13_14 ( // @[Stab.scala 85:60]
    .clock(cols_13_14_clock),
    .reset(cols_13_14_reset),
    .io_left_in_ready(cols_13_14_io_left_in_ready),
    .io_left_in_valid(cols_13_14_io_left_in_valid),
    .io_left_in_bits(cols_13_14_io_left_in_bits),
    .io_top_in_ready(cols_13_14_io_top_in_ready),
    .io_top_in_valid(cols_13_14_io_top_in_valid),
    .io_top_in_bits(cols_13_14_io_top_in_bits),
    .io_sum_ready(cols_13_14_io_sum_ready),
    .io_sum_valid(cols_13_14_io_sum_valid),
    .io_sum_bits(cols_13_14_io_sum_bits),
    .io_right_out_ready(cols_13_14_io_right_out_ready),
    .io_right_out_valid(cols_13_14_io_right_out_valid),
    .io_right_out_bits(cols_13_14_io_right_out_bits),
    .io_bottom_out_ready(cols_13_14_io_bottom_out_ready),
    .io_bottom_out_valid(cols_13_14_io_bottom_out_valid),
    .io_bottom_out_bits(cols_13_14_io_bottom_out_bits)
  );
  ProcessingElement cols_14_14 ( // @[Stab.scala 85:60]
    .clock(cols_14_14_clock),
    .reset(cols_14_14_reset),
    .io_left_in_ready(cols_14_14_io_left_in_ready),
    .io_left_in_valid(cols_14_14_io_left_in_valid),
    .io_left_in_bits(cols_14_14_io_left_in_bits),
    .io_top_in_ready(cols_14_14_io_top_in_ready),
    .io_top_in_valid(cols_14_14_io_top_in_valid),
    .io_top_in_bits(cols_14_14_io_top_in_bits),
    .io_sum_ready(cols_14_14_io_sum_ready),
    .io_sum_valid(cols_14_14_io_sum_valid),
    .io_sum_bits(cols_14_14_io_sum_bits),
    .io_right_out_ready(cols_14_14_io_right_out_ready),
    .io_right_out_valid(cols_14_14_io_right_out_valid),
    .io_right_out_bits(cols_14_14_io_right_out_bits),
    .io_bottom_out_ready(cols_14_14_io_bottom_out_ready),
    .io_bottom_out_valid(cols_14_14_io_bottom_out_valid),
    .io_bottom_out_bits(cols_14_14_io_bottom_out_bits)
  );
  ProcessingElement cols_15_14 ( // @[Stab.scala 85:60]
    .clock(cols_15_14_clock),
    .reset(cols_15_14_reset),
    .io_left_in_ready(cols_15_14_io_left_in_ready),
    .io_left_in_valid(cols_15_14_io_left_in_valid),
    .io_left_in_bits(cols_15_14_io_left_in_bits),
    .io_top_in_ready(cols_15_14_io_top_in_ready),
    .io_top_in_valid(cols_15_14_io_top_in_valid),
    .io_top_in_bits(cols_15_14_io_top_in_bits),
    .io_sum_ready(cols_15_14_io_sum_ready),
    .io_sum_valid(cols_15_14_io_sum_valid),
    .io_sum_bits(cols_15_14_io_sum_bits),
    .io_right_out_ready(cols_15_14_io_right_out_ready),
    .io_right_out_valid(cols_15_14_io_right_out_valid),
    .io_right_out_bits(cols_15_14_io_right_out_bits),
    .io_bottom_out_ready(cols_15_14_io_bottom_out_ready),
    .io_bottom_out_valid(cols_15_14_io_bottom_out_valid),
    .io_bottom_out_bits(cols_15_14_io_bottom_out_bits)
  );
  ProcessingElement cols_0_15 ( // @[Stab.scala 85:60]
    .clock(cols_0_15_clock),
    .reset(cols_0_15_reset),
    .io_left_in_ready(cols_0_15_io_left_in_ready),
    .io_left_in_valid(cols_0_15_io_left_in_valid),
    .io_left_in_bits(cols_0_15_io_left_in_bits),
    .io_top_in_ready(cols_0_15_io_top_in_ready),
    .io_top_in_valid(cols_0_15_io_top_in_valid),
    .io_top_in_bits(cols_0_15_io_top_in_bits),
    .io_sum_ready(cols_0_15_io_sum_ready),
    .io_sum_valid(cols_0_15_io_sum_valid),
    .io_sum_bits(cols_0_15_io_sum_bits),
    .io_right_out_ready(cols_0_15_io_right_out_ready),
    .io_right_out_valid(cols_0_15_io_right_out_valid),
    .io_right_out_bits(cols_0_15_io_right_out_bits),
    .io_bottom_out_ready(cols_0_15_io_bottom_out_ready),
    .io_bottom_out_valid(cols_0_15_io_bottom_out_valid),
    .io_bottom_out_bits(cols_0_15_io_bottom_out_bits)
  );
  ProcessingElement cols_1_15 ( // @[Stab.scala 85:60]
    .clock(cols_1_15_clock),
    .reset(cols_1_15_reset),
    .io_left_in_ready(cols_1_15_io_left_in_ready),
    .io_left_in_valid(cols_1_15_io_left_in_valid),
    .io_left_in_bits(cols_1_15_io_left_in_bits),
    .io_top_in_ready(cols_1_15_io_top_in_ready),
    .io_top_in_valid(cols_1_15_io_top_in_valid),
    .io_top_in_bits(cols_1_15_io_top_in_bits),
    .io_sum_ready(cols_1_15_io_sum_ready),
    .io_sum_valid(cols_1_15_io_sum_valid),
    .io_sum_bits(cols_1_15_io_sum_bits),
    .io_right_out_ready(cols_1_15_io_right_out_ready),
    .io_right_out_valid(cols_1_15_io_right_out_valid),
    .io_right_out_bits(cols_1_15_io_right_out_bits),
    .io_bottom_out_ready(cols_1_15_io_bottom_out_ready),
    .io_bottom_out_valid(cols_1_15_io_bottom_out_valid),
    .io_bottom_out_bits(cols_1_15_io_bottom_out_bits)
  );
  ProcessingElement cols_2_15 ( // @[Stab.scala 85:60]
    .clock(cols_2_15_clock),
    .reset(cols_2_15_reset),
    .io_left_in_ready(cols_2_15_io_left_in_ready),
    .io_left_in_valid(cols_2_15_io_left_in_valid),
    .io_left_in_bits(cols_2_15_io_left_in_bits),
    .io_top_in_ready(cols_2_15_io_top_in_ready),
    .io_top_in_valid(cols_2_15_io_top_in_valid),
    .io_top_in_bits(cols_2_15_io_top_in_bits),
    .io_sum_ready(cols_2_15_io_sum_ready),
    .io_sum_valid(cols_2_15_io_sum_valid),
    .io_sum_bits(cols_2_15_io_sum_bits),
    .io_right_out_ready(cols_2_15_io_right_out_ready),
    .io_right_out_valid(cols_2_15_io_right_out_valid),
    .io_right_out_bits(cols_2_15_io_right_out_bits),
    .io_bottom_out_ready(cols_2_15_io_bottom_out_ready),
    .io_bottom_out_valid(cols_2_15_io_bottom_out_valid),
    .io_bottom_out_bits(cols_2_15_io_bottom_out_bits)
  );
  ProcessingElement cols_3_15 ( // @[Stab.scala 85:60]
    .clock(cols_3_15_clock),
    .reset(cols_3_15_reset),
    .io_left_in_ready(cols_3_15_io_left_in_ready),
    .io_left_in_valid(cols_3_15_io_left_in_valid),
    .io_left_in_bits(cols_3_15_io_left_in_bits),
    .io_top_in_ready(cols_3_15_io_top_in_ready),
    .io_top_in_valid(cols_3_15_io_top_in_valid),
    .io_top_in_bits(cols_3_15_io_top_in_bits),
    .io_sum_ready(cols_3_15_io_sum_ready),
    .io_sum_valid(cols_3_15_io_sum_valid),
    .io_sum_bits(cols_3_15_io_sum_bits),
    .io_right_out_ready(cols_3_15_io_right_out_ready),
    .io_right_out_valid(cols_3_15_io_right_out_valid),
    .io_right_out_bits(cols_3_15_io_right_out_bits),
    .io_bottom_out_ready(cols_3_15_io_bottom_out_ready),
    .io_bottom_out_valid(cols_3_15_io_bottom_out_valid),
    .io_bottom_out_bits(cols_3_15_io_bottom_out_bits)
  );
  ProcessingElement cols_4_15 ( // @[Stab.scala 85:60]
    .clock(cols_4_15_clock),
    .reset(cols_4_15_reset),
    .io_left_in_ready(cols_4_15_io_left_in_ready),
    .io_left_in_valid(cols_4_15_io_left_in_valid),
    .io_left_in_bits(cols_4_15_io_left_in_bits),
    .io_top_in_ready(cols_4_15_io_top_in_ready),
    .io_top_in_valid(cols_4_15_io_top_in_valid),
    .io_top_in_bits(cols_4_15_io_top_in_bits),
    .io_sum_ready(cols_4_15_io_sum_ready),
    .io_sum_valid(cols_4_15_io_sum_valid),
    .io_sum_bits(cols_4_15_io_sum_bits),
    .io_right_out_ready(cols_4_15_io_right_out_ready),
    .io_right_out_valid(cols_4_15_io_right_out_valid),
    .io_right_out_bits(cols_4_15_io_right_out_bits),
    .io_bottom_out_ready(cols_4_15_io_bottom_out_ready),
    .io_bottom_out_valid(cols_4_15_io_bottom_out_valid),
    .io_bottom_out_bits(cols_4_15_io_bottom_out_bits)
  );
  ProcessingElement cols_5_15 ( // @[Stab.scala 85:60]
    .clock(cols_5_15_clock),
    .reset(cols_5_15_reset),
    .io_left_in_ready(cols_5_15_io_left_in_ready),
    .io_left_in_valid(cols_5_15_io_left_in_valid),
    .io_left_in_bits(cols_5_15_io_left_in_bits),
    .io_top_in_ready(cols_5_15_io_top_in_ready),
    .io_top_in_valid(cols_5_15_io_top_in_valid),
    .io_top_in_bits(cols_5_15_io_top_in_bits),
    .io_sum_ready(cols_5_15_io_sum_ready),
    .io_sum_valid(cols_5_15_io_sum_valid),
    .io_sum_bits(cols_5_15_io_sum_bits),
    .io_right_out_ready(cols_5_15_io_right_out_ready),
    .io_right_out_valid(cols_5_15_io_right_out_valid),
    .io_right_out_bits(cols_5_15_io_right_out_bits),
    .io_bottom_out_ready(cols_5_15_io_bottom_out_ready),
    .io_bottom_out_valid(cols_5_15_io_bottom_out_valid),
    .io_bottom_out_bits(cols_5_15_io_bottom_out_bits)
  );
  ProcessingElement cols_6_15 ( // @[Stab.scala 85:60]
    .clock(cols_6_15_clock),
    .reset(cols_6_15_reset),
    .io_left_in_ready(cols_6_15_io_left_in_ready),
    .io_left_in_valid(cols_6_15_io_left_in_valid),
    .io_left_in_bits(cols_6_15_io_left_in_bits),
    .io_top_in_ready(cols_6_15_io_top_in_ready),
    .io_top_in_valid(cols_6_15_io_top_in_valid),
    .io_top_in_bits(cols_6_15_io_top_in_bits),
    .io_sum_ready(cols_6_15_io_sum_ready),
    .io_sum_valid(cols_6_15_io_sum_valid),
    .io_sum_bits(cols_6_15_io_sum_bits),
    .io_right_out_ready(cols_6_15_io_right_out_ready),
    .io_right_out_valid(cols_6_15_io_right_out_valid),
    .io_right_out_bits(cols_6_15_io_right_out_bits),
    .io_bottom_out_ready(cols_6_15_io_bottom_out_ready),
    .io_bottom_out_valid(cols_6_15_io_bottom_out_valid),
    .io_bottom_out_bits(cols_6_15_io_bottom_out_bits)
  );
  ProcessingElement cols_7_15 ( // @[Stab.scala 85:60]
    .clock(cols_7_15_clock),
    .reset(cols_7_15_reset),
    .io_left_in_ready(cols_7_15_io_left_in_ready),
    .io_left_in_valid(cols_7_15_io_left_in_valid),
    .io_left_in_bits(cols_7_15_io_left_in_bits),
    .io_top_in_ready(cols_7_15_io_top_in_ready),
    .io_top_in_valid(cols_7_15_io_top_in_valid),
    .io_top_in_bits(cols_7_15_io_top_in_bits),
    .io_sum_ready(cols_7_15_io_sum_ready),
    .io_sum_valid(cols_7_15_io_sum_valid),
    .io_sum_bits(cols_7_15_io_sum_bits),
    .io_right_out_ready(cols_7_15_io_right_out_ready),
    .io_right_out_valid(cols_7_15_io_right_out_valid),
    .io_right_out_bits(cols_7_15_io_right_out_bits),
    .io_bottom_out_ready(cols_7_15_io_bottom_out_ready),
    .io_bottom_out_valid(cols_7_15_io_bottom_out_valid),
    .io_bottom_out_bits(cols_7_15_io_bottom_out_bits)
  );
  ProcessingElement cols_8_15 ( // @[Stab.scala 85:60]
    .clock(cols_8_15_clock),
    .reset(cols_8_15_reset),
    .io_left_in_ready(cols_8_15_io_left_in_ready),
    .io_left_in_valid(cols_8_15_io_left_in_valid),
    .io_left_in_bits(cols_8_15_io_left_in_bits),
    .io_top_in_ready(cols_8_15_io_top_in_ready),
    .io_top_in_valid(cols_8_15_io_top_in_valid),
    .io_top_in_bits(cols_8_15_io_top_in_bits),
    .io_sum_ready(cols_8_15_io_sum_ready),
    .io_sum_valid(cols_8_15_io_sum_valid),
    .io_sum_bits(cols_8_15_io_sum_bits),
    .io_right_out_ready(cols_8_15_io_right_out_ready),
    .io_right_out_valid(cols_8_15_io_right_out_valid),
    .io_right_out_bits(cols_8_15_io_right_out_bits),
    .io_bottom_out_ready(cols_8_15_io_bottom_out_ready),
    .io_bottom_out_valid(cols_8_15_io_bottom_out_valid),
    .io_bottom_out_bits(cols_8_15_io_bottom_out_bits)
  );
  ProcessingElement cols_9_15 ( // @[Stab.scala 85:60]
    .clock(cols_9_15_clock),
    .reset(cols_9_15_reset),
    .io_left_in_ready(cols_9_15_io_left_in_ready),
    .io_left_in_valid(cols_9_15_io_left_in_valid),
    .io_left_in_bits(cols_9_15_io_left_in_bits),
    .io_top_in_ready(cols_9_15_io_top_in_ready),
    .io_top_in_valid(cols_9_15_io_top_in_valid),
    .io_top_in_bits(cols_9_15_io_top_in_bits),
    .io_sum_ready(cols_9_15_io_sum_ready),
    .io_sum_valid(cols_9_15_io_sum_valid),
    .io_sum_bits(cols_9_15_io_sum_bits),
    .io_right_out_ready(cols_9_15_io_right_out_ready),
    .io_right_out_valid(cols_9_15_io_right_out_valid),
    .io_right_out_bits(cols_9_15_io_right_out_bits),
    .io_bottom_out_ready(cols_9_15_io_bottom_out_ready),
    .io_bottom_out_valid(cols_9_15_io_bottom_out_valid),
    .io_bottom_out_bits(cols_9_15_io_bottom_out_bits)
  );
  ProcessingElement cols_10_15 ( // @[Stab.scala 85:60]
    .clock(cols_10_15_clock),
    .reset(cols_10_15_reset),
    .io_left_in_ready(cols_10_15_io_left_in_ready),
    .io_left_in_valid(cols_10_15_io_left_in_valid),
    .io_left_in_bits(cols_10_15_io_left_in_bits),
    .io_top_in_ready(cols_10_15_io_top_in_ready),
    .io_top_in_valid(cols_10_15_io_top_in_valid),
    .io_top_in_bits(cols_10_15_io_top_in_bits),
    .io_sum_ready(cols_10_15_io_sum_ready),
    .io_sum_valid(cols_10_15_io_sum_valid),
    .io_sum_bits(cols_10_15_io_sum_bits),
    .io_right_out_ready(cols_10_15_io_right_out_ready),
    .io_right_out_valid(cols_10_15_io_right_out_valid),
    .io_right_out_bits(cols_10_15_io_right_out_bits),
    .io_bottom_out_ready(cols_10_15_io_bottom_out_ready),
    .io_bottom_out_valid(cols_10_15_io_bottom_out_valid),
    .io_bottom_out_bits(cols_10_15_io_bottom_out_bits)
  );
  ProcessingElement cols_11_15 ( // @[Stab.scala 85:60]
    .clock(cols_11_15_clock),
    .reset(cols_11_15_reset),
    .io_left_in_ready(cols_11_15_io_left_in_ready),
    .io_left_in_valid(cols_11_15_io_left_in_valid),
    .io_left_in_bits(cols_11_15_io_left_in_bits),
    .io_top_in_ready(cols_11_15_io_top_in_ready),
    .io_top_in_valid(cols_11_15_io_top_in_valid),
    .io_top_in_bits(cols_11_15_io_top_in_bits),
    .io_sum_ready(cols_11_15_io_sum_ready),
    .io_sum_valid(cols_11_15_io_sum_valid),
    .io_sum_bits(cols_11_15_io_sum_bits),
    .io_right_out_ready(cols_11_15_io_right_out_ready),
    .io_right_out_valid(cols_11_15_io_right_out_valid),
    .io_right_out_bits(cols_11_15_io_right_out_bits),
    .io_bottom_out_ready(cols_11_15_io_bottom_out_ready),
    .io_bottom_out_valid(cols_11_15_io_bottom_out_valid),
    .io_bottom_out_bits(cols_11_15_io_bottom_out_bits)
  );
  ProcessingElement cols_12_15 ( // @[Stab.scala 85:60]
    .clock(cols_12_15_clock),
    .reset(cols_12_15_reset),
    .io_left_in_ready(cols_12_15_io_left_in_ready),
    .io_left_in_valid(cols_12_15_io_left_in_valid),
    .io_left_in_bits(cols_12_15_io_left_in_bits),
    .io_top_in_ready(cols_12_15_io_top_in_ready),
    .io_top_in_valid(cols_12_15_io_top_in_valid),
    .io_top_in_bits(cols_12_15_io_top_in_bits),
    .io_sum_ready(cols_12_15_io_sum_ready),
    .io_sum_valid(cols_12_15_io_sum_valid),
    .io_sum_bits(cols_12_15_io_sum_bits),
    .io_right_out_ready(cols_12_15_io_right_out_ready),
    .io_right_out_valid(cols_12_15_io_right_out_valid),
    .io_right_out_bits(cols_12_15_io_right_out_bits),
    .io_bottom_out_ready(cols_12_15_io_bottom_out_ready),
    .io_bottom_out_valid(cols_12_15_io_bottom_out_valid),
    .io_bottom_out_bits(cols_12_15_io_bottom_out_bits)
  );
  ProcessingElement cols_13_15 ( // @[Stab.scala 85:60]
    .clock(cols_13_15_clock),
    .reset(cols_13_15_reset),
    .io_left_in_ready(cols_13_15_io_left_in_ready),
    .io_left_in_valid(cols_13_15_io_left_in_valid),
    .io_left_in_bits(cols_13_15_io_left_in_bits),
    .io_top_in_ready(cols_13_15_io_top_in_ready),
    .io_top_in_valid(cols_13_15_io_top_in_valid),
    .io_top_in_bits(cols_13_15_io_top_in_bits),
    .io_sum_ready(cols_13_15_io_sum_ready),
    .io_sum_valid(cols_13_15_io_sum_valid),
    .io_sum_bits(cols_13_15_io_sum_bits),
    .io_right_out_ready(cols_13_15_io_right_out_ready),
    .io_right_out_valid(cols_13_15_io_right_out_valid),
    .io_right_out_bits(cols_13_15_io_right_out_bits),
    .io_bottom_out_ready(cols_13_15_io_bottom_out_ready),
    .io_bottom_out_valid(cols_13_15_io_bottom_out_valid),
    .io_bottom_out_bits(cols_13_15_io_bottom_out_bits)
  );
  ProcessingElement cols_14_15 ( // @[Stab.scala 85:60]
    .clock(cols_14_15_clock),
    .reset(cols_14_15_reset),
    .io_left_in_ready(cols_14_15_io_left_in_ready),
    .io_left_in_valid(cols_14_15_io_left_in_valid),
    .io_left_in_bits(cols_14_15_io_left_in_bits),
    .io_top_in_ready(cols_14_15_io_top_in_ready),
    .io_top_in_valid(cols_14_15_io_top_in_valid),
    .io_top_in_bits(cols_14_15_io_top_in_bits),
    .io_sum_ready(cols_14_15_io_sum_ready),
    .io_sum_valid(cols_14_15_io_sum_valid),
    .io_sum_bits(cols_14_15_io_sum_bits),
    .io_right_out_ready(cols_14_15_io_right_out_ready),
    .io_right_out_valid(cols_14_15_io_right_out_valid),
    .io_right_out_bits(cols_14_15_io_right_out_bits),
    .io_bottom_out_ready(cols_14_15_io_bottom_out_ready),
    .io_bottom_out_valid(cols_14_15_io_bottom_out_valid),
    .io_bottom_out_bits(cols_14_15_io_bottom_out_bits)
  );
  ProcessingElement cols_15_15 ( // @[Stab.scala 85:60]
    .clock(cols_15_15_clock),
    .reset(cols_15_15_reset),
    .io_left_in_ready(cols_15_15_io_left_in_ready),
    .io_left_in_valid(cols_15_15_io_left_in_valid),
    .io_left_in_bits(cols_15_15_io_left_in_bits),
    .io_top_in_ready(cols_15_15_io_top_in_ready),
    .io_top_in_valid(cols_15_15_io_top_in_valid),
    .io_top_in_bits(cols_15_15_io_top_in_bits),
    .io_sum_ready(cols_15_15_io_sum_ready),
    .io_sum_valid(cols_15_15_io_sum_valid),
    .io_sum_bits(cols_15_15_io_sum_bits),
    .io_right_out_ready(cols_15_15_io_right_out_ready),
    .io_right_out_valid(cols_15_15_io_right_out_valid),
    .io_right_out_bits(cols_15_15_io_right_out_bits),
    .io_bottom_out_ready(cols_15_15_io_bottom_out_ready),
    .io_bottom_out_valid(cols_15_15_io_bottom_out_valid),
    .io_bottom_out_bits(cols_15_15_io_bottom_out_bits)
  );
  Queue q ( // @[Decoupled.scala 361:21]
    .clock(q_clock),
    .reset(q_reset),
    .io_enq_ready(q_io_enq_ready),
    .io_enq_valid(q_io_enq_valid),
    .io_enq_bits(q_io_enq_bits),
    .io_deq_ready(q_io_deq_ready),
    .io_deq_valid(q_io_deq_valid),
    .io_deq_bits(q_io_deq_bits)
  );
  Queue q_1 ( // @[Decoupled.scala 361:21]
    .clock(q_1_clock),
    .reset(q_1_reset),
    .io_enq_ready(q_1_io_enq_ready),
    .io_enq_valid(q_1_io_enq_valid),
    .io_enq_bits(q_1_io_enq_bits),
    .io_deq_ready(q_1_io_deq_ready),
    .io_deq_valid(q_1_io_deq_valid),
    .io_deq_bits(q_1_io_deq_bits)
  );
  Queue q_2 ( // @[Decoupled.scala 361:21]
    .clock(q_2_clock),
    .reset(q_2_reset),
    .io_enq_ready(q_2_io_enq_ready),
    .io_enq_valid(q_2_io_enq_valid),
    .io_enq_bits(q_2_io_enq_bits),
    .io_deq_ready(q_2_io_deq_ready),
    .io_deq_valid(q_2_io_deq_valid),
    .io_deq_bits(q_2_io_deq_bits)
  );
  Queue q_3 ( // @[Decoupled.scala 361:21]
    .clock(q_3_clock),
    .reset(q_3_reset),
    .io_enq_ready(q_3_io_enq_ready),
    .io_enq_valid(q_3_io_enq_valid),
    .io_enq_bits(q_3_io_enq_bits),
    .io_deq_ready(q_3_io_deq_ready),
    .io_deq_valid(q_3_io_deq_valid),
    .io_deq_bits(q_3_io_deq_bits)
  );
  Queue q_4 ( // @[Decoupled.scala 361:21]
    .clock(q_4_clock),
    .reset(q_4_reset),
    .io_enq_ready(q_4_io_enq_ready),
    .io_enq_valid(q_4_io_enq_valid),
    .io_enq_bits(q_4_io_enq_bits),
    .io_deq_ready(q_4_io_deq_ready),
    .io_deq_valid(q_4_io_deq_valid),
    .io_deq_bits(q_4_io_deq_bits)
  );
  Queue q_5 ( // @[Decoupled.scala 361:21]
    .clock(q_5_clock),
    .reset(q_5_reset),
    .io_enq_ready(q_5_io_enq_ready),
    .io_enq_valid(q_5_io_enq_valid),
    .io_enq_bits(q_5_io_enq_bits),
    .io_deq_ready(q_5_io_deq_ready),
    .io_deq_valid(q_5_io_deq_valid),
    .io_deq_bits(q_5_io_deq_bits)
  );
  Queue q_6 ( // @[Decoupled.scala 361:21]
    .clock(q_6_clock),
    .reset(q_6_reset),
    .io_enq_ready(q_6_io_enq_ready),
    .io_enq_valid(q_6_io_enq_valid),
    .io_enq_bits(q_6_io_enq_bits),
    .io_deq_ready(q_6_io_deq_ready),
    .io_deq_valid(q_6_io_deq_valid),
    .io_deq_bits(q_6_io_deq_bits)
  );
  Queue q_7 ( // @[Decoupled.scala 361:21]
    .clock(q_7_clock),
    .reset(q_7_reset),
    .io_enq_ready(q_7_io_enq_ready),
    .io_enq_valid(q_7_io_enq_valid),
    .io_enq_bits(q_7_io_enq_bits),
    .io_deq_ready(q_7_io_deq_ready),
    .io_deq_valid(q_7_io_deq_valid),
    .io_deq_bits(q_7_io_deq_bits)
  );
  Queue q_8 ( // @[Decoupled.scala 361:21]
    .clock(q_8_clock),
    .reset(q_8_reset),
    .io_enq_ready(q_8_io_enq_ready),
    .io_enq_valid(q_8_io_enq_valid),
    .io_enq_bits(q_8_io_enq_bits),
    .io_deq_ready(q_8_io_deq_ready),
    .io_deq_valid(q_8_io_deq_valid),
    .io_deq_bits(q_8_io_deq_bits)
  );
  Queue q_9 ( // @[Decoupled.scala 361:21]
    .clock(q_9_clock),
    .reset(q_9_reset),
    .io_enq_ready(q_9_io_enq_ready),
    .io_enq_valid(q_9_io_enq_valid),
    .io_enq_bits(q_9_io_enq_bits),
    .io_deq_ready(q_9_io_deq_ready),
    .io_deq_valid(q_9_io_deq_valid),
    .io_deq_bits(q_9_io_deq_bits)
  );
  Queue q_10 ( // @[Decoupled.scala 361:21]
    .clock(q_10_clock),
    .reset(q_10_reset),
    .io_enq_ready(q_10_io_enq_ready),
    .io_enq_valid(q_10_io_enq_valid),
    .io_enq_bits(q_10_io_enq_bits),
    .io_deq_ready(q_10_io_deq_ready),
    .io_deq_valid(q_10_io_deq_valid),
    .io_deq_bits(q_10_io_deq_bits)
  );
  Queue q_11 ( // @[Decoupled.scala 361:21]
    .clock(q_11_clock),
    .reset(q_11_reset),
    .io_enq_ready(q_11_io_enq_ready),
    .io_enq_valid(q_11_io_enq_valid),
    .io_enq_bits(q_11_io_enq_bits),
    .io_deq_ready(q_11_io_deq_ready),
    .io_deq_valid(q_11_io_deq_valid),
    .io_deq_bits(q_11_io_deq_bits)
  );
  Queue q_12 ( // @[Decoupled.scala 361:21]
    .clock(q_12_clock),
    .reset(q_12_reset),
    .io_enq_ready(q_12_io_enq_ready),
    .io_enq_valid(q_12_io_enq_valid),
    .io_enq_bits(q_12_io_enq_bits),
    .io_deq_ready(q_12_io_deq_ready),
    .io_deq_valid(q_12_io_deq_valid),
    .io_deq_bits(q_12_io_deq_bits)
  );
  Queue q_13 ( // @[Decoupled.scala 361:21]
    .clock(q_13_clock),
    .reset(q_13_reset),
    .io_enq_ready(q_13_io_enq_ready),
    .io_enq_valid(q_13_io_enq_valid),
    .io_enq_bits(q_13_io_enq_bits),
    .io_deq_ready(q_13_io_deq_ready),
    .io_deq_valid(q_13_io_deq_valid),
    .io_deq_bits(q_13_io_deq_bits)
  );
  Queue q_14 ( // @[Decoupled.scala 361:21]
    .clock(q_14_clock),
    .reset(q_14_reset),
    .io_enq_ready(q_14_io_enq_ready),
    .io_enq_valid(q_14_io_enq_valid),
    .io_enq_bits(q_14_io_enq_bits),
    .io_deq_ready(q_14_io_deq_ready),
    .io_deq_valid(q_14_io_deq_valid),
    .io_deq_bits(q_14_io_deq_bits)
  );
  Queue q_15 ( // @[Decoupled.scala 361:21]
    .clock(q_15_clock),
    .reset(q_15_reset),
    .io_enq_ready(q_15_io_enq_ready),
    .io_enq_valid(q_15_io_enq_valid),
    .io_enq_bits(q_15_io_enq_bits),
    .io_deq_ready(q_15_io_deq_ready),
    .io_deq_valid(q_15_io_deq_valid),
    .io_deq_bits(q_15_io_deq_bits)
  );
  Queue q_16 ( // @[Decoupled.scala 361:21]
    .clock(q_16_clock),
    .reset(q_16_reset),
    .io_enq_ready(q_16_io_enq_ready),
    .io_enq_valid(q_16_io_enq_valid),
    .io_enq_bits(q_16_io_enq_bits),
    .io_deq_ready(q_16_io_deq_ready),
    .io_deq_valid(q_16_io_deq_valid),
    .io_deq_bits(q_16_io_deq_bits)
  );
  Queue q_17 ( // @[Decoupled.scala 361:21]
    .clock(q_17_clock),
    .reset(q_17_reset),
    .io_enq_ready(q_17_io_enq_ready),
    .io_enq_valid(q_17_io_enq_valid),
    .io_enq_bits(q_17_io_enq_bits),
    .io_deq_ready(q_17_io_deq_ready),
    .io_deq_valid(q_17_io_deq_valid),
    .io_deq_bits(q_17_io_deq_bits)
  );
  Queue q_18 ( // @[Decoupled.scala 361:21]
    .clock(q_18_clock),
    .reset(q_18_reset),
    .io_enq_ready(q_18_io_enq_ready),
    .io_enq_valid(q_18_io_enq_valid),
    .io_enq_bits(q_18_io_enq_bits),
    .io_deq_ready(q_18_io_deq_ready),
    .io_deq_valid(q_18_io_deq_valid),
    .io_deq_bits(q_18_io_deq_bits)
  );
  Queue q_19 ( // @[Decoupled.scala 361:21]
    .clock(q_19_clock),
    .reset(q_19_reset),
    .io_enq_ready(q_19_io_enq_ready),
    .io_enq_valid(q_19_io_enq_valid),
    .io_enq_bits(q_19_io_enq_bits),
    .io_deq_ready(q_19_io_deq_ready),
    .io_deq_valid(q_19_io_deq_valid),
    .io_deq_bits(q_19_io_deq_bits)
  );
  Queue q_20 ( // @[Decoupled.scala 361:21]
    .clock(q_20_clock),
    .reset(q_20_reset),
    .io_enq_ready(q_20_io_enq_ready),
    .io_enq_valid(q_20_io_enq_valid),
    .io_enq_bits(q_20_io_enq_bits),
    .io_deq_ready(q_20_io_deq_ready),
    .io_deq_valid(q_20_io_deq_valid),
    .io_deq_bits(q_20_io_deq_bits)
  );
  Queue q_21 ( // @[Decoupled.scala 361:21]
    .clock(q_21_clock),
    .reset(q_21_reset),
    .io_enq_ready(q_21_io_enq_ready),
    .io_enq_valid(q_21_io_enq_valid),
    .io_enq_bits(q_21_io_enq_bits),
    .io_deq_ready(q_21_io_deq_ready),
    .io_deq_valid(q_21_io_deq_valid),
    .io_deq_bits(q_21_io_deq_bits)
  );
  Queue q_22 ( // @[Decoupled.scala 361:21]
    .clock(q_22_clock),
    .reset(q_22_reset),
    .io_enq_ready(q_22_io_enq_ready),
    .io_enq_valid(q_22_io_enq_valid),
    .io_enq_bits(q_22_io_enq_bits),
    .io_deq_ready(q_22_io_deq_ready),
    .io_deq_valid(q_22_io_deq_valid),
    .io_deq_bits(q_22_io_deq_bits)
  );
  Queue q_23 ( // @[Decoupled.scala 361:21]
    .clock(q_23_clock),
    .reset(q_23_reset),
    .io_enq_ready(q_23_io_enq_ready),
    .io_enq_valid(q_23_io_enq_valid),
    .io_enq_bits(q_23_io_enq_bits),
    .io_deq_ready(q_23_io_deq_ready),
    .io_deq_valid(q_23_io_deq_valid),
    .io_deq_bits(q_23_io_deq_bits)
  );
  Queue q_24 ( // @[Decoupled.scala 361:21]
    .clock(q_24_clock),
    .reset(q_24_reset),
    .io_enq_ready(q_24_io_enq_ready),
    .io_enq_valid(q_24_io_enq_valid),
    .io_enq_bits(q_24_io_enq_bits),
    .io_deq_ready(q_24_io_deq_ready),
    .io_deq_valid(q_24_io_deq_valid),
    .io_deq_bits(q_24_io_deq_bits)
  );
  Queue q_25 ( // @[Decoupled.scala 361:21]
    .clock(q_25_clock),
    .reset(q_25_reset),
    .io_enq_ready(q_25_io_enq_ready),
    .io_enq_valid(q_25_io_enq_valid),
    .io_enq_bits(q_25_io_enq_bits),
    .io_deq_ready(q_25_io_deq_ready),
    .io_deq_valid(q_25_io_deq_valid),
    .io_deq_bits(q_25_io_deq_bits)
  );
  Queue q_26 ( // @[Decoupled.scala 361:21]
    .clock(q_26_clock),
    .reset(q_26_reset),
    .io_enq_ready(q_26_io_enq_ready),
    .io_enq_valid(q_26_io_enq_valid),
    .io_enq_bits(q_26_io_enq_bits),
    .io_deq_ready(q_26_io_deq_ready),
    .io_deq_valid(q_26_io_deq_valid),
    .io_deq_bits(q_26_io_deq_bits)
  );
  Queue q_27 ( // @[Decoupled.scala 361:21]
    .clock(q_27_clock),
    .reset(q_27_reset),
    .io_enq_ready(q_27_io_enq_ready),
    .io_enq_valid(q_27_io_enq_valid),
    .io_enq_bits(q_27_io_enq_bits),
    .io_deq_ready(q_27_io_deq_ready),
    .io_deq_valid(q_27_io_deq_valid),
    .io_deq_bits(q_27_io_deq_bits)
  );
  Queue q_28 ( // @[Decoupled.scala 361:21]
    .clock(q_28_clock),
    .reset(q_28_reset),
    .io_enq_ready(q_28_io_enq_ready),
    .io_enq_valid(q_28_io_enq_valid),
    .io_enq_bits(q_28_io_enq_bits),
    .io_deq_ready(q_28_io_deq_ready),
    .io_deq_valid(q_28_io_deq_valid),
    .io_deq_bits(q_28_io_deq_bits)
  );
  Queue q_29 ( // @[Decoupled.scala 361:21]
    .clock(q_29_clock),
    .reset(q_29_reset),
    .io_enq_ready(q_29_io_enq_ready),
    .io_enq_valid(q_29_io_enq_valid),
    .io_enq_bits(q_29_io_enq_bits),
    .io_deq_ready(q_29_io_deq_ready),
    .io_deq_valid(q_29_io_deq_valid),
    .io_deq_bits(q_29_io_deq_bits)
  );
  Queue q_30 ( // @[Decoupled.scala 361:21]
    .clock(q_30_clock),
    .reset(q_30_reset),
    .io_enq_ready(q_30_io_enq_ready),
    .io_enq_valid(q_30_io_enq_valid),
    .io_enq_bits(q_30_io_enq_bits),
    .io_deq_ready(q_30_io_deq_ready),
    .io_deq_valid(q_30_io_deq_valid),
    .io_deq_bits(q_30_io_deq_bits)
  );
  Queue q_31 ( // @[Decoupled.scala 361:21]
    .clock(q_31_clock),
    .reset(q_31_reset),
    .io_enq_ready(q_31_io_enq_ready),
    .io_enq_valid(q_31_io_enq_valid),
    .io_enq_bits(q_31_io_enq_bits),
    .io_deq_ready(q_31_io_deq_ready),
    .io_deq_valid(q_31_io_deq_valid),
    .io_deq_bits(q_31_io_deq_bits)
  );
  Queue q_32 ( // @[Decoupled.scala 361:21]
    .clock(q_32_clock),
    .reset(q_32_reset),
    .io_enq_ready(q_32_io_enq_ready),
    .io_enq_valid(q_32_io_enq_valid),
    .io_enq_bits(q_32_io_enq_bits),
    .io_deq_ready(q_32_io_deq_ready),
    .io_deq_valid(q_32_io_deq_valid),
    .io_deq_bits(q_32_io_deq_bits)
  );
  Queue q_33 ( // @[Decoupled.scala 361:21]
    .clock(q_33_clock),
    .reset(q_33_reset),
    .io_enq_ready(q_33_io_enq_ready),
    .io_enq_valid(q_33_io_enq_valid),
    .io_enq_bits(q_33_io_enq_bits),
    .io_deq_ready(q_33_io_deq_ready),
    .io_deq_valid(q_33_io_deq_valid),
    .io_deq_bits(q_33_io_deq_bits)
  );
  Queue q_34 ( // @[Decoupled.scala 361:21]
    .clock(q_34_clock),
    .reset(q_34_reset),
    .io_enq_ready(q_34_io_enq_ready),
    .io_enq_valid(q_34_io_enq_valid),
    .io_enq_bits(q_34_io_enq_bits),
    .io_deq_ready(q_34_io_deq_ready),
    .io_deq_valid(q_34_io_deq_valid),
    .io_deq_bits(q_34_io_deq_bits)
  );
  Queue q_35 ( // @[Decoupled.scala 361:21]
    .clock(q_35_clock),
    .reset(q_35_reset),
    .io_enq_ready(q_35_io_enq_ready),
    .io_enq_valid(q_35_io_enq_valid),
    .io_enq_bits(q_35_io_enq_bits),
    .io_deq_ready(q_35_io_deq_ready),
    .io_deq_valid(q_35_io_deq_valid),
    .io_deq_bits(q_35_io_deq_bits)
  );
  Queue q_36 ( // @[Decoupled.scala 361:21]
    .clock(q_36_clock),
    .reset(q_36_reset),
    .io_enq_ready(q_36_io_enq_ready),
    .io_enq_valid(q_36_io_enq_valid),
    .io_enq_bits(q_36_io_enq_bits),
    .io_deq_ready(q_36_io_deq_ready),
    .io_deq_valid(q_36_io_deq_valid),
    .io_deq_bits(q_36_io_deq_bits)
  );
  Queue q_37 ( // @[Decoupled.scala 361:21]
    .clock(q_37_clock),
    .reset(q_37_reset),
    .io_enq_ready(q_37_io_enq_ready),
    .io_enq_valid(q_37_io_enq_valid),
    .io_enq_bits(q_37_io_enq_bits),
    .io_deq_ready(q_37_io_deq_ready),
    .io_deq_valid(q_37_io_deq_valid),
    .io_deq_bits(q_37_io_deq_bits)
  );
  Queue q_38 ( // @[Decoupled.scala 361:21]
    .clock(q_38_clock),
    .reset(q_38_reset),
    .io_enq_ready(q_38_io_enq_ready),
    .io_enq_valid(q_38_io_enq_valid),
    .io_enq_bits(q_38_io_enq_bits),
    .io_deq_ready(q_38_io_deq_ready),
    .io_deq_valid(q_38_io_deq_valid),
    .io_deq_bits(q_38_io_deq_bits)
  );
  Queue q_39 ( // @[Decoupled.scala 361:21]
    .clock(q_39_clock),
    .reset(q_39_reset),
    .io_enq_ready(q_39_io_enq_ready),
    .io_enq_valid(q_39_io_enq_valid),
    .io_enq_bits(q_39_io_enq_bits),
    .io_deq_ready(q_39_io_deq_ready),
    .io_deq_valid(q_39_io_deq_valid),
    .io_deq_bits(q_39_io_deq_bits)
  );
  Queue q_40 ( // @[Decoupled.scala 361:21]
    .clock(q_40_clock),
    .reset(q_40_reset),
    .io_enq_ready(q_40_io_enq_ready),
    .io_enq_valid(q_40_io_enq_valid),
    .io_enq_bits(q_40_io_enq_bits),
    .io_deq_ready(q_40_io_deq_ready),
    .io_deq_valid(q_40_io_deq_valid),
    .io_deq_bits(q_40_io_deq_bits)
  );
  Queue q_41 ( // @[Decoupled.scala 361:21]
    .clock(q_41_clock),
    .reset(q_41_reset),
    .io_enq_ready(q_41_io_enq_ready),
    .io_enq_valid(q_41_io_enq_valid),
    .io_enq_bits(q_41_io_enq_bits),
    .io_deq_ready(q_41_io_deq_ready),
    .io_deq_valid(q_41_io_deq_valid),
    .io_deq_bits(q_41_io_deq_bits)
  );
  Queue q_42 ( // @[Decoupled.scala 361:21]
    .clock(q_42_clock),
    .reset(q_42_reset),
    .io_enq_ready(q_42_io_enq_ready),
    .io_enq_valid(q_42_io_enq_valid),
    .io_enq_bits(q_42_io_enq_bits),
    .io_deq_ready(q_42_io_deq_ready),
    .io_deq_valid(q_42_io_deq_valid),
    .io_deq_bits(q_42_io_deq_bits)
  );
  Queue q_43 ( // @[Decoupled.scala 361:21]
    .clock(q_43_clock),
    .reset(q_43_reset),
    .io_enq_ready(q_43_io_enq_ready),
    .io_enq_valid(q_43_io_enq_valid),
    .io_enq_bits(q_43_io_enq_bits),
    .io_deq_ready(q_43_io_deq_ready),
    .io_deq_valid(q_43_io_deq_valid),
    .io_deq_bits(q_43_io_deq_bits)
  );
  Queue q_44 ( // @[Decoupled.scala 361:21]
    .clock(q_44_clock),
    .reset(q_44_reset),
    .io_enq_ready(q_44_io_enq_ready),
    .io_enq_valid(q_44_io_enq_valid),
    .io_enq_bits(q_44_io_enq_bits),
    .io_deq_ready(q_44_io_deq_ready),
    .io_deq_valid(q_44_io_deq_valid),
    .io_deq_bits(q_44_io_deq_bits)
  );
  Queue q_45 ( // @[Decoupled.scala 361:21]
    .clock(q_45_clock),
    .reset(q_45_reset),
    .io_enq_ready(q_45_io_enq_ready),
    .io_enq_valid(q_45_io_enq_valid),
    .io_enq_bits(q_45_io_enq_bits),
    .io_deq_ready(q_45_io_deq_ready),
    .io_deq_valid(q_45_io_deq_valid),
    .io_deq_bits(q_45_io_deq_bits)
  );
  Queue q_46 ( // @[Decoupled.scala 361:21]
    .clock(q_46_clock),
    .reset(q_46_reset),
    .io_enq_ready(q_46_io_enq_ready),
    .io_enq_valid(q_46_io_enq_valid),
    .io_enq_bits(q_46_io_enq_bits),
    .io_deq_ready(q_46_io_deq_ready),
    .io_deq_valid(q_46_io_deq_valid),
    .io_deq_bits(q_46_io_deq_bits)
  );
  Queue q_47 ( // @[Decoupled.scala 361:21]
    .clock(q_47_clock),
    .reset(q_47_reset),
    .io_enq_ready(q_47_io_enq_ready),
    .io_enq_valid(q_47_io_enq_valid),
    .io_enq_bits(q_47_io_enq_bits),
    .io_deq_ready(q_47_io_deq_ready),
    .io_deq_valid(q_47_io_deq_valid),
    .io_deq_bits(q_47_io_deq_bits)
  );
  Queue q_48 ( // @[Decoupled.scala 361:21]
    .clock(q_48_clock),
    .reset(q_48_reset),
    .io_enq_ready(q_48_io_enq_ready),
    .io_enq_valid(q_48_io_enq_valid),
    .io_enq_bits(q_48_io_enq_bits),
    .io_deq_ready(q_48_io_deq_ready),
    .io_deq_valid(q_48_io_deq_valid),
    .io_deq_bits(q_48_io_deq_bits)
  );
  Queue q_49 ( // @[Decoupled.scala 361:21]
    .clock(q_49_clock),
    .reset(q_49_reset),
    .io_enq_ready(q_49_io_enq_ready),
    .io_enq_valid(q_49_io_enq_valid),
    .io_enq_bits(q_49_io_enq_bits),
    .io_deq_ready(q_49_io_deq_ready),
    .io_deq_valid(q_49_io_deq_valid),
    .io_deq_bits(q_49_io_deq_bits)
  );
  Queue q_50 ( // @[Decoupled.scala 361:21]
    .clock(q_50_clock),
    .reset(q_50_reset),
    .io_enq_ready(q_50_io_enq_ready),
    .io_enq_valid(q_50_io_enq_valid),
    .io_enq_bits(q_50_io_enq_bits),
    .io_deq_ready(q_50_io_deq_ready),
    .io_deq_valid(q_50_io_deq_valid),
    .io_deq_bits(q_50_io_deq_bits)
  );
  Queue q_51 ( // @[Decoupled.scala 361:21]
    .clock(q_51_clock),
    .reset(q_51_reset),
    .io_enq_ready(q_51_io_enq_ready),
    .io_enq_valid(q_51_io_enq_valid),
    .io_enq_bits(q_51_io_enq_bits),
    .io_deq_ready(q_51_io_deq_ready),
    .io_deq_valid(q_51_io_deq_valid),
    .io_deq_bits(q_51_io_deq_bits)
  );
  Queue q_52 ( // @[Decoupled.scala 361:21]
    .clock(q_52_clock),
    .reset(q_52_reset),
    .io_enq_ready(q_52_io_enq_ready),
    .io_enq_valid(q_52_io_enq_valid),
    .io_enq_bits(q_52_io_enq_bits),
    .io_deq_ready(q_52_io_deq_ready),
    .io_deq_valid(q_52_io_deq_valid),
    .io_deq_bits(q_52_io_deq_bits)
  );
  Queue q_53 ( // @[Decoupled.scala 361:21]
    .clock(q_53_clock),
    .reset(q_53_reset),
    .io_enq_ready(q_53_io_enq_ready),
    .io_enq_valid(q_53_io_enq_valid),
    .io_enq_bits(q_53_io_enq_bits),
    .io_deq_ready(q_53_io_deq_ready),
    .io_deq_valid(q_53_io_deq_valid),
    .io_deq_bits(q_53_io_deq_bits)
  );
  Queue q_54 ( // @[Decoupled.scala 361:21]
    .clock(q_54_clock),
    .reset(q_54_reset),
    .io_enq_ready(q_54_io_enq_ready),
    .io_enq_valid(q_54_io_enq_valid),
    .io_enq_bits(q_54_io_enq_bits),
    .io_deq_ready(q_54_io_deq_ready),
    .io_deq_valid(q_54_io_deq_valid),
    .io_deq_bits(q_54_io_deq_bits)
  );
  Queue q_55 ( // @[Decoupled.scala 361:21]
    .clock(q_55_clock),
    .reset(q_55_reset),
    .io_enq_ready(q_55_io_enq_ready),
    .io_enq_valid(q_55_io_enq_valid),
    .io_enq_bits(q_55_io_enq_bits),
    .io_deq_ready(q_55_io_deq_ready),
    .io_deq_valid(q_55_io_deq_valid),
    .io_deq_bits(q_55_io_deq_bits)
  );
  Queue q_56 ( // @[Decoupled.scala 361:21]
    .clock(q_56_clock),
    .reset(q_56_reset),
    .io_enq_ready(q_56_io_enq_ready),
    .io_enq_valid(q_56_io_enq_valid),
    .io_enq_bits(q_56_io_enq_bits),
    .io_deq_ready(q_56_io_deq_ready),
    .io_deq_valid(q_56_io_deq_valid),
    .io_deq_bits(q_56_io_deq_bits)
  );
  Queue q_57 ( // @[Decoupled.scala 361:21]
    .clock(q_57_clock),
    .reset(q_57_reset),
    .io_enq_ready(q_57_io_enq_ready),
    .io_enq_valid(q_57_io_enq_valid),
    .io_enq_bits(q_57_io_enq_bits),
    .io_deq_ready(q_57_io_deq_ready),
    .io_deq_valid(q_57_io_deq_valid),
    .io_deq_bits(q_57_io_deq_bits)
  );
  Queue q_58 ( // @[Decoupled.scala 361:21]
    .clock(q_58_clock),
    .reset(q_58_reset),
    .io_enq_ready(q_58_io_enq_ready),
    .io_enq_valid(q_58_io_enq_valid),
    .io_enq_bits(q_58_io_enq_bits),
    .io_deq_ready(q_58_io_deq_ready),
    .io_deq_valid(q_58_io_deq_valid),
    .io_deq_bits(q_58_io_deq_bits)
  );
  Queue q_59 ( // @[Decoupled.scala 361:21]
    .clock(q_59_clock),
    .reset(q_59_reset),
    .io_enq_ready(q_59_io_enq_ready),
    .io_enq_valid(q_59_io_enq_valid),
    .io_enq_bits(q_59_io_enq_bits),
    .io_deq_ready(q_59_io_deq_ready),
    .io_deq_valid(q_59_io_deq_valid),
    .io_deq_bits(q_59_io_deq_bits)
  );
  Queue q_60 ( // @[Decoupled.scala 361:21]
    .clock(q_60_clock),
    .reset(q_60_reset),
    .io_enq_ready(q_60_io_enq_ready),
    .io_enq_valid(q_60_io_enq_valid),
    .io_enq_bits(q_60_io_enq_bits),
    .io_deq_ready(q_60_io_deq_ready),
    .io_deq_valid(q_60_io_deq_valid),
    .io_deq_bits(q_60_io_deq_bits)
  );
  Queue q_61 ( // @[Decoupled.scala 361:21]
    .clock(q_61_clock),
    .reset(q_61_reset),
    .io_enq_ready(q_61_io_enq_ready),
    .io_enq_valid(q_61_io_enq_valid),
    .io_enq_bits(q_61_io_enq_bits),
    .io_deq_ready(q_61_io_deq_ready),
    .io_deq_valid(q_61_io_deq_valid),
    .io_deq_bits(q_61_io_deq_bits)
  );
  Queue q_62 ( // @[Decoupled.scala 361:21]
    .clock(q_62_clock),
    .reset(q_62_reset),
    .io_enq_ready(q_62_io_enq_ready),
    .io_enq_valid(q_62_io_enq_valid),
    .io_enq_bits(q_62_io_enq_bits),
    .io_deq_ready(q_62_io_deq_ready),
    .io_deq_valid(q_62_io_deq_valid),
    .io_deq_bits(q_62_io_deq_bits)
  );
  Queue q_63 ( // @[Decoupled.scala 361:21]
    .clock(q_63_clock),
    .reset(q_63_reset),
    .io_enq_ready(q_63_io_enq_ready),
    .io_enq_valid(q_63_io_enq_valid),
    .io_enq_bits(q_63_io_enq_bits),
    .io_deq_ready(q_63_io_deq_ready),
    .io_deq_valid(q_63_io_deq_valid),
    .io_deq_bits(q_63_io_deq_bits)
  );
  Queue q_64 ( // @[Decoupled.scala 361:21]
    .clock(q_64_clock),
    .reset(q_64_reset),
    .io_enq_ready(q_64_io_enq_ready),
    .io_enq_valid(q_64_io_enq_valid),
    .io_enq_bits(q_64_io_enq_bits),
    .io_deq_ready(q_64_io_deq_ready),
    .io_deq_valid(q_64_io_deq_valid),
    .io_deq_bits(q_64_io_deq_bits)
  );
  Queue q_65 ( // @[Decoupled.scala 361:21]
    .clock(q_65_clock),
    .reset(q_65_reset),
    .io_enq_ready(q_65_io_enq_ready),
    .io_enq_valid(q_65_io_enq_valid),
    .io_enq_bits(q_65_io_enq_bits),
    .io_deq_ready(q_65_io_deq_ready),
    .io_deq_valid(q_65_io_deq_valid),
    .io_deq_bits(q_65_io_deq_bits)
  );
  Queue q_66 ( // @[Decoupled.scala 361:21]
    .clock(q_66_clock),
    .reset(q_66_reset),
    .io_enq_ready(q_66_io_enq_ready),
    .io_enq_valid(q_66_io_enq_valid),
    .io_enq_bits(q_66_io_enq_bits),
    .io_deq_ready(q_66_io_deq_ready),
    .io_deq_valid(q_66_io_deq_valid),
    .io_deq_bits(q_66_io_deq_bits)
  );
  Queue q_67 ( // @[Decoupled.scala 361:21]
    .clock(q_67_clock),
    .reset(q_67_reset),
    .io_enq_ready(q_67_io_enq_ready),
    .io_enq_valid(q_67_io_enq_valid),
    .io_enq_bits(q_67_io_enq_bits),
    .io_deq_ready(q_67_io_deq_ready),
    .io_deq_valid(q_67_io_deq_valid),
    .io_deq_bits(q_67_io_deq_bits)
  );
  Queue q_68 ( // @[Decoupled.scala 361:21]
    .clock(q_68_clock),
    .reset(q_68_reset),
    .io_enq_ready(q_68_io_enq_ready),
    .io_enq_valid(q_68_io_enq_valid),
    .io_enq_bits(q_68_io_enq_bits),
    .io_deq_ready(q_68_io_deq_ready),
    .io_deq_valid(q_68_io_deq_valid),
    .io_deq_bits(q_68_io_deq_bits)
  );
  Queue q_69 ( // @[Decoupled.scala 361:21]
    .clock(q_69_clock),
    .reset(q_69_reset),
    .io_enq_ready(q_69_io_enq_ready),
    .io_enq_valid(q_69_io_enq_valid),
    .io_enq_bits(q_69_io_enq_bits),
    .io_deq_ready(q_69_io_deq_ready),
    .io_deq_valid(q_69_io_deq_valid),
    .io_deq_bits(q_69_io_deq_bits)
  );
  Queue q_70 ( // @[Decoupled.scala 361:21]
    .clock(q_70_clock),
    .reset(q_70_reset),
    .io_enq_ready(q_70_io_enq_ready),
    .io_enq_valid(q_70_io_enq_valid),
    .io_enq_bits(q_70_io_enq_bits),
    .io_deq_ready(q_70_io_deq_ready),
    .io_deq_valid(q_70_io_deq_valid),
    .io_deq_bits(q_70_io_deq_bits)
  );
  Queue q_71 ( // @[Decoupled.scala 361:21]
    .clock(q_71_clock),
    .reset(q_71_reset),
    .io_enq_ready(q_71_io_enq_ready),
    .io_enq_valid(q_71_io_enq_valid),
    .io_enq_bits(q_71_io_enq_bits),
    .io_deq_ready(q_71_io_deq_ready),
    .io_deq_valid(q_71_io_deq_valid),
    .io_deq_bits(q_71_io_deq_bits)
  );
  Queue q_72 ( // @[Decoupled.scala 361:21]
    .clock(q_72_clock),
    .reset(q_72_reset),
    .io_enq_ready(q_72_io_enq_ready),
    .io_enq_valid(q_72_io_enq_valid),
    .io_enq_bits(q_72_io_enq_bits),
    .io_deq_ready(q_72_io_deq_ready),
    .io_deq_valid(q_72_io_deq_valid),
    .io_deq_bits(q_72_io_deq_bits)
  );
  Queue q_73 ( // @[Decoupled.scala 361:21]
    .clock(q_73_clock),
    .reset(q_73_reset),
    .io_enq_ready(q_73_io_enq_ready),
    .io_enq_valid(q_73_io_enq_valid),
    .io_enq_bits(q_73_io_enq_bits),
    .io_deq_ready(q_73_io_deq_ready),
    .io_deq_valid(q_73_io_deq_valid),
    .io_deq_bits(q_73_io_deq_bits)
  );
  Queue q_74 ( // @[Decoupled.scala 361:21]
    .clock(q_74_clock),
    .reset(q_74_reset),
    .io_enq_ready(q_74_io_enq_ready),
    .io_enq_valid(q_74_io_enq_valid),
    .io_enq_bits(q_74_io_enq_bits),
    .io_deq_ready(q_74_io_deq_ready),
    .io_deq_valid(q_74_io_deq_valid),
    .io_deq_bits(q_74_io_deq_bits)
  );
  Queue q_75 ( // @[Decoupled.scala 361:21]
    .clock(q_75_clock),
    .reset(q_75_reset),
    .io_enq_ready(q_75_io_enq_ready),
    .io_enq_valid(q_75_io_enq_valid),
    .io_enq_bits(q_75_io_enq_bits),
    .io_deq_ready(q_75_io_deq_ready),
    .io_deq_valid(q_75_io_deq_valid),
    .io_deq_bits(q_75_io_deq_bits)
  );
  Queue q_76 ( // @[Decoupled.scala 361:21]
    .clock(q_76_clock),
    .reset(q_76_reset),
    .io_enq_ready(q_76_io_enq_ready),
    .io_enq_valid(q_76_io_enq_valid),
    .io_enq_bits(q_76_io_enq_bits),
    .io_deq_ready(q_76_io_deq_ready),
    .io_deq_valid(q_76_io_deq_valid),
    .io_deq_bits(q_76_io_deq_bits)
  );
  Queue q_77 ( // @[Decoupled.scala 361:21]
    .clock(q_77_clock),
    .reset(q_77_reset),
    .io_enq_ready(q_77_io_enq_ready),
    .io_enq_valid(q_77_io_enq_valid),
    .io_enq_bits(q_77_io_enq_bits),
    .io_deq_ready(q_77_io_deq_ready),
    .io_deq_valid(q_77_io_deq_valid),
    .io_deq_bits(q_77_io_deq_bits)
  );
  Queue q_78 ( // @[Decoupled.scala 361:21]
    .clock(q_78_clock),
    .reset(q_78_reset),
    .io_enq_ready(q_78_io_enq_ready),
    .io_enq_valid(q_78_io_enq_valid),
    .io_enq_bits(q_78_io_enq_bits),
    .io_deq_ready(q_78_io_deq_ready),
    .io_deq_valid(q_78_io_deq_valid),
    .io_deq_bits(q_78_io_deq_bits)
  );
  Queue q_79 ( // @[Decoupled.scala 361:21]
    .clock(q_79_clock),
    .reset(q_79_reset),
    .io_enq_ready(q_79_io_enq_ready),
    .io_enq_valid(q_79_io_enq_valid),
    .io_enq_bits(q_79_io_enq_bits),
    .io_deq_ready(q_79_io_deq_ready),
    .io_deq_valid(q_79_io_deq_valid),
    .io_deq_bits(q_79_io_deq_bits)
  );
  Queue q_80 ( // @[Decoupled.scala 361:21]
    .clock(q_80_clock),
    .reset(q_80_reset),
    .io_enq_ready(q_80_io_enq_ready),
    .io_enq_valid(q_80_io_enq_valid),
    .io_enq_bits(q_80_io_enq_bits),
    .io_deq_ready(q_80_io_deq_ready),
    .io_deq_valid(q_80_io_deq_valid),
    .io_deq_bits(q_80_io_deq_bits)
  );
  Queue q_81 ( // @[Decoupled.scala 361:21]
    .clock(q_81_clock),
    .reset(q_81_reset),
    .io_enq_ready(q_81_io_enq_ready),
    .io_enq_valid(q_81_io_enq_valid),
    .io_enq_bits(q_81_io_enq_bits),
    .io_deq_ready(q_81_io_deq_ready),
    .io_deq_valid(q_81_io_deq_valid),
    .io_deq_bits(q_81_io_deq_bits)
  );
  Queue q_82 ( // @[Decoupled.scala 361:21]
    .clock(q_82_clock),
    .reset(q_82_reset),
    .io_enq_ready(q_82_io_enq_ready),
    .io_enq_valid(q_82_io_enq_valid),
    .io_enq_bits(q_82_io_enq_bits),
    .io_deq_ready(q_82_io_deq_ready),
    .io_deq_valid(q_82_io_deq_valid),
    .io_deq_bits(q_82_io_deq_bits)
  );
  Queue q_83 ( // @[Decoupled.scala 361:21]
    .clock(q_83_clock),
    .reset(q_83_reset),
    .io_enq_ready(q_83_io_enq_ready),
    .io_enq_valid(q_83_io_enq_valid),
    .io_enq_bits(q_83_io_enq_bits),
    .io_deq_ready(q_83_io_deq_ready),
    .io_deq_valid(q_83_io_deq_valid),
    .io_deq_bits(q_83_io_deq_bits)
  );
  Queue q_84 ( // @[Decoupled.scala 361:21]
    .clock(q_84_clock),
    .reset(q_84_reset),
    .io_enq_ready(q_84_io_enq_ready),
    .io_enq_valid(q_84_io_enq_valid),
    .io_enq_bits(q_84_io_enq_bits),
    .io_deq_ready(q_84_io_deq_ready),
    .io_deq_valid(q_84_io_deq_valid),
    .io_deq_bits(q_84_io_deq_bits)
  );
  Queue q_85 ( // @[Decoupled.scala 361:21]
    .clock(q_85_clock),
    .reset(q_85_reset),
    .io_enq_ready(q_85_io_enq_ready),
    .io_enq_valid(q_85_io_enq_valid),
    .io_enq_bits(q_85_io_enq_bits),
    .io_deq_ready(q_85_io_deq_ready),
    .io_deq_valid(q_85_io_deq_valid),
    .io_deq_bits(q_85_io_deq_bits)
  );
  Queue q_86 ( // @[Decoupled.scala 361:21]
    .clock(q_86_clock),
    .reset(q_86_reset),
    .io_enq_ready(q_86_io_enq_ready),
    .io_enq_valid(q_86_io_enq_valid),
    .io_enq_bits(q_86_io_enq_bits),
    .io_deq_ready(q_86_io_deq_ready),
    .io_deq_valid(q_86_io_deq_valid),
    .io_deq_bits(q_86_io_deq_bits)
  );
  Queue q_87 ( // @[Decoupled.scala 361:21]
    .clock(q_87_clock),
    .reset(q_87_reset),
    .io_enq_ready(q_87_io_enq_ready),
    .io_enq_valid(q_87_io_enq_valid),
    .io_enq_bits(q_87_io_enq_bits),
    .io_deq_ready(q_87_io_deq_ready),
    .io_deq_valid(q_87_io_deq_valid),
    .io_deq_bits(q_87_io_deq_bits)
  );
  Queue q_88 ( // @[Decoupled.scala 361:21]
    .clock(q_88_clock),
    .reset(q_88_reset),
    .io_enq_ready(q_88_io_enq_ready),
    .io_enq_valid(q_88_io_enq_valid),
    .io_enq_bits(q_88_io_enq_bits),
    .io_deq_ready(q_88_io_deq_ready),
    .io_deq_valid(q_88_io_deq_valid),
    .io_deq_bits(q_88_io_deq_bits)
  );
  Queue q_89 ( // @[Decoupled.scala 361:21]
    .clock(q_89_clock),
    .reset(q_89_reset),
    .io_enq_ready(q_89_io_enq_ready),
    .io_enq_valid(q_89_io_enq_valid),
    .io_enq_bits(q_89_io_enq_bits),
    .io_deq_ready(q_89_io_deq_ready),
    .io_deq_valid(q_89_io_deq_valid),
    .io_deq_bits(q_89_io_deq_bits)
  );
  Queue q_90 ( // @[Decoupled.scala 361:21]
    .clock(q_90_clock),
    .reset(q_90_reset),
    .io_enq_ready(q_90_io_enq_ready),
    .io_enq_valid(q_90_io_enq_valid),
    .io_enq_bits(q_90_io_enq_bits),
    .io_deq_ready(q_90_io_deq_ready),
    .io_deq_valid(q_90_io_deq_valid),
    .io_deq_bits(q_90_io_deq_bits)
  );
  Queue q_91 ( // @[Decoupled.scala 361:21]
    .clock(q_91_clock),
    .reset(q_91_reset),
    .io_enq_ready(q_91_io_enq_ready),
    .io_enq_valid(q_91_io_enq_valid),
    .io_enq_bits(q_91_io_enq_bits),
    .io_deq_ready(q_91_io_deq_ready),
    .io_deq_valid(q_91_io_deq_valid),
    .io_deq_bits(q_91_io_deq_bits)
  );
  Queue q_92 ( // @[Decoupled.scala 361:21]
    .clock(q_92_clock),
    .reset(q_92_reset),
    .io_enq_ready(q_92_io_enq_ready),
    .io_enq_valid(q_92_io_enq_valid),
    .io_enq_bits(q_92_io_enq_bits),
    .io_deq_ready(q_92_io_deq_ready),
    .io_deq_valid(q_92_io_deq_valid),
    .io_deq_bits(q_92_io_deq_bits)
  );
  Queue q_93 ( // @[Decoupled.scala 361:21]
    .clock(q_93_clock),
    .reset(q_93_reset),
    .io_enq_ready(q_93_io_enq_ready),
    .io_enq_valid(q_93_io_enq_valid),
    .io_enq_bits(q_93_io_enq_bits),
    .io_deq_ready(q_93_io_deq_ready),
    .io_deq_valid(q_93_io_deq_valid),
    .io_deq_bits(q_93_io_deq_bits)
  );
  Queue q_94 ( // @[Decoupled.scala 361:21]
    .clock(q_94_clock),
    .reset(q_94_reset),
    .io_enq_ready(q_94_io_enq_ready),
    .io_enq_valid(q_94_io_enq_valid),
    .io_enq_bits(q_94_io_enq_bits),
    .io_deq_ready(q_94_io_deq_ready),
    .io_deq_valid(q_94_io_deq_valid),
    .io_deq_bits(q_94_io_deq_bits)
  );
  Queue q_95 ( // @[Decoupled.scala 361:21]
    .clock(q_95_clock),
    .reset(q_95_reset),
    .io_enq_ready(q_95_io_enq_ready),
    .io_enq_valid(q_95_io_enq_valid),
    .io_enq_bits(q_95_io_enq_bits),
    .io_deq_ready(q_95_io_deq_ready),
    .io_deq_valid(q_95_io_deq_valid),
    .io_deq_bits(q_95_io_deq_bits)
  );
  Queue q_96 ( // @[Decoupled.scala 361:21]
    .clock(q_96_clock),
    .reset(q_96_reset),
    .io_enq_ready(q_96_io_enq_ready),
    .io_enq_valid(q_96_io_enq_valid),
    .io_enq_bits(q_96_io_enq_bits),
    .io_deq_ready(q_96_io_deq_ready),
    .io_deq_valid(q_96_io_deq_valid),
    .io_deq_bits(q_96_io_deq_bits)
  );
  Queue q_97 ( // @[Decoupled.scala 361:21]
    .clock(q_97_clock),
    .reset(q_97_reset),
    .io_enq_ready(q_97_io_enq_ready),
    .io_enq_valid(q_97_io_enq_valid),
    .io_enq_bits(q_97_io_enq_bits),
    .io_deq_ready(q_97_io_deq_ready),
    .io_deq_valid(q_97_io_deq_valid),
    .io_deq_bits(q_97_io_deq_bits)
  );
  Queue q_98 ( // @[Decoupled.scala 361:21]
    .clock(q_98_clock),
    .reset(q_98_reset),
    .io_enq_ready(q_98_io_enq_ready),
    .io_enq_valid(q_98_io_enq_valid),
    .io_enq_bits(q_98_io_enq_bits),
    .io_deq_ready(q_98_io_deq_ready),
    .io_deq_valid(q_98_io_deq_valid),
    .io_deq_bits(q_98_io_deq_bits)
  );
  Queue q_99 ( // @[Decoupled.scala 361:21]
    .clock(q_99_clock),
    .reset(q_99_reset),
    .io_enq_ready(q_99_io_enq_ready),
    .io_enq_valid(q_99_io_enq_valid),
    .io_enq_bits(q_99_io_enq_bits),
    .io_deq_ready(q_99_io_deq_ready),
    .io_deq_valid(q_99_io_deq_valid),
    .io_deq_bits(q_99_io_deq_bits)
  );
  Queue q_100 ( // @[Decoupled.scala 361:21]
    .clock(q_100_clock),
    .reset(q_100_reset),
    .io_enq_ready(q_100_io_enq_ready),
    .io_enq_valid(q_100_io_enq_valid),
    .io_enq_bits(q_100_io_enq_bits),
    .io_deq_ready(q_100_io_deq_ready),
    .io_deq_valid(q_100_io_deq_valid),
    .io_deq_bits(q_100_io_deq_bits)
  );
  Queue q_101 ( // @[Decoupled.scala 361:21]
    .clock(q_101_clock),
    .reset(q_101_reset),
    .io_enq_ready(q_101_io_enq_ready),
    .io_enq_valid(q_101_io_enq_valid),
    .io_enq_bits(q_101_io_enq_bits),
    .io_deq_ready(q_101_io_deq_ready),
    .io_deq_valid(q_101_io_deq_valid),
    .io_deq_bits(q_101_io_deq_bits)
  );
  Queue q_102 ( // @[Decoupled.scala 361:21]
    .clock(q_102_clock),
    .reset(q_102_reset),
    .io_enq_ready(q_102_io_enq_ready),
    .io_enq_valid(q_102_io_enq_valid),
    .io_enq_bits(q_102_io_enq_bits),
    .io_deq_ready(q_102_io_deq_ready),
    .io_deq_valid(q_102_io_deq_valid),
    .io_deq_bits(q_102_io_deq_bits)
  );
  Queue q_103 ( // @[Decoupled.scala 361:21]
    .clock(q_103_clock),
    .reset(q_103_reset),
    .io_enq_ready(q_103_io_enq_ready),
    .io_enq_valid(q_103_io_enq_valid),
    .io_enq_bits(q_103_io_enq_bits),
    .io_deq_ready(q_103_io_deq_ready),
    .io_deq_valid(q_103_io_deq_valid),
    .io_deq_bits(q_103_io_deq_bits)
  );
  Queue q_104 ( // @[Decoupled.scala 361:21]
    .clock(q_104_clock),
    .reset(q_104_reset),
    .io_enq_ready(q_104_io_enq_ready),
    .io_enq_valid(q_104_io_enq_valid),
    .io_enq_bits(q_104_io_enq_bits),
    .io_deq_ready(q_104_io_deq_ready),
    .io_deq_valid(q_104_io_deq_valid),
    .io_deq_bits(q_104_io_deq_bits)
  );
  Queue q_105 ( // @[Decoupled.scala 361:21]
    .clock(q_105_clock),
    .reset(q_105_reset),
    .io_enq_ready(q_105_io_enq_ready),
    .io_enq_valid(q_105_io_enq_valid),
    .io_enq_bits(q_105_io_enq_bits),
    .io_deq_ready(q_105_io_deq_ready),
    .io_deq_valid(q_105_io_deq_valid),
    .io_deq_bits(q_105_io_deq_bits)
  );
  Queue q_106 ( // @[Decoupled.scala 361:21]
    .clock(q_106_clock),
    .reset(q_106_reset),
    .io_enq_ready(q_106_io_enq_ready),
    .io_enq_valid(q_106_io_enq_valid),
    .io_enq_bits(q_106_io_enq_bits),
    .io_deq_ready(q_106_io_deq_ready),
    .io_deq_valid(q_106_io_deq_valid),
    .io_deq_bits(q_106_io_deq_bits)
  );
  Queue q_107 ( // @[Decoupled.scala 361:21]
    .clock(q_107_clock),
    .reset(q_107_reset),
    .io_enq_ready(q_107_io_enq_ready),
    .io_enq_valid(q_107_io_enq_valid),
    .io_enq_bits(q_107_io_enq_bits),
    .io_deq_ready(q_107_io_deq_ready),
    .io_deq_valid(q_107_io_deq_valid),
    .io_deq_bits(q_107_io_deq_bits)
  );
  Queue q_108 ( // @[Decoupled.scala 361:21]
    .clock(q_108_clock),
    .reset(q_108_reset),
    .io_enq_ready(q_108_io_enq_ready),
    .io_enq_valid(q_108_io_enq_valid),
    .io_enq_bits(q_108_io_enq_bits),
    .io_deq_ready(q_108_io_deq_ready),
    .io_deq_valid(q_108_io_deq_valid),
    .io_deq_bits(q_108_io_deq_bits)
  );
  Queue q_109 ( // @[Decoupled.scala 361:21]
    .clock(q_109_clock),
    .reset(q_109_reset),
    .io_enq_ready(q_109_io_enq_ready),
    .io_enq_valid(q_109_io_enq_valid),
    .io_enq_bits(q_109_io_enq_bits),
    .io_deq_ready(q_109_io_deq_ready),
    .io_deq_valid(q_109_io_deq_valid),
    .io_deq_bits(q_109_io_deq_bits)
  );
  Queue q_110 ( // @[Decoupled.scala 361:21]
    .clock(q_110_clock),
    .reset(q_110_reset),
    .io_enq_ready(q_110_io_enq_ready),
    .io_enq_valid(q_110_io_enq_valid),
    .io_enq_bits(q_110_io_enq_bits),
    .io_deq_ready(q_110_io_deq_ready),
    .io_deq_valid(q_110_io_deq_valid),
    .io_deq_bits(q_110_io_deq_bits)
  );
  Queue q_111 ( // @[Decoupled.scala 361:21]
    .clock(q_111_clock),
    .reset(q_111_reset),
    .io_enq_ready(q_111_io_enq_ready),
    .io_enq_valid(q_111_io_enq_valid),
    .io_enq_bits(q_111_io_enq_bits),
    .io_deq_ready(q_111_io_deq_ready),
    .io_deq_valid(q_111_io_deq_valid),
    .io_deq_bits(q_111_io_deq_bits)
  );
  Queue q_112 ( // @[Decoupled.scala 361:21]
    .clock(q_112_clock),
    .reset(q_112_reset),
    .io_enq_ready(q_112_io_enq_ready),
    .io_enq_valid(q_112_io_enq_valid),
    .io_enq_bits(q_112_io_enq_bits),
    .io_deq_ready(q_112_io_deq_ready),
    .io_deq_valid(q_112_io_deq_valid),
    .io_deq_bits(q_112_io_deq_bits)
  );
  Queue q_113 ( // @[Decoupled.scala 361:21]
    .clock(q_113_clock),
    .reset(q_113_reset),
    .io_enq_ready(q_113_io_enq_ready),
    .io_enq_valid(q_113_io_enq_valid),
    .io_enq_bits(q_113_io_enq_bits),
    .io_deq_ready(q_113_io_deq_ready),
    .io_deq_valid(q_113_io_deq_valid),
    .io_deq_bits(q_113_io_deq_bits)
  );
  Queue q_114 ( // @[Decoupled.scala 361:21]
    .clock(q_114_clock),
    .reset(q_114_reset),
    .io_enq_ready(q_114_io_enq_ready),
    .io_enq_valid(q_114_io_enq_valid),
    .io_enq_bits(q_114_io_enq_bits),
    .io_deq_ready(q_114_io_deq_ready),
    .io_deq_valid(q_114_io_deq_valid),
    .io_deq_bits(q_114_io_deq_bits)
  );
  Queue q_115 ( // @[Decoupled.scala 361:21]
    .clock(q_115_clock),
    .reset(q_115_reset),
    .io_enq_ready(q_115_io_enq_ready),
    .io_enq_valid(q_115_io_enq_valid),
    .io_enq_bits(q_115_io_enq_bits),
    .io_deq_ready(q_115_io_deq_ready),
    .io_deq_valid(q_115_io_deq_valid),
    .io_deq_bits(q_115_io_deq_bits)
  );
  Queue q_116 ( // @[Decoupled.scala 361:21]
    .clock(q_116_clock),
    .reset(q_116_reset),
    .io_enq_ready(q_116_io_enq_ready),
    .io_enq_valid(q_116_io_enq_valid),
    .io_enq_bits(q_116_io_enq_bits),
    .io_deq_ready(q_116_io_deq_ready),
    .io_deq_valid(q_116_io_deq_valid),
    .io_deq_bits(q_116_io_deq_bits)
  );
  Queue q_117 ( // @[Decoupled.scala 361:21]
    .clock(q_117_clock),
    .reset(q_117_reset),
    .io_enq_ready(q_117_io_enq_ready),
    .io_enq_valid(q_117_io_enq_valid),
    .io_enq_bits(q_117_io_enq_bits),
    .io_deq_ready(q_117_io_deq_ready),
    .io_deq_valid(q_117_io_deq_valid),
    .io_deq_bits(q_117_io_deq_bits)
  );
  Queue q_118 ( // @[Decoupled.scala 361:21]
    .clock(q_118_clock),
    .reset(q_118_reset),
    .io_enq_ready(q_118_io_enq_ready),
    .io_enq_valid(q_118_io_enq_valid),
    .io_enq_bits(q_118_io_enq_bits),
    .io_deq_ready(q_118_io_deq_ready),
    .io_deq_valid(q_118_io_deq_valid),
    .io_deq_bits(q_118_io_deq_bits)
  );
  Queue q_119 ( // @[Decoupled.scala 361:21]
    .clock(q_119_clock),
    .reset(q_119_reset),
    .io_enq_ready(q_119_io_enq_ready),
    .io_enq_valid(q_119_io_enq_valid),
    .io_enq_bits(q_119_io_enq_bits),
    .io_deq_ready(q_119_io_deq_ready),
    .io_deq_valid(q_119_io_deq_valid),
    .io_deq_bits(q_119_io_deq_bits)
  );
  Queue q_120 ( // @[Decoupled.scala 361:21]
    .clock(q_120_clock),
    .reset(q_120_reset),
    .io_enq_ready(q_120_io_enq_ready),
    .io_enq_valid(q_120_io_enq_valid),
    .io_enq_bits(q_120_io_enq_bits),
    .io_deq_ready(q_120_io_deq_ready),
    .io_deq_valid(q_120_io_deq_valid),
    .io_deq_bits(q_120_io_deq_bits)
  );
  Queue q_121 ( // @[Decoupled.scala 361:21]
    .clock(q_121_clock),
    .reset(q_121_reset),
    .io_enq_ready(q_121_io_enq_ready),
    .io_enq_valid(q_121_io_enq_valid),
    .io_enq_bits(q_121_io_enq_bits),
    .io_deq_ready(q_121_io_deq_ready),
    .io_deq_valid(q_121_io_deq_valid),
    .io_deq_bits(q_121_io_deq_bits)
  );
  Queue q_122 ( // @[Decoupled.scala 361:21]
    .clock(q_122_clock),
    .reset(q_122_reset),
    .io_enq_ready(q_122_io_enq_ready),
    .io_enq_valid(q_122_io_enq_valid),
    .io_enq_bits(q_122_io_enq_bits),
    .io_deq_ready(q_122_io_deq_ready),
    .io_deq_valid(q_122_io_deq_valid),
    .io_deq_bits(q_122_io_deq_bits)
  );
  Queue q_123 ( // @[Decoupled.scala 361:21]
    .clock(q_123_clock),
    .reset(q_123_reset),
    .io_enq_ready(q_123_io_enq_ready),
    .io_enq_valid(q_123_io_enq_valid),
    .io_enq_bits(q_123_io_enq_bits),
    .io_deq_ready(q_123_io_deq_ready),
    .io_deq_valid(q_123_io_deq_valid),
    .io_deq_bits(q_123_io_deq_bits)
  );
  Queue q_124 ( // @[Decoupled.scala 361:21]
    .clock(q_124_clock),
    .reset(q_124_reset),
    .io_enq_ready(q_124_io_enq_ready),
    .io_enq_valid(q_124_io_enq_valid),
    .io_enq_bits(q_124_io_enq_bits),
    .io_deq_ready(q_124_io_deq_ready),
    .io_deq_valid(q_124_io_deq_valid),
    .io_deq_bits(q_124_io_deq_bits)
  );
  Queue q_125 ( // @[Decoupled.scala 361:21]
    .clock(q_125_clock),
    .reset(q_125_reset),
    .io_enq_ready(q_125_io_enq_ready),
    .io_enq_valid(q_125_io_enq_valid),
    .io_enq_bits(q_125_io_enq_bits),
    .io_deq_ready(q_125_io_deq_ready),
    .io_deq_valid(q_125_io_deq_valid),
    .io_deq_bits(q_125_io_deq_bits)
  );
  Queue q_126 ( // @[Decoupled.scala 361:21]
    .clock(q_126_clock),
    .reset(q_126_reset),
    .io_enq_ready(q_126_io_enq_ready),
    .io_enq_valid(q_126_io_enq_valid),
    .io_enq_bits(q_126_io_enq_bits),
    .io_deq_ready(q_126_io_deq_ready),
    .io_deq_valid(q_126_io_deq_valid),
    .io_deq_bits(q_126_io_deq_bits)
  );
  Queue q_127 ( // @[Decoupled.scala 361:21]
    .clock(q_127_clock),
    .reset(q_127_reset),
    .io_enq_ready(q_127_io_enq_ready),
    .io_enq_valid(q_127_io_enq_valid),
    .io_enq_bits(q_127_io_enq_bits),
    .io_deq_ready(q_127_io_deq_ready),
    .io_deq_valid(q_127_io_deq_valid),
    .io_deq_bits(q_127_io_deq_bits)
  );
  Queue q_128 ( // @[Decoupled.scala 361:21]
    .clock(q_128_clock),
    .reset(q_128_reset),
    .io_enq_ready(q_128_io_enq_ready),
    .io_enq_valid(q_128_io_enq_valid),
    .io_enq_bits(q_128_io_enq_bits),
    .io_deq_ready(q_128_io_deq_ready),
    .io_deq_valid(q_128_io_deq_valid),
    .io_deq_bits(q_128_io_deq_bits)
  );
  Queue q_129 ( // @[Decoupled.scala 361:21]
    .clock(q_129_clock),
    .reset(q_129_reset),
    .io_enq_ready(q_129_io_enq_ready),
    .io_enq_valid(q_129_io_enq_valid),
    .io_enq_bits(q_129_io_enq_bits),
    .io_deq_ready(q_129_io_deq_ready),
    .io_deq_valid(q_129_io_deq_valid),
    .io_deq_bits(q_129_io_deq_bits)
  );
  Queue q_130 ( // @[Decoupled.scala 361:21]
    .clock(q_130_clock),
    .reset(q_130_reset),
    .io_enq_ready(q_130_io_enq_ready),
    .io_enq_valid(q_130_io_enq_valid),
    .io_enq_bits(q_130_io_enq_bits),
    .io_deq_ready(q_130_io_deq_ready),
    .io_deq_valid(q_130_io_deq_valid),
    .io_deq_bits(q_130_io_deq_bits)
  );
  Queue q_131 ( // @[Decoupled.scala 361:21]
    .clock(q_131_clock),
    .reset(q_131_reset),
    .io_enq_ready(q_131_io_enq_ready),
    .io_enq_valid(q_131_io_enq_valid),
    .io_enq_bits(q_131_io_enq_bits),
    .io_deq_ready(q_131_io_deq_ready),
    .io_deq_valid(q_131_io_deq_valid),
    .io_deq_bits(q_131_io_deq_bits)
  );
  Queue q_132 ( // @[Decoupled.scala 361:21]
    .clock(q_132_clock),
    .reset(q_132_reset),
    .io_enq_ready(q_132_io_enq_ready),
    .io_enq_valid(q_132_io_enq_valid),
    .io_enq_bits(q_132_io_enq_bits),
    .io_deq_ready(q_132_io_deq_ready),
    .io_deq_valid(q_132_io_deq_valid),
    .io_deq_bits(q_132_io_deq_bits)
  );
  Queue q_133 ( // @[Decoupled.scala 361:21]
    .clock(q_133_clock),
    .reset(q_133_reset),
    .io_enq_ready(q_133_io_enq_ready),
    .io_enq_valid(q_133_io_enq_valid),
    .io_enq_bits(q_133_io_enq_bits),
    .io_deq_ready(q_133_io_deq_ready),
    .io_deq_valid(q_133_io_deq_valid),
    .io_deq_bits(q_133_io_deq_bits)
  );
  Queue q_134 ( // @[Decoupled.scala 361:21]
    .clock(q_134_clock),
    .reset(q_134_reset),
    .io_enq_ready(q_134_io_enq_ready),
    .io_enq_valid(q_134_io_enq_valid),
    .io_enq_bits(q_134_io_enq_bits),
    .io_deq_ready(q_134_io_deq_ready),
    .io_deq_valid(q_134_io_deq_valid),
    .io_deq_bits(q_134_io_deq_bits)
  );
  Queue q_135 ( // @[Decoupled.scala 361:21]
    .clock(q_135_clock),
    .reset(q_135_reset),
    .io_enq_ready(q_135_io_enq_ready),
    .io_enq_valid(q_135_io_enq_valid),
    .io_enq_bits(q_135_io_enq_bits),
    .io_deq_ready(q_135_io_deq_ready),
    .io_deq_valid(q_135_io_deq_valid),
    .io_deq_bits(q_135_io_deq_bits)
  );
  Queue q_136 ( // @[Decoupled.scala 361:21]
    .clock(q_136_clock),
    .reset(q_136_reset),
    .io_enq_ready(q_136_io_enq_ready),
    .io_enq_valid(q_136_io_enq_valid),
    .io_enq_bits(q_136_io_enq_bits),
    .io_deq_ready(q_136_io_deq_ready),
    .io_deq_valid(q_136_io_deq_valid),
    .io_deq_bits(q_136_io_deq_bits)
  );
  Queue q_137 ( // @[Decoupled.scala 361:21]
    .clock(q_137_clock),
    .reset(q_137_reset),
    .io_enq_ready(q_137_io_enq_ready),
    .io_enq_valid(q_137_io_enq_valid),
    .io_enq_bits(q_137_io_enq_bits),
    .io_deq_ready(q_137_io_deq_ready),
    .io_deq_valid(q_137_io_deq_valid),
    .io_deq_bits(q_137_io_deq_bits)
  );
  Queue q_138 ( // @[Decoupled.scala 361:21]
    .clock(q_138_clock),
    .reset(q_138_reset),
    .io_enq_ready(q_138_io_enq_ready),
    .io_enq_valid(q_138_io_enq_valid),
    .io_enq_bits(q_138_io_enq_bits),
    .io_deq_ready(q_138_io_deq_ready),
    .io_deq_valid(q_138_io_deq_valid),
    .io_deq_bits(q_138_io_deq_bits)
  );
  Queue q_139 ( // @[Decoupled.scala 361:21]
    .clock(q_139_clock),
    .reset(q_139_reset),
    .io_enq_ready(q_139_io_enq_ready),
    .io_enq_valid(q_139_io_enq_valid),
    .io_enq_bits(q_139_io_enq_bits),
    .io_deq_ready(q_139_io_deq_ready),
    .io_deq_valid(q_139_io_deq_valid),
    .io_deq_bits(q_139_io_deq_bits)
  );
  Queue q_140 ( // @[Decoupled.scala 361:21]
    .clock(q_140_clock),
    .reset(q_140_reset),
    .io_enq_ready(q_140_io_enq_ready),
    .io_enq_valid(q_140_io_enq_valid),
    .io_enq_bits(q_140_io_enq_bits),
    .io_deq_ready(q_140_io_deq_ready),
    .io_deq_valid(q_140_io_deq_valid),
    .io_deq_bits(q_140_io_deq_bits)
  );
  Queue q_141 ( // @[Decoupled.scala 361:21]
    .clock(q_141_clock),
    .reset(q_141_reset),
    .io_enq_ready(q_141_io_enq_ready),
    .io_enq_valid(q_141_io_enq_valid),
    .io_enq_bits(q_141_io_enq_bits),
    .io_deq_ready(q_141_io_deq_ready),
    .io_deq_valid(q_141_io_deq_valid),
    .io_deq_bits(q_141_io_deq_bits)
  );
  Queue q_142 ( // @[Decoupled.scala 361:21]
    .clock(q_142_clock),
    .reset(q_142_reset),
    .io_enq_ready(q_142_io_enq_ready),
    .io_enq_valid(q_142_io_enq_valid),
    .io_enq_bits(q_142_io_enq_bits),
    .io_deq_ready(q_142_io_deq_ready),
    .io_deq_valid(q_142_io_deq_valid),
    .io_deq_bits(q_142_io_deq_bits)
  );
  Queue q_143 ( // @[Decoupled.scala 361:21]
    .clock(q_143_clock),
    .reset(q_143_reset),
    .io_enq_ready(q_143_io_enq_ready),
    .io_enq_valid(q_143_io_enq_valid),
    .io_enq_bits(q_143_io_enq_bits),
    .io_deq_ready(q_143_io_deq_ready),
    .io_deq_valid(q_143_io_deq_valid),
    .io_deq_bits(q_143_io_deq_bits)
  );
  Queue q_144 ( // @[Decoupled.scala 361:21]
    .clock(q_144_clock),
    .reset(q_144_reset),
    .io_enq_ready(q_144_io_enq_ready),
    .io_enq_valid(q_144_io_enq_valid),
    .io_enq_bits(q_144_io_enq_bits),
    .io_deq_ready(q_144_io_deq_ready),
    .io_deq_valid(q_144_io_deq_valid),
    .io_deq_bits(q_144_io_deq_bits)
  );
  Queue q_145 ( // @[Decoupled.scala 361:21]
    .clock(q_145_clock),
    .reset(q_145_reset),
    .io_enq_ready(q_145_io_enq_ready),
    .io_enq_valid(q_145_io_enq_valid),
    .io_enq_bits(q_145_io_enq_bits),
    .io_deq_ready(q_145_io_deq_ready),
    .io_deq_valid(q_145_io_deq_valid),
    .io_deq_bits(q_145_io_deq_bits)
  );
  Queue q_146 ( // @[Decoupled.scala 361:21]
    .clock(q_146_clock),
    .reset(q_146_reset),
    .io_enq_ready(q_146_io_enq_ready),
    .io_enq_valid(q_146_io_enq_valid),
    .io_enq_bits(q_146_io_enq_bits),
    .io_deq_ready(q_146_io_deq_ready),
    .io_deq_valid(q_146_io_deq_valid),
    .io_deq_bits(q_146_io_deq_bits)
  );
  Queue q_147 ( // @[Decoupled.scala 361:21]
    .clock(q_147_clock),
    .reset(q_147_reset),
    .io_enq_ready(q_147_io_enq_ready),
    .io_enq_valid(q_147_io_enq_valid),
    .io_enq_bits(q_147_io_enq_bits),
    .io_deq_ready(q_147_io_deq_ready),
    .io_deq_valid(q_147_io_deq_valid),
    .io_deq_bits(q_147_io_deq_bits)
  );
  Queue q_148 ( // @[Decoupled.scala 361:21]
    .clock(q_148_clock),
    .reset(q_148_reset),
    .io_enq_ready(q_148_io_enq_ready),
    .io_enq_valid(q_148_io_enq_valid),
    .io_enq_bits(q_148_io_enq_bits),
    .io_deq_ready(q_148_io_deq_ready),
    .io_deq_valid(q_148_io_deq_valid),
    .io_deq_bits(q_148_io_deq_bits)
  );
  Queue q_149 ( // @[Decoupled.scala 361:21]
    .clock(q_149_clock),
    .reset(q_149_reset),
    .io_enq_ready(q_149_io_enq_ready),
    .io_enq_valid(q_149_io_enq_valid),
    .io_enq_bits(q_149_io_enq_bits),
    .io_deq_ready(q_149_io_deq_ready),
    .io_deq_valid(q_149_io_deq_valid),
    .io_deq_bits(q_149_io_deq_bits)
  );
  Queue q_150 ( // @[Decoupled.scala 361:21]
    .clock(q_150_clock),
    .reset(q_150_reset),
    .io_enq_ready(q_150_io_enq_ready),
    .io_enq_valid(q_150_io_enq_valid),
    .io_enq_bits(q_150_io_enq_bits),
    .io_deq_ready(q_150_io_deq_ready),
    .io_deq_valid(q_150_io_deq_valid),
    .io_deq_bits(q_150_io_deq_bits)
  );
  Queue q_151 ( // @[Decoupled.scala 361:21]
    .clock(q_151_clock),
    .reset(q_151_reset),
    .io_enq_ready(q_151_io_enq_ready),
    .io_enq_valid(q_151_io_enq_valid),
    .io_enq_bits(q_151_io_enq_bits),
    .io_deq_ready(q_151_io_deq_ready),
    .io_deq_valid(q_151_io_deq_valid),
    .io_deq_bits(q_151_io_deq_bits)
  );
  Queue q_152 ( // @[Decoupled.scala 361:21]
    .clock(q_152_clock),
    .reset(q_152_reset),
    .io_enq_ready(q_152_io_enq_ready),
    .io_enq_valid(q_152_io_enq_valid),
    .io_enq_bits(q_152_io_enq_bits),
    .io_deq_ready(q_152_io_deq_ready),
    .io_deq_valid(q_152_io_deq_valid),
    .io_deq_bits(q_152_io_deq_bits)
  );
  Queue q_153 ( // @[Decoupled.scala 361:21]
    .clock(q_153_clock),
    .reset(q_153_reset),
    .io_enq_ready(q_153_io_enq_ready),
    .io_enq_valid(q_153_io_enq_valid),
    .io_enq_bits(q_153_io_enq_bits),
    .io_deq_ready(q_153_io_deq_ready),
    .io_deq_valid(q_153_io_deq_valid),
    .io_deq_bits(q_153_io_deq_bits)
  );
  Queue q_154 ( // @[Decoupled.scala 361:21]
    .clock(q_154_clock),
    .reset(q_154_reset),
    .io_enq_ready(q_154_io_enq_ready),
    .io_enq_valid(q_154_io_enq_valid),
    .io_enq_bits(q_154_io_enq_bits),
    .io_deq_ready(q_154_io_deq_ready),
    .io_deq_valid(q_154_io_deq_valid),
    .io_deq_bits(q_154_io_deq_bits)
  );
  Queue q_155 ( // @[Decoupled.scala 361:21]
    .clock(q_155_clock),
    .reset(q_155_reset),
    .io_enq_ready(q_155_io_enq_ready),
    .io_enq_valid(q_155_io_enq_valid),
    .io_enq_bits(q_155_io_enq_bits),
    .io_deq_ready(q_155_io_deq_ready),
    .io_deq_valid(q_155_io_deq_valid),
    .io_deq_bits(q_155_io_deq_bits)
  );
  Queue q_156 ( // @[Decoupled.scala 361:21]
    .clock(q_156_clock),
    .reset(q_156_reset),
    .io_enq_ready(q_156_io_enq_ready),
    .io_enq_valid(q_156_io_enq_valid),
    .io_enq_bits(q_156_io_enq_bits),
    .io_deq_ready(q_156_io_deq_ready),
    .io_deq_valid(q_156_io_deq_valid),
    .io_deq_bits(q_156_io_deq_bits)
  );
  Queue q_157 ( // @[Decoupled.scala 361:21]
    .clock(q_157_clock),
    .reset(q_157_reset),
    .io_enq_ready(q_157_io_enq_ready),
    .io_enq_valid(q_157_io_enq_valid),
    .io_enq_bits(q_157_io_enq_bits),
    .io_deq_ready(q_157_io_deq_ready),
    .io_deq_valid(q_157_io_deq_valid),
    .io_deq_bits(q_157_io_deq_bits)
  );
  Queue q_158 ( // @[Decoupled.scala 361:21]
    .clock(q_158_clock),
    .reset(q_158_reset),
    .io_enq_ready(q_158_io_enq_ready),
    .io_enq_valid(q_158_io_enq_valid),
    .io_enq_bits(q_158_io_enq_bits),
    .io_deq_ready(q_158_io_deq_ready),
    .io_deq_valid(q_158_io_deq_valid),
    .io_deq_bits(q_158_io_deq_bits)
  );
  Queue q_159 ( // @[Decoupled.scala 361:21]
    .clock(q_159_clock),
    .reset(q_159_reset),
    .io_enq_ready(q_159_io_enq_ready),
    .io_enq_valid(q_159_io_enq_valid),
    .io_enq_bits(q_159_io_enq_bits),
    .io_deq_ready(q_159_io_deq_ready),
    .io_deq_valid(q_159_io_deq_valid),
    .io_deq_bits(q_159_io_deq_bits)
  );
  Queue q_160 ( // @[Decoupled.scala 361:21]
    .clock(q_160_clock),
    .reset(q_160_reset),
    .io_enq_ready(q_160_io_enq_ready),
    .io_enq_valid(q_160_io_enq_valid),
    .io_enq_bits(q_160_io_enq_bits),
    .io_deq_ready(q_160_io_deq_ready),
    .io_deq_valid(q_160_io_deq_valid),
    .io_deq_bits(q_160_io_deq_bits)
  );
  Queue q_161 ( // @[Decoupled.scala 361:21]
    .clock(q_161_clock),
    .reset(q_161_reset),
    .io_enq_ready(q_161_io_enq_ready),
    .io_enq_valid(q_161_io_enq_valid),
    .io_enq_bits(q_161_io_enq_bits),
    .io_deq_ready(q_161_io_deq_ready),
    .io_deq_valid(q_161_io_deq_valid),
    .io_deq_bits(q_161_io_deq_bits)
  );
  Queue q_162 ( // @[Decoupled.scala 361:21]
    .clock(q_162_clock),
    .reset(q_162_reset),
    .io_enq_ready(q_162_io_enq_ready),
    .io_enq_valid(q_162_io_enq_valid),
    .io_enq_bits(q_162_io_enq_bits),
    .io_deq_ready(q_162_io_deq_ready),
    .io_deq_valid(q_162_io_deq_valid),
    .io_deq_bits(q_162_io_deq_bits)
  );
  Queue q_163 ( // @[Decoupled.scala 361:21]
    .clock(q_163_clock),
    .reset(q_163_reset),
    .io_enq_ready(q_163_io_enq_ready),
    .io_enq_valid(q_163_io_enq_valid),
    .io_enq_bits(q_163_io_enq_bits),
    .io_deq_ready(q_163_io_deq_ready),
    .io_deq_valid(q_163_io_deq_valid),
    .io_deq_bits(q_163_io_deq_bits)
  );
  Queue q_164 ( // @[Decoupled.scala 361:21]
    .clock(q_164_clock),
    .reset(q_164_reset),
    .io_enq_ready(q_164_io_enq_ready),
    .io_enq_valid(q_164_io_enq_valid),
    .io_enq_bits(q_164_io_enq_bits),
    .io_deq_ready(q_164_io_deq_ready),
    .io_deq_valid(q_164_io_deq_valid),
    .io_deq_bits(q_164_io_deq_bits)
  );
  Queue q_165 ( // @[Decoupled.scala 361:21]
    .clock(q_165_clock),
    .reset(q_165_reset),
    .io_enq_ready(q_165_io_enq_ready),
    .io_enq_valid(q_165_io_enq_valid),
    .io_enq_bits(q_165_io_enq_bits),
    .io_deq_ready(q_165_io_deq_ready),
    .io_deq_valid(q_165_io_deq_valid),
    .io_deq_bits(q_165_io_deq_bits)
  );
  Queue q_166 ( // @[Decoupled.scala 361:21]
    .clock(q_166_clock),
    .reset(q_166_reset),
    .io_enq_ready(q_166_io_enq_ready),
    .io_enq_valid(q_166_io_enq_valid),
    .io_enq_bits(q_166_io_enq_bits),
    .io_deq_ready(q_166_io_deq_ready),
    .io_deq_valid(q_166_io_deq_valid),
    .io_deq_bits(q_166_io_deq_bits)
  );
  Queue q_167 ( // @[Decoupled.scala 361:21]
    .clock(q_167_clock),
    .reset(q_167_reset),
    .io_enq_ready(q_167_io_enq_ready),
    .io_enq_valid(q_167_io_enq_valid),
    .io_enq_bits(q_167_io_enq_bits),
    .io_deq_ready(q_167_io_deq_ready),
    .io_deq_valid(q_167_io_deq_valid),
    .io_deq_bits(q_167_io_deq_bits)
  );
  Queue q_168 ( // @[Decoupled.scala 361:21]
    .clock(q_168_clock),
    .reset(q_168_reset),
    .io_enq_ready(q_168_io_enq_ready),
    .io_enq_valid(q_168_io_enq_valid),
    .io_enq_bits(q_168_io_enq_bits),
    .io_deq_ready(q_168_io_deq_ready),
    .io_deq_valid(q_168_io_deq_valid),
    .io_deq_bits(q_168_io_deq_bits)
  );
  Queue q_169 ( // @[Decoupled.scala 361:21]
    .clock(q_169_clock),
    .reset(q_169_reset),
    .io_enq_ready(q_169_io_enq_ready),
    .io_enq_valid(q_169_io_enq_valid),
    .io_enq_bits(q_169_io_enq_bits),
    .io_deq_ready(q_169_io_deq_ready),
    .io_deq_valid(q_169_io_deq_valid),
    .io_deq_bits(q_169_io_deq_bits)
  );
  Queue q_170 ( // @[Decoupled.scala 361:21]
    .clock(q_170_clock),
    .reset(q_170_reset),
    .io_enq_ready(q_170_io_enq_ready),
    .io_enq_valid(q_170_io_enq_valid),
    .io_enq_bits(q_170_io_enq_bits),
    .io_deq_ready(q_170_io_deq_ready),
    .io_deq_valid(q_170_io_deq_valid),
    .io_deq_bits(q_170_io_deq_bits)
  );
  Queue q_171 ( // @[Decoupled.scala 361:21]
    .clock(q_171_clock),
    .reset(q_171_reset),
    .io_enq_ready(q_171_io_enq_ready),
    .io_enq_valid(q_171_io_enq_valid),
    .io_enq_bits(q_171_io_enq_bits),
    .io_deq_ready(q_171_io_deq_ready),
    .io_deq_valid(q_171_io_deq_valid),
    .io_deq_bits(q_171_io_deq_bits)
  );
  Queue q_172 ( // @[Decoupled.scala 361:21]
    .clock(q_172_clock),
    .reset(q_172_reset),
    .io_enq_ready(q_172_io_enq_ready),
    .io_enq_valid(q_172_io_enq_valid),
    .io_enq_bits(q_172_io_enq_bits),
    .io_deq_ready(q_172_io_deq_ready),
    .io_deq_valid(q_172_io_deq_valid),
    .io_deq_bits(q_172_io_deq_bits)
  );
  Queue q_173 ( // @[Decoupled.scala 361:21]
    .clock(q_173_clock),
    .reset(q_173_reset),
    .io_enq_ready(q_173_io_enq_ready),
    .io_enq_valid(q_173_io_enq_valid),
    .io_enq_bits(q_173_io_enq_bits),
    .io_deq_ready(q_173_io_deq_ready),
    .io_deq_valid(q_173_io_deq_valid),
    .io_deq_bits(q_173_io_deq_bits)
  );
  Queue q_174 ( // @[Decoupled.scala 361:21]
    .clock(q_174_clock),
    .reset(q_174_reset),
    .io_enq_ready(q_174_io_enq_ready),
    .io_enq_valid(q_174_io_enq_valid),
    .io_enq_bits(q_174_io_enq_bits),
    .io_deq_ready(q_174_io_deq_ready),
    .io_deq_valid(q_174_io_deq_valid),
    .io_deq_bits(q_174_io_deq_bits)
  );
  Queue q_175 ( // @[Decoupled.scala 361:21]
    .clock(q_175_clock),
    .reset(q_175_reset),
    .io_enq_ready(q_175_io_enq_ready),
    .io_enq_valid(q_175_io_enq_valid),
    .io_enq_bits(q_175_io_enq_bits),
    .io_deq_ready(q_175_io_deq_ready),
    .io_deq_valid(q_175_io_deq_valid),
    .io_deq_bits(q_175_io_deq_bits)
  );
  Queue q_176 ( // @[Decoupled.scala 361:21]
    .clock(q_176_clock),
    .reset(q_176_reset),
    .io_enq_ready(q_176_io_enq_ready),
    .io_enq_valid(q_176_io_enq_valid),
    .io_enq_bits(q_176_io_enq_bits),
    .io_deq_ready(q_176_io_deq_ready),
    .io_deq_valid(q_176_io_deq_valid),
    .io_deq_bits(q_176_io_deq_bits)
  );
  Queue q_177 ( // @[Decoupled.scala 361:21]
    .clock(q_177_clock),
    .reset(q_177_reset),
    .io_enq_ready(q_177_io_enq_ready),
    .io_enq_valid(q_177_io_enq_valid),
    .io_enq_bits(q_177_io_enq_bits),
    .io_deq_ready(q_177_io_deq_ready),
    .io_deq_valid(q_177_io_deq_valid),
    .io_deq_bits(q_177_io_deq_bits)
  );
  Queue q_178 ( // @[Decoupled.scala 361:21]
    .clock(q_178_clock),
    .reset(q_178_reset),
    .io_enq_ready(q_178_io_enq_ready),
    .io_enq_valid(q_178_io_enq_valid),
    .io_enq_bits(q_178_io_enq_bits),
    .io_deq_ready(q_178_io_deq_ready),
    .io_deq_valid(q_178_io_deq_valid),
    .io_deq_bits(q_178_io_deq_bits)
  );
  Queue q_179 ( // @[Decoupled.scala 361:21]
    .clock(q_179_clock),
    .reset(q_179_reset),
    .io_enq_ready(q_179_io_enq_ready),
    .io_enq_valid(q_179_io_enq_valid),
    .io_enq_bits(q_179_io_enq_bits),
    .io_deq_ready(q_179_io_deq_ready),
    .io_deq_valid(q_179_io_deq_valid),
    .io_deq_bits(q_179_io_deq_bits)
  );
  Queue q_180 ( // @[Decoupled.scala 361:21]
    .clock(q_180_clock),
    .reset(q_180_reset),
    .io_enq_ready(q_180_io_enq_ready),
    .io_enq_valid(q_180_io_enq_valid),
    .io_enq_bits(q_180_io_enq_bits),
    .io_deq_ready(q_180_io_deq_ready),
    .io_deq_valid(q_180_io_deq_valid),
    .io_deq_bits(q_180_io_deq_bits)
  );
  Queue q_181 ( // @[Decoupled.scala 361:21]
    .clock(q_181_clock),
    .reset(q_181_reset),
    .io_enq_ready(q_181_io_enq_ready),
    .io_enq_valid(q_181_io_enq_valid),
    .io_enq_bits(q_181_io_enq_bits),
    .io_deq_ready(q_181_io_deq_ready),
    .io_deq_valid(q_181_io_deq_valid),
    .io_deq_bits(q_181_io_deq_bits)
  );
  Queue q_182 ( // @[Decoupled.scala 361:21]
    .clock(q_182_clock),
    .reset(q_182_reset),
    .io_enq_ready(q_182_io_enq_ready),
    .io_enq_valid(q_182_io_enq_valid),
    .io_enq_bits(q_182_io_enq_bits),
    .io_deq_ready(q_182_io_deq_ready),
    .io_deq_valid(q_182_io_deq_valid),
    .io_deq_bits(q_182_io_deq_bits)
  );
  Queue q_183 ( // @[Decoupled.scala 361:21]
    .clock(q_183_clock),
    .reset(q_183_reset),
    .io_enq_ready(q_183_io_enq_ready),
    .io_enq_valid(q_183_io_enq_valid),
    .io_enq_bits(q_183_io_enq_bits),
    .io_deq_ready(q_183_io_deq_ready),
    .io_deq_valid(q_183_io_deq_valid),
    .io_deq_bits(q_183_io_deq_bits)
  );
  Queue q_184 ( // @[Decoupled.scala 361:21]
    .clock(q_184_clock),
    .reset(q_184_reset),
    .io_enq_ready(q_184_io_enq_ready),
    .io_enq_valid(q_184_io_enq_valid),
    .io_enq_bits(q_184_io_enq_bits),
    .io_deq_ready(q_184_io_deq_ready),
    .io_deq_valid(q_184_io_deq_valid),
    .io_deq_bits(q_184_io_deq_bits)
  );
  Queue q_185 ( // @[Decoupled.scala 361:21]
    .clock(q_185_clock),
    .reset(q_185_reset),
    .io_enq_ready(q_185_io_enq_ready),
    .io_enq_valid(q_185_io_enq_valid),
    .io_enq_bits(q_185_io_enq_bits),
    .io_deq_ready(q_185_io_deq_ready),
    .io_deq_valid(q_185_io_deq_valid),
    .io_deq_bits(q_185_io_deq_bits)
  );
  Queue q_186 ( // @[Decoupled.scala 361:21]
    .clock(q_186_clock),
    .reset(q_186_reset),
    .io_enq_ready(q_186_io_enq_ready),
    .io_enq_valid(q_186_io_enq_valid),
    .io_enq_bits(q_186_io_enq_bits),
    .io_deq_ready(q_186_io_deq_ready),
    .io_deq_valid(q_186_io_deq_valid),
    .io_deq_bits(q_186_io_deq_bits)
  );
  Queue q_187 ( // @[Decoupled.scala 361:21]
    .clock(q_187_clock),
    .reset(q_187_reset),
    .io_enq_ready(q_187_io_enq_ready),
    .io_enq_valid(q_187_io_enq_valid),
    .io_enq_bits(q_187_io_enq_bits),
    .io_deq_ready(q_187_io_deq_ready),
    .io_deq_valid(q_187_io_deq_valid),
    .io_deq_bits(q_187_io_deq_bits)
  );
  Queue q_188 ( // @[Decoupled.scala 361:21]
    .clock(q_188_clock),
    .reset(q_188_reset),
    .io_enq_ready(q_188_io_enq_ready),
    .io_enq_valid(q_188_io_enq_valid),
    .io_enq_bits(q_188_io_enq_bits),
    .io_deq_ready(q_188_io_deq_ready),
    .io_deq_valid(q_188_io_deq_valid),
    .io_deq_bits(q_188_io_deq_bits)
  );
  Queue q_189 ( // @[Decoupled.scala 361:21]
    .clock(q_189_clock),
    .reset(q_189_reset),
    .io_enq_ready(q_189_io_enq_ready),
    .io_enq_valid(q_189_io_enq_valid),
    .io_enq_bits(q_189_io_enq_bits),
    .io_deq_ready(q_189_io_deq_ready),
    .io_deq_valid(q_189_io_deq_valid),
    .io_deq_bits(q_189_io_deq_bits)
  );
  Queue q_190 ( // @[Decoupled.scala 361:21]
    .clock(q_190_clock),
    .reset(q_190_reset),
    .io_enq_ready(q_190_io_enq_ready),
    .io_enq_valid(q_190_io_enq_valid),
    .io_enq_bits(q_190_io_enq_bits),
    .io_deq_ready(q_190_io_deq_ready),
    .io_deq_valid(q_190_io_deq_valid),
    .io_deq_bits(q_190_io_deq_bits)
  );
  Queue q_191 ( // @[Decoupled.scala 361:21]
    .clock(q_191_clock),
    .reset(q_191_reset),
    .io_enq_ready(q_191_io_enq_ready),
    .io_enq_valid(q_191_io_enq_valid),
    .io_enq_bits(q_191_io_enq_bits),
    .io_deq_ready(q_191_io_deq_ready),
    .io_deq_valid(q_191_io_deq_valid),
    .io_deq_bits(q_191_io_deq_bits)
  );
  Queue q_192 ( // @[Decoupled.scala 361:21]
    .clock(q_192_clock),
    .reset(q_192_reset),
    .io_enq_ready(q_192_io_enq_ready),
    .io_enq_valid(q_192_io_enq_valid),
    .io_enq_bits(q_192_io_enq_bits),
    .io_deq_ready(q_192_io_deq_ready),
    .io_deq_valid(q_192_io_deq_valid),
    .io_deq_bits(q_192_io_deq_bits)
  );
  Queue q_193 ( // @[Decoupled.scala 361:21]
    .clock(q_193_clock),
    .reset(q_193_reset),
    .io_enq_ready(q_193_io_enq_ready),
    .io_enq_valid(q_193_io_enq_valid),
    .io_enq_bits(q_193_io_enq_bits),
    .io_deq_ready(q_193_io_deq_ready),
    .io_deq_valid(q_193_io_deq_valid),
    .io_deq_bits(q_193_io_deq_bits)
  );
  Queue q_194 ( // @[Decoupled.scala 361:21]
    .clock(q_194_clock),
    .reset(q_194_reset),
    .io_enq_ready(q_194_io_enq_ready),
    .io_enq_valid(q_194_io_enq_valid),
    .io_enq_bits(q_194_io_enq_bits),
    .io_deq_ready(q_194_io_deq_ready),
    .io_deq_valid(q_194_io_deq_valid),
    .io_deq_bits(q_194_io_deq_bits)
  );
  Queue q_195 ( // @[Decoupled.scala 361:21]
    .clock(q_195_clock),
    .reset(q_195_reset),
    .io_enq_ready(q_195_io_enq_ready),
    .io_enq_valid(q_195_io_enq_valid),
    .io_enq_bits(q_195_io_enq_bits),
    .io_deq_ready(q_195_io_deq_ready),
    .io_deq_valid(q_195_io_deq_valid),
    .io_deq_bits(q_195_io_deq_bits)
  );
  Queue q_196 ( // @[Decoupled.scala 361:21]
    .clock(q_196_clock),
    .reset(q_196_reset),
    .io_enq_ready(q_196_io_enq_ready),
    .io_enq_valid(q_196_io_enq_valid),
    .io_enq_bits(q_196_io_enq_bits),
    .io_deq_ready(q_196_io_deq_ready),
    .io_deq_valid(q_196_io_deq_valid),
    .io_deq_bits(q_196_io_deq_bits)
  );
  Queue q_197 ( // @[Decoupled.scala 361:21]
    .clock(q_197_clock),
    .reset(q_197_reset),
    .io_enq_ready(q_197_io_enq_ready),
    .io_enq_valid(q_197_io_enq_valid),
    .io_enq_bits(q_197_io_enq_bits),
    .io_deq_ready(q_197_io_deq_ready),
    .io_deq_valid(q_197_io_deq_valid),
    .io_deq_bits(q_197_io_deq_bits)
  );
  Queue q_198 ( // @[Decoupled.scala 361:21]
    .clock(q_198_clock),
    .reset(q_198_reset),
    .io_enq_ready(q_198_io_enq_ready),
    .io_enq_valid(q_198_io_enq_valid),
    .io_enq_bits(q_198_io_enq_bits),
    .io_deq_ready(q_198_io_deq_ready),
    .io_deq_valid(q_198_io_deq_valid),
    .io_deq_bits(q_198_io_deq_bits)
  );
  Queue q_199 ( // @[Decoupled.scala 361:21]
    .clock(q_199_clock),
    .reset(q_199_reset),
    .io_enq_ready(q_199_io_enq_ready),
    .io_enq_valid(q_199_io_enq_valid),
    .io_enq_bits(q_199_io_enq_bits),
    .io_deq_ready(q_199_io_deq_ready),
    .io_deq_valid(q_199_io_deq_valid),
    .io_deq_bits(q_199_io_deq_bits)
  );
  Queue q_200 ( // @[Decoupled.scala 361:21]
    .clock(q_200_clock),
    .reset(q_200_reset),
    .io_enq_ready(q_200_io_enq_ready),
    .io_enq_valid(q_200_io_enq_valid),
    .io_enq_bits(q_200_io_enq_bits),
    .io_deq_ready(q_200_io_deq_ready),
    .io_deq_valid(q_200_io_deq_valid),
    .io_deq_bits(q_200_io_deq_bits)
  );
  Queue q_201 ( // @[Decoupled.scala 361:21]
    .clock(q_201_clock),
    .reset(q_201_reset),
    .io_enq_ready(q_201_io_enq_ready),
    .io_enq_valid(q_201_io_enq_valid),
    .io_enq_bits(q_201_io_enq_bits),
    .io_deq_ready(q_201_io_deq_ready),
    .io_deq_valid(q_201_io_deq_valid),
    .io_deq_bits(q_201_io_deq_bits)
  );
  Queue q_202 ( // @[Decoupled.scala 361:21]
    .clock(q_202_clock),
    .reset(q_202_reset),
    .io_enq_ready(q_202_io_enq_ready),
    .io_enq_valid(q_202_io_enq_valid),
    .io_enq_bits(q_202_io_enq_bits),
    .io_deq_ready(q_202_io_deq_ready),
    .io_deq_valid(q_202_io_deq_valid),
    .io_deq_bits(q_202_io_deq_bits)
  );
  Queue q_203 ( // @[Decoupled.scala 361:21]
    .clock(q_203_clock),
    .reset(q_203_reset),
    .io_enq_ready(q_203_io_enq_ready),
    .io_enq_valid(q_203_io_enq_valid),
    .io_enq_bits(q_203_io_enq_bits),
    .io_deq_ready(q_203_io_deq_ready),
    .io_deq_valid(q_203_io_deq_valid),
    .io_deq_bits(q_203_io_deq_bits)
  );
  Queue q_204 ( // @[Decoupled.scala 361:21]
    .clock(q_204_clock),
    .reset(q_204_reset),
    .io_enq_ready(q_204_io_enq_ready),
    .io_enq_valid(q_204_io_enq_valid),
    .io_enq_bits(q_204_io_enq_bits),
    .io_deq_ready(q_204_io_deq_ready),
    .io_deq_valid(q_204_io_deq_valid),
    .io_deq_bits(q_204_io_deq_bits)
  );
  Queue q_205 ( // @[Decoupled.scala 361:21]
    .clock(q_205_clock),
    .reset(q_205_reset),
    .io_enq_ready(q_205_io_enq_ready),
    .io_enq_valid(q_205_io_enq_valid),
    .io_enq_bits(q_205_io_enq_bits),
    .io_deq_ready(q_205_io_deq_ready),
    .io_deq_valid(q_205_io_deq_valid),
    .io_deq_bits(q_205_io_deq_bits)
  );
  Queue q_206 ( // @[Decoupled.scala 361:21]
    .clock(q_206_clock),
    .reset(q_206_reset),
    .io_enq_ready(q_206_io_enq_ready),
    .io_enq_valid(q_206_io_enq_valid),
    .io_enq_bits(q_206_io_enq_bits),
    .io_deq_ready(q_206_io_deq_ready),
    .io_deq_valid(q_206_io_deq_valid),
    .io_deq_bits(q_206_io_deq_bits)
  );
  Queue q_207 ( // @[Decoupled.scala 361:21]
    .clock(q_207_clock),
    .reset(q_207_reset),
    .io_enq_ready(q_207_io_enq_ready),
    .io_enq_valid(q_207_io_enq_valid),
    .io_enq_bits(q_207_io_enq_bits),
    .io_deq_ready(q_207_io_deq_ready),
    .io_deq_valid(q_207_io_deq_valid),
    .io_deq_bits(q_207_io_deq_bits)
  );
  Queue q_208 ( // @[Decoupled.scala 361:21]
    .clock(q_208_clock),
    .reset(q_208_reset),
    .io_enq_ready(q_208_io_enq_ready),
    .io_enq_valid(q_208_io_enq_valid),
    .io_enq_bits(q_208_io_enq_bits),
    .io_deq_ready(q_208_io_deq_ready),
    .io_deq_valid(q_208_io_deq_valid),
    .io_deq_bits(q_208_io_deq_bits)
  );
  Queue q_209 ( // @[Decoupled.scala 361:21]
    .clock(q_209_clock),
    .reset(q_209_reset),
    .io_enq_ready(q_209_io_enq_ready),
    .io_enq_valid(q_209_io_enq_valid),
    .io_enq_bits(q_209_io_enq_bits),
    .io_deq_ready(q_209_io_deq_ready),
    .io_deq_valid(q_209_io_deq_valid),
    .io_deq_bits(q_209_io_deq_bits)
  );
  Queue q_210 ( // @[Decoupled.scala 361:21]
    .clock(q_210_clock),
    .reset(q_210_reset),
    .io_enq_ready(q_210_io_enq_ready),
    .io_enq_valid(q_210_io_enq_valid),
    .io_enq_bits(q_210_io_enq_bits),
    .io_deq_ready(q_210_io_deq_ready),
    .io_deq_valid(q_210_io_deq_valid),
    .io_deq_bits(q_210_io_deq_bits)
  );
  Queue q_211 ( // @[Decoupled.scala 361:21]
    .clock(q_211_clock),
    .reset(q_211_reset),
    .io_enq_ready(q_211_io_enq_ready),
    .io_enq_valid(q_211_io_enq_valid),
    .io_enq_bits(q_211_io_enq_bits),
    .io_deq_ready(q_211_io_deq_ready),
    .io_deq_valid(q_211_io_deq_valid),
    .io_deq_bits(q_211_io_deq_bits)
  );
  Queue q_212 ( // @[Decoupled.scala 361:21]
    .clock(q_212_clock),
    .reset(q_212_reset),
    .io_enq_ready(q_212_io_enq_ready),
    .io_enq_valid(q_212_io_enq_valid),
    .io_enq_bits(q_212_io_enq_bits),
    .io_deq_ready(q_212_io_deq_ready),
    .io_deq_valid(q_212_io_deq_valid),
    .io_deq_bits(q_212_io_deq_bits)
  );
  Queue q_213 ( // @[Decoupled.scala 361:21]
    .clock(q_213_clock),
    .reset(q_213_reset),
    .io_enq_ready(q_213_io_enq_ready),
    .io_enq_valid(q_213_io_enq_valid),
    .io_enq_bits(q_213_io_enq_bits),
    .io_deq_ready(q_213_io_deq_ready),
    .io_deq_valid(q_213_io_deq_valid),
    .io_deq_bits(q_213_io_deq_bits)
  );
  Queue q_214 ( // @[Decoupled.scala 361:21]
    .clock(q_214_clock),
    .reset(q_214_reset),
    .io_enq_ready(q_214_io_enq_ready),
    .io_enq_valid(q_214_io_enq_valid),
    .io_enq_bits(q_214_io_enq_bits),
    .io_deq_ready(q_214_io_deq_ready),
    .io_deq_valid(q_214_io_deq_valid),
    .io_deq_bits(q_214_io_deq_bits)
  );
  Queue q_215 ( // @[Decoupled.scala 361:21]
    .clock(q_215_clock),
    .reset(q_215_reset),
    .io_enq_ready(q_215_io_enq_ready),
    .io_enq_valid(q_215_io_enq_valid),
    .io_enq_bits(q_215_io_enq_bits),
    .io_deq_ready(q_215_io_deq_ready),
    .io_deq_valid(q_215_io_deq_valid),
    .io_deq_bits(q_215_io_deq_bits)
  );
  Queue q_216 ( // @[Decoupled.scala 361:21]
    .clock(q_216_clock),
    .reset(q_216_reset),
    .io_enq_ready(q_216_io_enq_ready),
    .io_enq_valid(q_216_io_enq_valid),
    .io_enq_bits(q_216_io_enq_bits),
    .io_deq_ready(q_216_io_deq_ready),
    .io_deq_valid(q_216_io_deq_valid),
    .io_deq_bits(q_216_io_deq_bits)
  );
  Queue q_217 ( // @[Decoupled.scala 361:21]
    .clock(q_217_clock),
    .reset(q_217_reset),
    .io_enq_ready(q_217_io_enq_ready),
    .io_enq_valid(q_217_io_enq_valid),
    .io_enq_bits(q_217_io_enq_bits),
    .io_deq_ready(q_217_io_deq_ready),
    .io_deq_valid(q_217_io_deq_valid),
    .io_deq_bits(q_217_io_deq_bits)
  );
  Queue q_218 ( // @[Decoupled.scala 361:21]
    .clock(q_218_clock),
    .reset(q_218_reset),
    .io_enq_ready(q_218_io_enq_ready),
    .io_enq_valid(q_218_io_enq_valid),
    .io_enq_bits(q_218_io_enq_bits),
    .io_deq_ready(q_218_io_deq_ready),
    .io_deq_valid(q_218_io_deq_valid),
    .io_deq_bits(q_218_io_deq_bits)
  );
  Queue q_219 ( // @[Decoupled.scala 361:21]
    .clock(q_219_clock),
    .reset(q_219_reset),
    .io_enq_ready(q_219_io_enq_ready),
    .io_enq_valid(q_219_io_enq_valid),
    .io_enq_bits(q_219_io_enq_bits),
    .io_deq_ready(q_219_io_deq_ready),
    .io_deq_valid(q_219_io_deq_valid),
    .io_deq_bits(q_219_io_deq_bits)
  );
  Queue q_220 ( // @[Decoupled.scala 361:21]
    .clock(q_220_clock),
    .reset(q_220_reset),
    .io_enq_ready(q_220_io_enq_ready),
    .io_enq_valid(q_220_io_enq_valid),
    .io_enq_bits(q_220_io_enq_bits),
    .io_deq_ready(q_220_io_deq_ready),
    .io_deq_valid(q_220_io_deq_valid),
    .io_deq_bits(q_220_io_deq_bits)
  );
  Queue q_221 ( // @[Decoupled.scala 361:21]
    .clock(q_221_clock),
    .reset(q_221_reset),
    .io_enq_ready(q_221_io_enq_ready),
    .io_enq_valid(q_221_io_enq_valid),
    .io_enq_bits(q_221_io_enq_bits),
    .io_deq_ready(q_221_io_deq_ready),
    .io_deq_valid(q_221_io_deq_valid),
    .io_deq_bits(q_221_io_deq_bits)
  );
  Queue q_222 ( // @[Decoupled.scala 361:21]
    .clock(q_222_clock),
    .reset(q_222_reset),
    .io_enq_ready(q_222_io_enq_ready),
    .io_enq_valid(q_222_io_enq_valid),
    .io_enq_bits(q_222_io_enq_bits),
    .io_deq_ready(q_222_io_deq_ready),
    .io_deq_valid(q_222_io_deq_valid),
    .io_deq_bits(q_222_io_deq_bits)
  );
  Queue q_223 ( // @[Decoupled.scala 361:21]
    .clock(q_223_clock),
    .reset(q_223_reset),
    .io_enq_ready(q_223_io_enq_ready),
    .io_enq_valid(q_223_io_enq_valid),
    .io_enq_bits(q_223_io_enq_bits),
    .io_deq_ready(q_223_io_deq_ready),
    .io_deq_valid(q_223_io_deq_valid),
    .io_deq_bits(q_223_io_deq_bits)
  );
  Queue q_224 ( // @[Decoupled.scala 361:21]
    .clock(q_224_clock),
    .reset(q_224_reset),
    .io_enq_ready(q_224_io_enq_ready),
    .io_enq_valid(q_224_io_enq_valid),
    .io_enq_bits(q_224_io_enq_bits),
    .io_deq_ready(q_224_io_deq_ready),
    .io_deq_valid(q_224_io_deq_valid),
    .io_deq_bits(q_224_io_deq_bits)
  );
  Queue q_225 ( // @[Decoupled.scala 361:21]
    .clock(q_225_clock),
    .reset(q_225_reset),
    .io_enq_ready(q_225_io_enq_ready),
    .io_enq_valid(q_225_io_enq_valid),
    .io_enq_bits(q_225_io_enq_bits),
    .io_deq_ready(q_225_io_deq_ready),
    .io_deq_valid(q_225_io_deq_valid),
    .io_deq_bits(q_225_io_deq_bits)
  );
  Queue q_226 ( // @[Decoupled.scala 361:21]
    .clock(q_226_clock),
    .reset(q_226_reset),
    .io_enq_ready(q_226_io_enq_ready),
    .io_enq_valid(q_226_io_enq_valid),
    .io_enq_bits(q_226_io_enq_bits),
    .io_deq_ready(q_226_io_deq_ready),
    .io_deq_valid(q_226_io_deq_valid),
    .io_deq_bits(q_226_io_deq_bits)
  );
  Queue q_227 ( // @[Decoupled.scala 361:21]
    .clock(q_227_clock),
    .reset(q_227_reset),
    .io_enq_ready(q_227_io_enq_ready),
    .io_enq_valid(q_227_io_enq_valid),
    .io_enq_bits(q_227_io_enq_bits),
    .io_deq_ready(q_227_io_deq_ready),
    .io_deq_valid(q_227_io_deq_valid),
    .io_deq_bits(q_227_io_deq_bits)
  );
  Queue q_228 ( // @[Decoupled.scala 361:21]
    .clock(q_228_clock),
    .reset(q_228_reset),
    .io_enq_ready(q_228_io_enq_ready),
    .io_enq_valid(q_228_io_enq_valid),
    .io_enq_bits(q_228_io_enq_bits),
    .io_deq_ready(q_228_io_deq_ready),
    .io_deq_valid(q_228_io_deq_valid),
    .io_deq_bits(q_228_io_deq_bits)
  );
  Queue q_229 ( // @[Decoupled.scala 361:21]
    .clock(q_229_clock),
    .reset(q_229_reset),
    .io_enq_ready(q_229_io_enq_ready),
    .io_enq_valid(q_229_io_enq_valid),
    .io_enq_bits(q_229_io_enq_bits),
    .io_deq_ready(q_229_io_deq_ready),
    .io_deq_valid(q_229_io_deq_valid),
    .io_deq_bits(q_229_io_deq_bits)
  );
  Queue q_230 ( // @[Decoupled.scala 361:21]
    .clock(q_230_clock),
    .reset(q_230_reset),
    .io_enq_ready(q_230_io_enq_ready),
    .io_enq_valid(q_230_io_enq_valid),
    .io_enq_bits(q_230_io_enq_bits),
    .io_deq_ready(q_230_io_deq_ready),
    .io_deq_valid(q_230_io_deq_valid),
    .io_deq_bits(q_230_io_deq_bits)
  );
  Queue q_231 ( // @[Decoupled.scala 361:21]
    .clock(q_231_clock),
    .reset(q_231_reset),
    .io_enq_ready(q_231_io_enq_ready),
    .io_enq_valid(q_231_io_enq_valid),
    .io_enq_bits(q_231_io_enq_bits),
    .io_deq_ready(q_231_io_deq_ready),
    .io_deq_valid(q_231_io_deq_valid),
    .io_deq_bits(q_231_io_deq_bits)
  );
  Queue q_232 ( // @[Decoupled.scala 361:21]
    .clock(q_232_clock),
    .reset(q_232_reset),
    .io_enq_ready(q_232_io_enq_ready),
    .io_enq_valid(q_232_io_enq_valid),
    .io_enq_bits(q_232_io_enq_bits),
    .io_deq_ready(q_232_io_deq_ready),
    .io_deq_valid(q_232_io_deq_valid),
    .io_deq_bits(q_232_io_deq_bits)
  );
  Queue q_233 ( // @[Decoupled.scala 361:21]
    .clock(q_233_clock),
    .reset(q_233_reset),
    .io_enq_ready(q_233_io_enq_ready),
    .io_enq_valid(q_233_io_enq_valid),
    .io_enq_bits(q_233_io_enq_bits),
    .io_deq_ready(q_233_io_deq_ready),
    .io_deq_valid(q_233_io_deq_valid),
    .io_deq_bits(q_233_io_deq_bits)
  );
  Queue q_234 ( // @[Decoupled.scala 361:21]
    .clock(q_234_clock),
    .reset(q_234_reset),
    .io_enq_ready(q_234_io_enq_ready),
    .io_enq_valid(q_234_io_enq_valid),
    .io_enq_bits(q_234_io_enq_bits),
    .io_deq_ready(q_234_io_deq_ready),
    .io_deq_valid(q_234_io_deq_valid),
    .io_deq_bits(q_234_io_deq_bits)
  );
  Queue q_235 ( // @[Decoupled.scala 361:21]
    .clock(q_235_clock),
    .reset(q_235_reset),
    .io_enq_ready(q_235_io_enq_ready),
    .io_enq_valid(q_235_io_enq_valid),
    .io_enq_bits(q_235_io_enq_bits),
    .io_deq_ready(q_235_io_deq_ready),
    .io_deq_valid(q_235_io_deq_valid),
    .io_deq_bits(q_235_io_deq_bits)
  );
  Queue q_236 ( // @[Decoupled.scala 361:21]
    .clock(q_236_clock),
    .reset(q_236_reset),
    .io_enq_ready(q_236_io_enq_ready),
    .io_enq_valid(q_236_io_enq_valid),
    .io_enq_bits(q_236_io_enq_bits),
    .io_deq_ready(q_236_io_deq_ready),
    .io_deq_valid(q_236_io_deq_valid),
    .io_deq_bits(q_236_io_deq_bits)
  );
  Queue q_237 ( // @[Decoupled.scala 361:21]
    .clock(q_237_clock),
    .reset(q_237_reset),
    .io_enq_ready(q_237_io_enq_ready),
    .io_enq_valid(q_237_io_enq_valid),
    .io_enq_bits(q_237_io_enq_bits),
    .io_deq_ready(q_237_io_deq_ready),
    .io_deq_valid(q_237_io_deq_valid),
    .io_deq_bits(q_237_io_deq_bits)
  );
  Queue q_238 ( // @[Decoupled.scala 361:21]
    .clock(q_238_clock),
    .reset(q_238_reset),
    .io_enq_ready(q_238_io_enq_ready),
    .io_enq_valid(q_238_io_enq_valid),
    .io_enq_bits(q_238_io_enq_bits),
    .io_deq_ready(q_238_io_deq_ready),
    .io_deq_valid(q_238_io_deq_valid),
    .io_deq_bits(q_238_io_deq_bits)
  );
  Queue q_239 ( // @[Decoupled.scala 361:21]
    .clock(q_239_clock),
    .reset(q_239_reset),
    .io_enq_ready(q_239_io_enq_ready),
    .io_enq_valid(q_239_io_enq_valid),
    .io_enq_bits(q_239_io_enq_bits),
    .io_deq_ready(q_239_io_deq_ready),
    .io_deq_valid(q_239_io_deq_valid),
    .io_deq_bits(q_239_io_deq_bits)
  );
  Queue q_240 ( // @[Decoupled.scala 361:21]
    .clock(q_240_clock),
    .reset(q_240_reset),
    .io_enq_ready(q_240_io_enq_ready),
    .io_enq_valid(q_240_io_enq_valid),
    .io_enq_bits(q_240_io_enq_bits),
    .io_deq_ready(q_240_io_deq_ready),
    .io_deq_valid(q_240_io_deq_valid),
    .io_deq_bits(q_240_io_deq_bits)
  );
  Queue q_241 ( // @[Decoupled.scala 361:21]
    .clock(q_241_clock),
    .reset(q_241_reset),
    .io_enq_ready(q_241_io_enq_ready),
    .io_enq_valid(q_241_io_enq_valid),
    .io_enq_bits(q_241_io_enq_bits),
    .io_deq_ready(q_241_io_deq_ready),
    .io_deq_valid(q_241_io_deq_valid),
    .io_deq_bits(q_241_io_deq_bits)
  );
  Queue q_242 ( // @[Decoupled.scala 361:21]
    .clock(q_242_clock),
    .reset(q_242_reset),
    .io_enq_ready(q_242_io_enq_ready),
    .io_enq_valid(q_242_io_enq_valid),
    .io_enq_bits(q_242_io_enq_bits),
    .io_deq_ready(q_242_io_deq_ready),
    .io_deq_valid(q_242_io_deq_valid),
    .io_deq_bits(q_242_io_deq_bits)
  );
  Queue q_243 ( // @[Decoupled.scala 361:21]
    .clock(q_243_clock),
    .reset(q_243_reset),
    .io_enq_ready(q_243_io_enq_ready),
    .io_enq_valid(q_243_io_enq_valid),
    .io_enq_bits(q_243_io_enq_bits),
    .io_deq_ready(q_243_io_deq_ready),
    .io_deq_valid(q_243_io_deq_valid),
    .io_deq_bits(q_243_io_deq_bits)
  );
  Queue q_244 ( // @[Decoupled.scala 361:21]
    .clock(q_244_clock),
    .reset(q_244_reset),
    .io_enq_ready(q_244_io_enq_ready),
    .io_enq_valid(q_244_io_enq_valid),
    .io_enq_bits(q_244_io_enq_bits),
    .io_deq_ready(q_244_io_deq_ready),
    .io_deq_valid(q_244_io_deq_valid),
    .io_deq_bits(q_244_io_deq_bits)
  );
  Queue q_245 ( // @[Decoupled.scala 361:21]
    .clock(q_245_clock),
    .reset(q_245_reset),
    .io_enq_ready(q_245_io_enq_ready),
    .io_enq_valid(q_245_io_enq_valid),
    .io_enq_bits(q_245_io_enq_bits),
    .io_deq_ready(q_245_io_deq_ready),
    .io_deq_valid(q_245_io_deq_valid),
    .io_deq_bits(q_245_io_deq_bits)
  );
  Queue q_246 ( // @[Decoupled.scala 361:21]
    .clock(q_246_clock),
    .reset(q_246_reset),
    .io_enq_ready(q_246_io_enq_ready),
    .io_enq_valid(q_246_io_enq_valid),
    .io_enq_bits(q_246_io_enq_bits),
    .io_deq_ready(q_246_io_deq_ready),
    .io_deq_valid(q_246_io_deq_valid),
    .io_deq_bits(q_246_io_deq_bits)
  );
  Queue q_247 ( // @[Decoupled.scala 361:21]
    .clock(q_247_clock),
    .reset(q_247_reset),
    .io_enq_ready(q_247_io_enq_ready),
    .io_enq_valid(q_247_io_enq_valid),
    .io_enq_bits(q_247_io_enq_bits),
    .io_deq_ready(q_247_io_deq_ready),
    .io_deq_valid(q_247_io_deq_valid),
    .io_deq_bits(q_247_io_deq_bits)
  );
  Queue q_248 ( // @[Decoupled.scala 361:21]
    .clock(q_248_clock),
    .reset(q_248_reset),
    .io_enq_ready(q_248_io_enq_ready),
    .io_enq_valid(q_248_io_enq_valid),
    .io_enq_bits(q_248_io_enq_bits),
    .io_deq_ready(q_248_io_deq_ready),
    .io_deq_valid(q_248_io_deq_valid),
    .io_deq_bits(q_248_io_deq_bits)
  );
  Queue q_249 ( // @[Decoupled.scala 361:21]
    .clock(q_249_clock),
    .reset(q_249_reset),
    .io_enq_ready(q_249_io_enq_ready),
    .io_enq_valid(q_249_io_enq_valid),
    .io_enq_bits(q_249_io_enq_bits),
    .io_deq_ready(q_249_io_deq_ready),
    .io_deq_valid(q_249_io_deq_valid),
    .io_deq_bits(q_249_io_deq_bits)
  );
  Queue q_250 ( // @[Decoupled.scala 361:21]
    .clock(q_250_clock),
    .reset(q_250_reset),
    .io_enq_ready(q_250_io_enq_ready),
    .io_enq_valid(q_250_io_enq_valid),
    .io_enq_bits(q_250_io_enq_bits),
    .io_deq_ready(q_250_io_deq_ready),
    .io_deq_valid(q_250_io_deq_valid),
    .io_deq_bits(q_250_io_deq_bits)
  );
  Queue q_251 ( // @[Decoupled.scala 361:21]
    .clock(q_251_clock),
    .reset(q_251_reset),
    .io_enq_ready(q_251_io_enq_ready),
    .io_enq_valid(q_251_io_enq_valid),
    .io_enq_bits(q_251_io_enq_bits),
    .io_deq_ready(q_251_io_deq_ready),
    .io_deq_valid(q_251_io_deq_valid),
    .io_deq_bits(q_251_io_deq_bits)
  );
  Queue q_252 ( // @[Decoupled.scala 361:21]
    .clock(q_252_clock),
    .reset(q_252_reset),
    .io_enq_ready(q_252_io_enq_ready),
    .io_enq_valid(q_252_io_enq_valid),
    .io_enq_bits(q_252_io_enq_bits),
    .io_deq_ready(q_252_io_deq_ready),
    .io_deq_valid(q_252_io_deq_valid),
    .io_deq_bits(q_252_io_deq_bits)
  );
  Queue q_253 ( // @[Decoupled.scala 361:21]
    .clock(q_253_clock),
    .reset(q_253_reset),
    .io_enq_ready(q_253_io_enq_ready),
    .io_enq_valid(q_253_io_enq_valid),
    .io_enq_bits(q_253_io_enq_bits),
    .io_deq_ready(q_253_io_deq_ready),
    .io_deq_valid(q_253_io_deq_valid),
    .io_deq_bits(q_253_io_deq_bits)
  );
  Queue q_254 ( // @[Decoupled.scala 361:21]
    .clock(q_254_clock),
    .reset(q_254_reset),
    .io_enq_ready(q_254_io_enq_ready),
    .io_enq_valid(q_254_io_enq_valid),
    .io_enq_bits(q_254_io_enq_bits),
    .io_deq_ready(q_254_io_deq_ready),
    .io_deq_valid(q_254_io_deq_valid),
    .io_deq_bits(q_254_io_deq_bits)
  );
  Queue q_255 ( // @[Decoupled.scala 361:21]
    .clock(q_255_clock),
    .reset(q_255_reset),
    .io_enq_ready(q_255_io_enq_ready),
    .io_enq_valid(q_255_io_enq_valid),
    .io_enq_bits(q_255_io_enq_bits),
    .io_deq_ready(q_255_io_deq_ready),
    .io_deq_valid(q_255_io_deq_valid),
    .io_deq_bits(q_255_io_deq_bits)
  );
  Queue q_256 ( // @[Decoupled.scala 361:21]
    .clock(q_256_clock),
    .reset(q_256_reset),
    .io_enq_ready(q_256_io_enq_ready),
    .io_enq_valid(q_256_io_enq_valid),
    .io_enq_bits(q_256_io_enq_bits),
    .io_deq_ready(q_256_io_deq_ready),
    .io_deq_valid(q_256_io_deq_valid),
    .io_deq_bits(q_256_io_deq_bits)
  );
  Queue q_257 ( // @[Decoupled.scala 361:21]
    .clock(q_257_clock),
    .reset(q_257_reset),
    .io_enq_ready(q_257_io_enq_ready),
    .io_enq_valid(q_257_io_enq_valid),
    .io_enq_bits(q_257_io_enq_bits),
    .io_deq_ready(q_257_io_deq_ready),
    .io_deq_valid(q_257_io_deq_valid),
    .io_deq_bits(q_257_io_deq_bits)
  );
  Queue q_258 ( // @[Decoupled.scala 361:21]
    .clock(q_258_clock),
    .reset(q_258_reset),
    .io_enq_ready(q_258_io_enq_ready),
    .io_enq_valid(q_258_io_enq_valid),
    .io_enq_bits(q_258_io_enq_bits),
    .io_deq_ready(q_258_io_deq_ready),
    .io_deq_valid(q_258_io_deq_valid),
    .io_deq_bits(q_258_io_deq_bits)
  );
  Queue q_259 ( // @[Decoupled.scala 361:21]
    .clock(q_259_clock),
    .reset(q_259_reset),
    .io_enq_ready(q_259_io_enq_ready),
    .io_enq_valid(q_259_io_enq_valid),
    .io_enq_bits(q_259_io_enq_bits),
    .io_deq_ready(q_259_io_deq_ready),
    .io_deq_valid(q_259_io_deq_valid),
    .io_deq_bits(q_259_io_deq_bits)
  );
  Queue q_260 ( // @[Decoupled.scala 361:21]
    .clock(q_260_clock),
    .reset(q_260_reset),
    .io_enq_ready(q_260_io_enq_ready),
    .io_enq_valid(q_260_io_enq_valid),
    .io_enq_bits(q_260_io_enq_bits),
    .io_deq_ready(q_260_io_deq_ready),
    .io_deq_valid(q_260_io_deq_valid),
    .io_deq_bits(q_260_io_deq_bits)
  );
  Queue q_261 ( // @[Decoupled.scala 361:21]
    .clock(q_261_clock),
    .reset(q_261_reset),
    .io_enq_ready(q_261_io_enq_ready),
    .io_enq_valid(q_261_io_enq_valid),
    .io_enq_bits(q_261_io_enq_bits),
    .io_deq_ready(q_261_io_deq_ready),
    .io_deq_valid(q_261_io_deq_valid),
    .io_deq_bits(q_261_io_deq_bits)
  );
  Queue q_262 ( // @[Decoupled.scala 361:21]
    .clock(q_262_clock),
    .reset(q_262_reset),
    .io_enq_ready(q_262_io_enq_ready),
    .io_enq_valid(q_262_io_enq_valid),
    .io_enq_bits(q_262_io_enq_bits),
    .io_deq_ready(q_262_io_deq_ready),
    .io_deq_valid(q_262_io_deq_valid),
    .io_deq_bits(q_262_io_deq_bits)
  );
  Queue q_263 ( // @[Decoupled.scala 361:21]
    .clock(q_263_clock),
    .reset(q_263_reset),
    .io_enq_ready(q_263_io_enq_ready),
    .io_enq_valid(q_263_io_enq_valid),
    .io_enq_bits(q_263_io_enq_bits),
    .io_deq_ready(q_263_io_deq_ready),
    .io_deq_valid(q_263_io_deq_valid),
    .io_deq_bits(q_263_io_deq_bits)
  );
  Queue q_264 ( // @[Decoupled.scala 361:21]
    .clock(q_264_clock),
    .reset(q_264_reset),
    .io_enq_ready(q_264_io_enq_ready),
    .io_enq_valid(q_264_io_enq_valid),
    .io_enq_bits(q_264_io_enq_bits),
    .io_deq_ready(q_264_io_deq_ready),
    .io_deq_valid(q_264_io_deq_valid),
    .io_deq_bits(q_264_io_deq_bits)
  );
  Queue q_265 ( // @[Decoupled.scala 361:21]
    .clock(q_265_clock),
    .reset(q_265_reset),
    .io_enq_ready(q_265_io_enq_ready),
    .io_enq_valid(q_265_io_enq_valid),
    .io_enq_bits(q_265_io_enq_bits),
    .io_deq_ready(q_265_io_deq_ready),
    .io_deq_valid(q_265_io_deq_valid),
    .io_deq_bits(q_265_io_deq_bits)
  );
  Queue q_266 ( // @[Decoupled.scala 361:21]
    .clock(q_266_clock),
    .reset(q_266_reset),
    .io_enq_ready(q_266_io_enq_ready),
    .io_enq_valid(q_266_io_enq_valid),
    .io_enq_bits(q_266_io_enq_bits),
    .io_deq_ready(q_266_io_deq_ready),
    .io_deq_valid(q_266_io_deq_valid),
    .io_deq_bits(q_266_io_deq_bits)
  );
  Queue q_267 ( // @[Decoupled.scala 361:21]
    .clock(q_267_clock),
    .reset(q_267_reset),
    .io_enq_ready(q_267_io_enq_ready),
    .io_enq_valid(q_267_io_enq_valid),
    .io_enq_bits(q_267_io_enq_bits),
    .io_deq_ready(q_267_io_deq_ready),
    .io_deq_valid(q_267_io_deq_valid),
    .io_deq_bits(q_267_io_deq_bits)
  );
  Queue q_268 ( // @[Decoupled.scala 361:21]
    .clock(q_268_clock),
    .reset(q_268_reset),
    .io_enq_ready(q_268_io_enq_ready),
    .io_enq_valid(q_268_io_enq_valid),
    .io_enq_bits(q_268_io_enq_bits),
    .io_deq_ready(q_268_io_deq_ready),
    .io_deq_valid(q_268_io_deq_valid),
    .io_deq_bits(q_268_io_deq_bits)
  );
  Queue q_269 ( // @[Decoupled.scala 361:21]
    .clock(q_269_clock),
    .reset(q_269_reset),
    .io_enq_ready(q_269_io_enq_ready),
    .io_enq_valid(q_269_io_enq_valid),
    .io_enq_bits(q_269_io_enq_bits),
    .io_deq_ready(q_269_io_deq_ready),
    .io_deq_valid(q_269_io_deq_valid),
    .io_deq_bits(q_269_io_deq_bits)
  );
  Queue q_270 ( // @[Decoupled.scala 361:21]
    .clock(q_270_clock),
    .reset(q_270_reset),
    .io_enq_ready(q_270_io_enq_ready),
    .io_enq_valid(q_270_io_enq_valid),
    .io_enq_bits(q_270_io_enq_bits),
    .io_deq_ready(q_270_io_deq_ready),
    .io_deq_valid(q_270_io_deq_valid),
    .io_deq_bits(q_270_io_deq_bits)
  );
  Queue q_271 ( // @[Decoupled.scala 361:21]
    .clock(q_271_clock),
    .reset(q_271_reset),
    .io_enq_ready(q_271_io_enq_ready),
    .io_enq_valid(q_271_io_enq_valid),
    .io_enq_bits(q_271_io_enq_bits),
    .io_deq_ready(q_271_io_deq_ready),
    .io_deq_valid(q_271_io_deq_valid),
    .io_deq_bits(q_271_io_deq_bits)
  );
  Queue q_272 ( // @[Decoupled.scala 361:21]
    .clock(q_272_clock),
    .reset(q_272_reset),
    .io_enq_ready(q_272_io_enq_ready),
    .io_enq_valid(q_272_io_enq_valid),
    .io_enq_bits(q_272_io_enq_bits),
    .io_deq_ready(q_272_io_deq_ready),
    .io_deq_valid(q_272_io_deq_valid),
    .io_deq_bits(q_272_io_deq_bits)
  );
  Queue q_273 ( // @[Decoupled.scala 361:21]
    .clock(q_273_clock),
    .reset(q_273_reset),
    .io_enq_ready(q_273_io_enq_ready),
    .io_enq_valid(q_273_io_enq_valid),
    .io_enq_bits(q_273_io_enq_bits),
    .io_deq_ready(q_273_io_deq_ready),
    .io_deq_valid(q_273_io_deq_valid),
    .io_deq_bits(q_273_io_deq_bits)
  );
  Queue q_274 ( // @[Decoupled.scala 361:21]
    .clock(q_274_clock),
    .reset(q_274_reset),
    .io_enq_ready(q_274_io_enq_ready),
    .io_enq_valid(q_274_io_enq_valid),
    .io_enq_bits(q_274_io_enq_bits),
    .io_deq_ready(q_274_io_deq_ready),
    .io_deq_valid(q_274_io_deq_valid),
    .io_deq_bits(q_274_io_deq_bits)
  );
  Queue q_275 ( // @[Decoupled.scala 361:21]
    .clock(q_275_clock),
    .reset(q_275_reset),
    .io_enq_ready(q_275_io_enq_ready),
    .io_enq_valid(q_275_io_enq_valid),
    .io_enq_bits(q_275_io_enq_bits),
    .io_deq_ready(q_275_io_deq_ready),
    .io_deq_valid(q_275_io_deq_valid),
    .io_deq_bits(q_275_io_deq_bits)
  );
  Queue q_276 ( // @[Decoupled.scala 361:21]
    .clock(q_276_clock),
    .reset(q_276_reset),
    .io_enq_ready(q_276_io_enq_ready),
    .io_enq_valid(q_276_io_enq_valid),
    .io_enq_bits(q_276_io_enq_bits),
    .io_deq_ready(q_276_io_deq_ready),
    .io_deq_valid(q_276_io_deq_valid),
    .io_deq_bits(q_276_io_deq_bits)
  );
  Queue q_277 ( // @[Decoupled.scala 361:21]
    .clock(q_277_clock),
    .reset(q_277_reset),
    .io_enq_ready(q_277_io_enq_ready),
    .io_enq_valid(q_277_io_enq_valid),
    .io_enq_bits(q_277_io_enq_bits),
    .io_deq_ready(q_277_io_deq_ready),
    .io_deq_valid(q_277_io_deq_valid),
    .io_deq_bits(q_277_io_deq_bits)
  );
  Queue q_278 ( // @[Decoupled.scala 361:21]
    .clock(q_278_clock),
    .reset(q_278_reset),
    .io_enq_ready(q_278_io_enq_ready),
    .io_enq_valid(q_278_io_enq_valid),
    .io_enq_bits(q_278_io_enq_bits),
    .io_deq_ready(q_278_io_deq_ready),
    .io_deq_valid(q_278_io_deq_valid),
    .io_deq_bits(q_278_io_deq_bits)
  );
  Queue q_279 ( // @[Decoupled.scala 361:21]
    .clock(q_279_clock),
    .reset(q_279_reset),
    .io_enq_ready(q_279_io_enq_ready),
    .io_enq_valid(q_279_io_enq_valid),
    .io_enq_bits(q_279_io_enq_bits),
    .io_deq_ready(q_279_io_deq_ready),
    .io_deq_valid(q_279_io_deq_valid),
    .io_deq_bits(q_279_io_deq_bits)
  );
  Queue q_280 ( // @[Decoupled.scala 361:21]
    .clock(q_280_clock),
    .reset(q_280_reset),
    .io_enq_ready(q_280_io_enq_ready),
    .io_enq_valid(q_280_io_enq_valid),
    .io_enq_bits(q_280_io_enq_bits),
    .io_deq_ready(q_280_io_deq_ready),
    .io_deq_valid(q_280_io_deq_valid),
    .io_deq_bits(q_280_io_deq_bits)
  );
  Queue q_281 ( // @[Decoupled.scala 361:21]
    .clock(q_281_clock),
    .reset(q_281_reset),
    .io_enq_ready(q_281_io_enq_ready),
    .io_enq_valid(q_281_io_enq_valid),
    .io_enq_bits(q_281_io_enq_bits),
    .io_deq_ready(q_281_io_deq_ready),
    .io_deq_valid(q_281_io_deq_valid),
    .io_deq_bits(q_281_io_deq_bits)
  );
  Queue q_282 ( // @[Decoupled.scala 361:21]
    .clock(q_282_clock),
    .reset(q_282_reset),
    .io_enq_ready(q_282_io_enq_ready),
    .io_enq_valid(q_282_io_enq_valid),
    .io_enq_bits(q_282_io_enq_bits),
    .io_deq_ready(q_282_io_deq_ready),
    .io_deq_valid(q_282_io_deq_valid),
    .io_deq_bits(q_282_io_deq_bits)
  );
  Queue q_283 ( // @[Decoupled.scala 361:21]
    .clock(q_283_clock),
    .reset(q_283_reset),
    .io_enq_ready(q_283_io_enq_ready),
    .io_enq_valid(q_283_io_enq_valid),
    .io_enq_bits(q_283_io_enq_bits),
    .io_deq_ready(q_283_io_deq_ready),
    .io_deq_valid(q_283_io_deq_valid),
    .io_deq_bits(q_283_io_deq_bits)
  );
  Queue q_284 ( // @[Decoupled.scala 361:21]
    .clock(q_284_clock),
    .reset(q_284_reset),
    .io_enq_ready(q_284_io_enq_ready),
    .io_enq_valid(q_284_io_enq_valid),
    .io_enq_bits(q_284_io_enq_bits),
    .io_deq_ready(q_284_io_deq_ready),
    .io_deq_valid(q_284_io_deq_valid),
    .io_deq_bits(q_284_io_deq_bits)
  );
  Queue q_285 ( // @[Decoupled.scala 361:21]
    .clock(q_285_clock),
    .reset(q_285_reset),
    .io_enq_ready(q_285_io_enq_ready),
    .io_enq_valid(q_285_io_enq_valid),
    .io_enq_bits(q_285_io_enq_bits),
    .io_deq_ready(q_285_io_deq_ready),
    .io_deq_valid(q_285_io_deq_valid),
    .io_deq_bits(q_285_io_deq_bits)
  );
  Queue q_286 ( // @[Decoupled.scala 361:21]
    .clock(q_286_clock),
    .reset(q_286_reset),
    .io_enq_ready(q_286_io_enq_ready),
    .io_enq_valid(q_286_io_enq_valid),
    .io_enq_bits(q_286_io_enq_bits),
    .io_deq_ready(q_286_io_deq_ready),
    .io_deq_valid(q_286_io_deq_valid),
    .io_deq_bits(q_286_io_deq_bits)
  );
  Queue q_287 ( // @[Decoupled.scala 361:21]
    .clock(q_287_clock),
    .reset(q_287_reset),
    .io_enq_ready(q_287_io_enq_ready),
    .io_enq_valid(q_287_io_enq_valid),
    .io_enq_bits(q_287_io_enq_bits),
    .io_deq_ready(q_287_io_deq_ready),
    .io_deq_valid(q_287_io_deq_valid),
    .io_deq_bits(q_287_io_deq_bits)
  );
  Queue q_288 ( // @[Decoupled.scala 361:21]
    .clock(q_288_clock),
    .reset(q_288_reset),
    .io_enq_ready(q_288_io_enq_ready),
    .io_enq_valid(q_288_io_enq_valid),
    .io_enq_bits(q_288_io_enq_bits),
    .io_deq_ready(q_288_io_deq_ready),
    .io_deq_valid(q_288_io_deq_valid),
    .io_deq_bits(q_288_io_deq_bits)
  );
  Queue q_289 ( // @[Decoupled.scala 361:21]
    .clock(q_289_clock),
    .reset(q_289_reset),
    .io_enq_ready(q_289_io_enq_ready),
    .io_enq_valid(q_289_io_enq_valid),
    .io_enq_bits(q_289_io_enq_bits),
    .io_deq_ready(q_289_io_deq_ready),
    .io_deq_valid(q_289_io_deq_valid),
    .io_deq_bits(q_289_io_deq_bits)
  );
  Queue q_290 ( // @[Decoupled.scala 361:21]
    .clock(q_290_clock),
    .reset(q_290_reset),
    .io_enq_ready(q_290_io_enq_ready),
    .io_enq_valid(q_290_io_enq_valid),
    .io_enq_bits(q_290_io_enq_bits),
    .io_deq_ready(q_290_io_deq_ready),
    .io_deq_valid(q_290_io_deq_valid),
    .io_deq_bits(q_290_io_deq_bits)
  );
  Queue q_291 ( // @[Decoupled.scala 361:21]
    .clock(q_291_clock),
    .reset(q_291_reset),
    .io_enq_ready(q_291_io_enq_ready),
    .io_enq_valid(q_291_io_enq_valid),
    .io_enq_bits(q_291_io_enq_bits),
    .io_deq_ready(q_291_io_deq_ready),
    .io_deq_valid(q_291_io_deq_valid),
    .io_deq_bits(q_291_io_deq_bits)
  );
  Queue q_292 ( // @[Decoupled.scala 361:21]
    .clock(q_292_clock),
    .reset(q_292_reset),
    .io_enq_ready(q_292_io_enq_ready),
    .io_enq_valid(q_292_io_enq_valid),
    .io_enq_bits(q_292_io_enq_bits),
    .io_deq_ready(q_292_io_deq_ready),
    .io_deq_valid(q_292_io_deq_valid),
    .io_deq_bits(q_292_io_deq_bits)
  );
  Queue q_293 ( // @[Decoupled.scala 361:21]
    .clock(q_293_clock),
    .reset(q_293_reset),
    .io_enq_ready(q_293_io_enq_ready),
    .io_enq_valid(q_293_io_enq_valid),
    .io_enq_bits(q_293_io_enq_bits),
    .io_deq_ready(q_293_io_deq_ready),
    .io_deq_valid(q_293_io_deq_valid),
    .io_deq_bits(q_293_io_deq_bits)
  );
  Queue q_294 ( // @[Decoupled.scala 361:21]
    .clock(q_294_clock),
    .reset(q_294_reset),
    .io_enq_ready(q_294_io_enq_ready),
    .io_enq_valid(q_294_io_enq_valid),
    .io_enq_bits(q_294_io_enq_bits),
    .io_deq_ready(q_294_io_deq_ready),
    .io_deq_valid(q_294_io_deq_valid),
    .io_deq_bits(q_294_io_deq_bits)
  );
  Queue q_295 ( // @[Decoupled.scala 361:21]
    .clock(q_295_clock),
    .reset(q_295_reset),
    .io_enq_ready(q_295_io_enq_ready),
    .io_enq_valid(q_295_io_enq_valid),
    .io_enq_bits(q_295_io_enq_bits),
    .io_deq_ready(q_295_io_deq_ready),
    .io_deq_valid(q_295_io_deq_valid),
    .io_deq_bits(q_295_io_deq_bits)
  );
  Queue q_296 ( // @[Decoupled.scala 361:21]
    .clock(q_296_clock),
    .reset(q_296_reset),
    .io_enq_ready(q_296_io_enq_ready),
    .io_enq_valid(q_296_io_enq_valid),
    .io_enq_bits(q_296_io_enq_bits),
    .io_deq_ready(q_296_io_deq_ready),
    .io_deq_valid(q_296_io_deq_valid),
    .io_deq_bits(q_296_io_deq_bits)
  );
  Queue q_297 ( // @[Decoupled.scala 361:21]
    .clock(q_297_clock),
    .reset(q_297_reset),
    .io_enq_ready(q_297_io_enq_ready),
    .io_enq_valid(q_297_io_enq_valid),
    .io_enq_bits(q_297_io_enq_bits),
    .io_deq_ready(q_297_io_deq_ready),
    .io_deq_valid(q_297_io_deq_valid),
    .io_deq_bits(q_297_io_deq_bits)
  );
  Queue q_298 ( // @[Decoupled.scala 361:21]
    .clock(q_298_clock),
    .reset(q_298_reset),
    .io_enq_ready(q_298_io_enq_ready),
    .io_enq_valid(q_298_io_enq_valid),
    .io_enq_bits(q_298_io_enq_bits),
    .io_deq_ready(q_298_io_deq_ready),
    .io_deq_valid(q_298_io_deq_valid),
    .io_deq_bits(q_298_io_deq_bits)
  );
  Queue q_299 ( // @[Decoupled.scala 361:21]
    .clock(q_299_clock),
    .reset(q_299_reset),
    .io_enq_ready(q_299_io_enq_ready),
    .io_enq_valid(q_299_io_enq_valid),
    .io_enq_bits(q_299_io_enq_bits),
    .io_deq_ready(q_299_io_deq_ready),
    .io_deq_valid(q_299_io_deq_valid),
    .io_deq_bits(q_299_io_deq_bits)
  );
  Queue q_300 ( // @[Decoupled.scala 361:21]
    .clock(q_300_clock),
    .reset(q_300_reset),
    .io_enq_ready(q_300_io_enq_ready),
    .io_enq_valid(q_300_io_enq_valid),
    .io_enq_bits(q_300_io_enq_bits),
    .io_deq_ready(q_300_io_deq_ready),
    .io_deq_valid(q_300_io_deq_valid),
    .io_deq_bits(q_300_io_deq_bits)
  );
  Queue q_301 ( // @[Decoupled.scala 361:21]
    .clock(q_301_clock),
    .reset(q_301_reset),
    .io_enq_ready(q_301_io_enq_ready),
    .io_enq_valid(q_301_io_enq_valid),
    .io_enq_bits(q_301_io_enq_bits),
    .io_deq_ready(q_301_io_deq_ready),
    .io_deq_valid(q_301_io_deq_valid),
    .io_deq_bits(q_301_io_deq_bits)
  );
  Queue q_302 ( // @[Decoupled.scala 361:21]
    .clock(q_302_clock),
    .reset(q_302_reset),
    .io_enq_ready(q_302_io_enq_ready),
    .io_enq_valid(q_302_io_enq_valid),
    .io_enq_bits(q_302_io_enq_bits),
    .io_deq_ready(q_302_io_deq_ready),
    .io_deq_valid(q_302_io_deq_valid),
    .io_deq_bits(q_302_io_deq_bits)
  );
  Queue q_303 ( // @[Decoupled.scala 361:21]
    .clock(q_303_clock),
    .reset(q_303_reset),
    .io_enq_ready(q_303_io_enq_ready),
    .io_enq_valid(q_303_io_enq_valid),
    .io_enq_bits(q_303_io_enq_bits),
    .io_deq_ready(q_303_io_deq_ready),
    .io_deq_valid(q_303_io_deq_valid),
    .io_deq_bits(q_303_io_deq_bits)
  );
  Queue q_304 ( // @[Decoupled.scala 361:21]
    .clock(q_304_clock),
    .reset(q_304_reset),
    .io_enq_ready(q_304_io_enq_ready),
    .io_enq_valid(q_304_io_enq_valid),
    .io_enq_bits(q_304_io_enq_bits),
    .io_deq_ready(q_304_io_deq_ready),
    .io_deq_valid(q_304_io_deq_valid),
    .io_deq_bits(q_304_io_deq_bits)
  );
  Queue q_305 ( // @[Decoupled.scala 361:21]
    .clock(q_305_clock),
    .reset(q_305_reset),
    .io_enq_ready(q_305_io_enq_ready),
    .io_enq_valid(q_305_io_enq_valid),
    .io_enq_bits(q_305_io_enq_bits),
    .io_deq_ready(q_305_io_deq_ready),
    .io_deq_valid(q_305_io_deq_valid),
    .io_deq_bits(q_305_io_deq_bits)
  );
  Queue q_306 ( // @[Decoupled.scala 361:21]
    .clock(q_306_clock),
    .reset(q_306_reset),
    .io_enq_ready(q_306_io_enq_ready),
    .io_enq_valid(q_306_io_enq_valid),
    .io_enq_bits(q_306_io_enq_bits),
    .io_deq_ready(q_306_io_deq_ready),
    .io_deq_valid(q_306_io_deq_valid),
    .io_deq_bits(q_306_io_deq_bits)
  );
  Queue q_307 ( // @[Decoupled.scala 361:21]
    .clock(q_307_clock),
    .reset(q_307_reset),
    .io_enq_ready(q_307_io_enq_ready),
    .io_enq_valid(q_307_io_enq_valid),
    .io_enq_bits(q_307_io_enq_bits),
    .io_deq_ready(q_307_io_deq_ready),
    .io_deq_valid(q_307_io_deq_valid),
    .io_deq_bits(q_307_io_deq_bits)
  );
  Queue q_308 ( // @[Decoupled.scala 361:21]
    .clock(q_308_clock),
    .reset(q_308_reset),
    .io_enq_ready(q_308_io_enq_ready),
    .io_enq_valid(q_308_io_enq_valid),
    .io_enq_bits(q_308_io_enq_bits),
    .io_deq_ready(q_308_io_deq_ready),
    .io_deq_valid(q_308_io_deq_valid),
    .io_deq_bits(q_308_io_deq_bits)
  );
  Queue q_309 ( // @[Decoupled.scala 361:21]
    .clock(q_309_clock),
    .reset(q_309_reset),
    .io_enq_ready(q_309_io_enq_ready),
    .io_enq_valid(q_309_io_enq_valid),
    .io_enq_bits(q_309_io_enq_bits),
    .io_deq_ready(q_309_io_deq_ready),
    .io_deq_valid(q_309_io_deq_valid),
    .io_deq_bits(q_309_io_deq_bits)
  );
  Queue q_310 ( // @[Decoupled.scala 361:21]
    .clock(q_310_clock),
    .reset(q_310_reset),
    .io_enq_ready(q_310_io_enq_ready),
    .io_enq_valid(q_310_io_enq_valid),
    .io_enq_bits(q_310_io_enq_bits),
    .io_deq_ready(q_310_io_deq_ready),
    .io_deq_valid(q_310_io_deq_valid),
    .io_deq_bits(q_310_io_deq_bits)
  );
  Queue q_311 ( // @[Decoupled.scala 361:21]
    .clock(q_311_clock),
    .reset(q_311_reset),
    .io_enq_ready(q_311_io_enq_ready),
    .io_enq_valid(q_311_io_enq_valid),
    .io_enq_bits(q_311_io_enq_bits),
    .io_deq_ready(q_311_io_deq_ready),
    .io_deq_valid(q_311_io_deq_valid),
    .io_deq_bits(q_311_io_deq_bits)
  );
  Queue q_312 ( // @[Decoupled.scala 361:21]
    .clock(q_312_clock),
    .reset(q_312_reset),
    .io_enq_ready(q_312_io_enq_ready),
    .io_enq_valid(q_312_io_enq_valid),
    .io_enq_bits(q_312_io_enq_bits),
    .io_deq_ready(q_312_io_deq_ready),
    .io_deq_valid(q_312_io_deq_valid),
    .io_deq_bits(q_312_io_deq_bits)
  );
  Queue q_313 ( // @[Decoupled.scala 361:21]
    .clock(q_313_clock),
    .reset(q_313_reset),
    .io_enq_ready(q_313_io_enq_ready),
    .io_enq_valid(q_313_io_enq_valid),
    .io_enq_bits(q_313_io_enq_bits),
    .io_deq_ready(q_313_io_deq_ready),
    .io_deq_valid(q_313_io_deq_valid),
    .io_deq_bits(q_313_io_deq_bits)
  );
  Queue q_314 ( // @[Decoupled.scala 361:21]
    .clock(q_314_clock),
    .reset(q_314_reset),
    .io_enq_ready(q_314_io_enq_ready),
    .io_enq_valid(q_314_io_enq_valid),
    .io_enq_bits(q_314_io_enq_bits),
    .io_deq_ready(q_314_io_deq_ready),
    .io_deq_valid(q_314_io_deq_valid),
    .io_deq_bits(q_314_io_deq_bits)
  );
  Queue q_315 ( // @[Decoupled.scala 361:21]
    .clock(q_315_clock),
    .reset(q_315_reset),
    .io_enq_ready(q_315_io_enq_ready),
    .io_enq_valid(q_315_io_enq_valid),
    .io_enq_bits(q_315_io_enq_bits),
    .io_deq_ready(q_315_io_deq_ready),
    .io_deq_valid(q_315_io_deq_valid),
    .io_deq_bits(q_315_io_deq_bits)
  );
  Queue q_316 ( // @[Decoupled.scala 361:21]
    .clock(q_316_clock),
    .reset(q_316_reset),
    .io_enq_ready(q_316_io_enq_ready),
    .io_enq_valid(q_316_io_enq_valid),
    .io_enq_bits(q_316_io_enq_bits),
    .io_deq_ready(q_316_io_deq_ready),
    .io_deq_valid(q_316_io_deq_valid),
    .io_deq_bits(q_316_io_deq_bits)
  );
  Queue q_317 ( // @[Decoupled.scala 361:21]
    .clock(q_317_clock),
    .reset(q_317_reset),
    .io_enq_ready(q_317_io_enq_ready),
    .io_enq_valid(q_317_io_enq_valid),
    .io_enq_bits(q_317_io_enq_bits),
    .io_deq_ready(q_317_io_deq_ready),
    .io_deq_valid(q_317_io_deq_valid),
    .io_deq_bits(q_317_io_deq_bits)
  );
  Queue q_318 ( // @[Decoupled.scala 361:21]
    .clock(q_318_clock),
    .reset(q_318_reset),
    .io_enq_ready(q_318_io_enq_ready),
    .io_enq_valid(q_318_io_enq_valid),
    .io_enq_bits(q_318_io_enq_bits),
    .io_deq_ready(q_318_io_deq_ready),
    .io_deq_valid(q_318_io_deq_valid),
    .io_deq_bits(q_318_io_deq_bits)
  );
  Queue q_319 ( // @[Decoupled.scala 361:21]
    .clock(q_319_clock),
    .reset(q_319_reset),
    .io_enq_ready(q_319_io_enq_ready),
    .io_enq_valid(q_319_io_enq_valid),
    .io_enq_bits(q_319_io_enq_bits),
    .io_deq_ready(q_319_io_deq_ready),
    .io_deq_valid(q_319_io_deq_valid),
    .io_deq_bits(q_319_io_deq_bits)
  );
  Queue q_320 ( // @[Decoupled.scala 361:21]
    .clock(q_320_clock),
    .reset(q_320_reset),
    .io_enq_ready(q_320_io_enq_ready),
    .io_enq_valid(q_320_io_enq_valid),
    .io_enq_bits(q_320_io_enq_bits),
    .io_deq_ready(q_320_io_deq_ready),
    .io_deq_valid(q_320_io_deq_valid),
    .io_deq_bits(q_320_io_deq_bits)
  );
  Queue q_321 ( // @[Decoupled.scala 361:21]
    .clock(q_321_clock),
    .reset(q_321_reset),
    .io_enq_ready(q_321_io_enq_ready),
    .io_enq_valid(q_321_io_enq_valid),
    .io_enq_bits(q_321_io_enq_bits),
    .io_deq_ready(q_321_io_deq_ready),
    .io_deq_valid(q_321_io_deq_valid),
    .io_deq_bits(q_321_io_deq_bits)
  );
  Queue q_322 ( // @[Decoupled.scala 361:21]
    .clock(q_322_clock),
    .reset(q_322_reset),
    .io_enq_ready(q_322_io_enq_ready),
    .io_enq_valid(q_322_io_enq_valid),
    .io_enq_bits(q_322_io_enq_bits),
    .io_deq_ready(q_322_io_deq_ready),
    .io_deq_valid(q_322_io_deq_valid),
    .io_deq_bits(q_322_io_deq_bits)
  );
  Queue q_323 ( // @[Decoupled.scala 361:21]
    .clock(q_323_clock),
    .reset(q_323_reset),
    .io_enq_ready(q_323_io_enq_ready),
    .io_enq_valid(q_323_io_enq_valid),
    .io_enq_bits(q_323_io_enq_bits),
    .io_deq_ready(q_323_io_deq_ready),
    .io_deq_valid(q_323_io_deq_valid),
    .io_deq_bits(q_323_io_deq_bits)
  );
  Queue q_324 ( // @[Decoupled.scala 361:21]
    .clock(q_324_clock),
    .reset(q_324_reset),
    .io_enq_ready(q_324_io_enq_ready),
    .io_enq_valid(q_324_io_enq_valid),
    .io_enq_bits(q_324_io_enq_bits),
    .io_deq_ready(q_324_io_deq_ready),
    .io_deq_valid(q_324_io_deq_valid),
    .io_deq_bits(q_324_io_deq_bits)
  );
  Queue q_325 ( // @[Decoupled.scala 361:21]
    .clock(q_325_clock),
    .reset(q_325_reset),
    .io_enq_ready(q_325_io_enq_ready),
    .io_enq_valid(q_325_io_enq_valid),
    .io_enq_bits(q_325_io_enq_bits),
    .io_deq_ready(q_325_io_deq_ready),
    .io_deq_valid(q_325_io_deq_valid),
    .io_deq_bits(q_325_io_deq_bits)
  );
  Queue q_326 ( // @[Decoupled.scala 361:21]
    .clock(q_326_clock),
    .reset(q_326_reset),
    .io_enq_ready(q_326_io_enq_ready),
    .io_enq_valid(q_326_io_enq_valid),
    .io_enq_bits(q_326_io_enq_bits),
    .io_deq_ready(q_326_io_deq_ready),
    .io_deq_valid(q_326_io_deq_valid),
    .io_deq_bits(q_326_io_deq_bits)
  );
  Queue q_327 ( // @[Decoupled.scala 361:21]
    .clock(q_327_clock),
    .reset(q_327_reset),
    .io_enq_ready(q_327_io_enq_ready),
    .io_enq_valid(q_327_io_enq_valid),
    .io_enq_bits(q_327_io_enq_bits),
    .io_deq_ready(q_327_io_deq_ready),
    .io_deq_valid(q_327_io_deq_valid),
    .io_deq_bits(q_327_io_deq_bits)
  );
  Queue q_328 ( // @[Decoupled.scala 361:21]
    .clock(q_328_clock),
    .reset(q_328_reset),
    .io_enq_ready(q_328_io_enq_ready),
    .io_enq_valid(q_328_io_enq_valid),
    .io_enq_bits(q_328_io_enq_bits),
    .io_deq_ready(q_328_io_deq_ready),
    .io_deq_valid(q_328_io_deq_valid),
    .io_deq_bits(q_328_io_deq_bits)
  );
  Queue q_329 ( // @[Decoupled.scala 361:21]
    .clock(q_329_clock),
    .reset(q_329_reset),
    .io_enq_ready(q_329_io_enq_ready),
    .io_enq_valid(q_329_io_enq_valid),
    .io_enq_bits(q_329_io_enq_bits),
    .io_deq_ready(q_329_io_deq_ready),
    .io_deq_valid(q_329_io_deq_valid),
    .io_deq_bits(q_329_io_deq_bits)
  );
  Queue q_330 ( // @[Decoupled.scala 361:21]
    .clock(q_330_clock),
    .reset(q_330_reset),
    .io_enq_ready(q_330_io_enq_ready),
    .io_enq_valid(q_330_io_enq_valid),
    .io_enq_bits(q_330_io_enq_bits),
    .io_deq_ready(q_330_io_deq_ready),
    .io_deq_valid(q_330_io_deq_valid),
    .io_deq_bits(q_330_io_deq_bits)
  );
  Queue q_331 ( // @[Decoupled.scala 361:21]
    .clock(q_331_clock),
    .reset(q_331_reset),
    .io_enq_ready(q_331_io_enq_ready),
    .io_enq_valid(q_331_io_enq_valid),
    .io_enq_bits(q_331_io_enq_bits),
    .io_deq_ready(q_331_io_deq_ready),
    .io_deq_valid(q_331_io_deq_valid),
    .io_deq_bits(q_331_io_deq_bits)
  );
  Queue q_332 ( // @[Decoupled.scala 361:21]
    .clock(q_332_clock),
    .reset(q_332_reset),
    .io_enq_ready(q_332_io_enq_ready),
    .io_enq_valid(q_332_io_enq_valid),
    .io_enq_bits(q_332_io_enq_bits),
    .io_deq_ready(q_332_io_deq_ready),
    .io_deq_valid(q_332_io_deq_valid),
    .io_deq_bits(q_332_io_deq_bits)
  );
  Queue q_333 ( // @[Decoupled.scala 361:21]
    .clock(q_333_clock),
    .reset(q_333_reset),
    .io_enq_ready(q_333_io_enq_ready),
    .io_enq_valid(q_333_io_enq_valid),
    .io_enq_bits(q_333_io_enq_bits),
    .io_deq_ready(q_333_io_deq_ready),
    .io_deq_valid(q_333_io_deq_valid),
    .io_deq_bits(q_333_io_deq_bits)
  );
  Queue q_334 ( // @[Decoupled.scala 361:21]
    .clock(q_334_clock),
    .reset(q_334_reset),
    .io_enq_ready(q_334_io_enq_ready),
    .io_enq_valid(q_334_io_enq_valid),
    .io_enq_bits(q_334_io_enq_bits),
    .io_deq_ready(q_334_io_deq_ready),
    .io_deq_valid(q_334_io_deq_valid),
    .io_deq_bits(q_334_io_deq_bits)
  );
  Queue q_335 ( // @[Decoupled.scala 361:21]
    .clock(q_335_clock),
    .reset(q_335_reset),
    .io_enq_ready(q_335_io_enq_ready),
    .io_enq_valid(q_335_io_enq_valid),
    .io_enq_bits(q_335_io_enq_bits),
    .io_deq_ready(q_335_io_deq_ready),
    .io_deq_valid(q_335_io_deq_valid),
    .io_deq_bits(q_335_io_deq_bits)
  );
  Queue q_336 ( // @[Decoupled.scala 361:21]
    .clock(q_336_clock),
    .reset(q_336_reset),
    .io_enq_ready(q_336_io_enq_ready),
    .io_enq_valid(q_336_io_enq_valid),
    .io_enq_bits(q_336_io_enq_bits),
    .io_deq_ready(q_336_io_deq_ready),
    .io_deq_valid(q_336_io_deq_valid),
    .io_deq_bits(q_336_io_deq_bits)
  );
  Queue q_337 ( // @[Decoupled.scala 361:21]
    .clock(q_337_clock),
    .reset(q_337_reset),
    .io_enq_ready(q_337_io_enq_ready),
    .io_enq_valid(q_337_io_enq_valid),
    .io_enq_bits(q_337_io_enq_bits),
    .io_deq_ready(q_337_io_deq_ready),
    .io_deq_valid(q_337_io_deq_valid),
    .io_deq_bits(q_337_io_deq_bits)
  );
  Queue q_338 ( // @[Decoupled.scala 361:21]
    .clock(q_338_clock),
    .reset(q_338_reset),
    .io_enq_ready(q_338_io_enq_ready),
    .io_enq_valid(q_338_io_enq_valid),
    .io_enq_bits(q_338_io_enq_bits),
    .io_deq_ready(q_338_io_deq_ready),
    .io_deq_valid(q_338_io_deq_valid),
    .io_deq_bits(q_338_io_deq_bits)
  );
  Queue q_339 ( // @[Decoupled.scala 361:21]
    .clock(q_339_clock),
    .reset(q_339_reset),
    .io_enq_ready(q_339_io_enq_ready),
    .io_enq_valid(q_339_io_enq_valid),
    .io_enq_bits(q_339_io_enq_bits),
    .io_deq_ready(q_339_io_deq_ready),
    .io_deq_valid(q_339_io_deq_valid),
    .io_deq_bits(q_339_io_deq_bits)
  );
  Queue q_340 ( // @[Decoupled.scala 361:21]
    .clock(q_340_clock),
    .reset(q_340_reset),
    .io_enq_ready(q_340_io_enq_ready),
    .io_enq_valid(q_340_io_enq_valid),
    .io_enq_bits(q_340_io_enq_bits),
    .io_deq_ready(q_340_io_deq_ready),
    .io_deq_valid(q_340_io_deq_valid),
    .io_deq_bits(q_340_io_deq_bits)
  );
  Queue q_341 ( // @[Decoupled.scala 361:21]
    .clock(q_341_clock),
    .reset(q_341_reset),
    .io_enq_ready(q_341_io_enq_ready),
    .io_enq_valid(q_341_io_enq_valid),
    .io_enq_bits(q_341_io_enq_bits),
    .io_deq_ready(q_341_io_deq_ready),
    .io_deq_valid(q_341_io_deq_valid),
    .io_deq_bits(q_341_io_deq_bits)
  );
  Queue q_342 ( // @[Decoupled.scala 361:21]
    .clock(q_342_clock),
    .reset(q_342_reset),
    .io_enq_ready(q_342_io_enq_ready),
    .io_enq_valid(q_342_io_enq_valid),
    .io_enq_bits(q_342_io_enq_bits),
    .io_deq_ready(q_342_io_deq_ready),
    .io_deq_valid(q_342_io_deq_valid),
    .io_deq_bits(q_342_io_deq_bits)
  );
  Queue q_343 ( // @[Decoupled.scala 361:21]
    .clock(q_343_clock),
    .reset(q_343_reset),
    .io_enq_ready(q_343_io_enq_ready),
    .io_enq_valid(q_343_io_enq_valid),
    .io_enq_bits(q_343_io_enq_bits),
    .io_deq_ready(q_343_io_deq_ready),
    .io_deq_valid(q_343_io_deq_valid),
    .io_deq_bits(q_343_io_deq_bits)
  );
  Queue q_344 ( // @[Decoupled.scala 361:21]
    .clock(q_344_clock),
    .reset(q_344_reset),
    .io_enq_ready(q_344_io_enq_ready),
    .io_enq_valid(q_344_io_enq_valid),
    .io_enq_bits(q_344_io_enq_bits),
    .io_deq_ready(q_344_io_deq_ready),
    .io_deq_valid(q_344_io_deq_valid),
    .io_deq_bits(q_344_io_deq_bits)
  );
  Queue q_345 ( // @[Decoupled.scala 361:21]
    .clock(q_345_clock),
    .reset(q_345_reset),
    .io_enq_ready(q_345_io_enq_ready),
    .io_enq_valid(q_345_io_enq_valid),
    .io_enq_bits(q_345_io_enq_bits),
    .io_deq_ready(q_345_io_deq_ready),
    .io_deq_valid(q_345_io_deq_valid),
    .io_deq_bits(q_345_io_deq_bits)
  );
  Queue q_346 ( // @[Decoupled.scala 361:21]
    .clock(q_346_clock),
    .reset(q_346_reset),
    .io_enq_ready(q_346_io_enq_ready),
    .io_enq_valid(q_346_io_enq_valid),
    .io_enq_bits(q_346_io_enq_bits),
    .io_deq_ready(q_346_io_deq_ready),
    .io_deq_valid(q_346_io_deq_valid),
    .io_deq_bits(q_346_io_deq_bits)
  );
  Queue q_347 ( // @[Decoupled.scala 361:21]
    .clock(q_347_clock),
    .reset(q_347_reset),
    .io_enq_ready(q_347_io_enq_ready),
    .io_enq_valid(q_347_io_enq_valid),
    .io_enq_bits(q_347_io_enq_bits),
    .io_deq_ready(q_347_io_deq_ready),
    .io_deq_valid(q_347_io_deq_valid),
    .io_deq_bits(q_347_io_deq_bits)
  );
  Queue q_348 ( // @[Decoupled.scala 361:21]
    .clock(q_348_clock),
    .reset(q_348_reset),
    .io_enq_ready(q_348_io_enq_ready),
    .io_enq_valid(q_348_io_enq_valid),
    .io_enq_bits(q_348_io_enq_bits),
    .io_deq_ready(q_348_io_deq_ready),
    .io_deq_valid(q_348_io_deq_valid),
    .io_deq_bits(q_348_io_deq_bits)
  );
  Queue q_349 ( // @[Decoupled.scala 361:21]
    .clock(q_349_clock),
    .reset(q_349_reset),
    .io_enq_ready(q_349_io_enq_ready),
    .io_enq_valid(q_349_io_enq_valid),
    .io_enq_bits(q_349_io_enq_bits),
    .io_deq_ready(q_349_io_deq_ready),
    .io_deq_valid(q_349_io_deq_valid),
    .io_deq_bits(q_349_io_deq_bits)
  );
  Queue q_350 ( // @[Decoupled.scala 361:21]
    .clock(q_350_clock),
    .reset(q_350_reset),
    .io_enq_ready(q_350_io_enq_ready),
    .io_enq_valid(q_350_io_enq_valid),
    .io_enq_bits(q_350_io_enq_bits),
    .io_deq_ready(q_350_io_deq_ready),
    .io_deq_valid(q_350_io_deq_valid),
    .io_deq_bits(q_350_io_deq_bits)
  );
  Queue q_351 ( // @[Decoupled.scala 361:21]
    .clock(q_351_clock),
    .reset(q_351_reset),
    .io_enq_ready(q_351_io_enq_ready),
    .io_enq_valid(q_351_io_enq_valid),
    .io_enq_bits(q_351_io_enq_bits),
    .io_deq_ready(q_351_io_deq_ready),
    .io_deq_valid(q_351_io_deq_valid),
    .io_deq_bits(q_351_io_deq_bits)
  );
  Queue q_352 ( // @[Decoupled.scala 361:21]
    .clock(q_352_clock),
    .reset(q_352_reset),
    .io_enq_ready(q_352_io_enq_ready),
    .io_enq_valid(q_352_io_enq_valid),
    .io_enq_bits(q_352_io_enq_bits),
    .io_deq_ready(q_352_io_deq_ready),
    .io_deq_valid(q_352_io_deq_valid),
    .io_deq_bits(q_352_io_deq_bits)
  );
  Queue q_353 ( // @[Decoupled.scala 361:21]
    .clock(q_353_clock),
    .reset(q_353_reset),
    .io_enq_ready(q_353_io_enq_ready),
    .io_enq_valid(q_353_io_enq_valid),
    .io_enq_bits(q_353_io_enq_bits),
    .io_deq_ready(q_353_io_deq_ready),
    .io_deq_valid(q_353_io_deq_valid),
    .io_deq_bits(q_353_io_deq_bits)
  );
  Queue q_354 ( // @[Decoupled.scala 361:21]
    .clock(q_354_clock),
    .reset(q_354_reset),
    .io_enq_ready(q_354_io_enq_ready),
    .io_enq_valid(q_354_io_enq_valid),
    .io_enq_bits(q_354_io_enq_bits),
    .io_deq_ready(q_354_io_deq_ready),
    .io_deq_valid(q_354_io_deq_valid),
    .io_deq_bits(q_354_io_deq_bits)
  );
  Queue q_355 ( // @[Decoupled.scala 361:21]
    .clock(q_355_clock),
    .reset(q_355_reset),
    .io_enq_ready(q_355_io_enq_ready),
    .io_enq_valid(q_355_io_enq_valid),
    .io_enq_bits(q_355_io_enq_bits),
    .io_deq_ready(q_355_io_deq_ready),
    .io_deq_valid(q_355_io_deq_valid),
    .io_deq_bits(q_355_io_deq_bits)
  );
  Queue q_356 ( // @[Decoupled.scala 361:21]
    .clock(q_356_clock),
    .reset(q_356_reset),
    .io_enq_ready(q_356_io_enq_ready),
    .io_enq_valid(q_356_io_enq_valid),
    .io_enq_bits(q_356_io_enq_bits),
    .io_deq_ready(q_356_io_deq_ready),
    .io_deq_valid(q_356_io_deq_valid),
    .io_deq_bits(q_356_io_deq_bits)
  );
  Queue q_357 ( // @[Decoupled.scala 361:21]
    .clock(q_357_clock),
    .reset(q_357_reset),
    .io_enq_ready(q_357_io_enq_ready),
    .io_enq_valid(q_357_io_enq_valid),
    .io_enq_bits(q_357_io_enq_bits),
    .io_deq_ready(q_357_io_deq_ready),
    .io_deq_valid(q_357_io_deq_valid),
    .io_deq_bits(q_357_io_deq_bits)
  );
  Queue q_358 ( // @[Decoupled.scala 361:21]
    .clock(q_358_clock),
    .reset(q_358_reset),
    .io_enq_ready(q_358_io_enq_ready),
    .io_enq_valid(q_358_io_enq_valid),
    .io_enq_bits(q_358_io_enq_bits),
    .io_deq_ready(q_358_io_deq_ready),
    .io_deq_valid(q_358_io_deq_valid),
    .io_deq_bits(q_358_io_deq_bits)
  );
  Queue q_359 ( // @[Decoupled.scala 361:21]
    .clock(q_359_clock),
    .reset(q_359_reset),
    .io_enq_ready(q_359_io_enq_ready),
    .io_enq_valid(q_359_io_enq_valid),
    .io_enq_bits(q_359_io_enq_bits),
    .io_deq_ready(q_359_io_deq_ready),
    .io_deq_valid(q_359_io_deq_valid),
    .io_deq_bits(q_359_io_deq_bits)
  );
  Queue q_360 ( // @[Decoupled.scala 361:21]
    .clock(q_360_clock),
    .reset(q_360_reset),
    .io_enq_ready(q_360_io_enq_ready),
    .io_enq_valid(q_360_io_enq_valid),
    .io_enq_bits(q_360_io_enq_bits),
    .io_deq_ready(q_360_io_deq_ready),
    .io_deq_valid(q_360_io_deq_valid),
    .io_deq_bits(q_360_io_deq_bits)
  );
  Queue q_361 ( // @[Decoupled.scala 361:21]
    .clock(q_361_clock),
    .reset(q_361_reset),
    .io_enq_ready(q_361_io_enq_ready),
    .io_enq_valid(q_361_io_enq_valid),
    .io_enq_bits(q_361_io_enq_bits),
    .io_deq_ready(q_361_io_deq_ready),
    .io_deq_valid(q_361_io_deq_valid),
    .io_deq_bits(q_361_io_deq_bits)
  );
  Queue q_362 ( // @[Decoupled.scala 361:21]
    .clock(q_362_clock),
    .reset(q_362_reset),
    .io_enq_ready(q_362_io_enq_ready),
    .io_enq_valid(q_362_io_enq_valid),
    .io_enq_bits(q_362_io_enq_bits),
    .io_deq_ready(q_362_io_deq_ready),
    .io_deq_valid(q_362_io_deq_valid),
    .io_deq_bits(q_362_io_deq_bits)
  );
  Queue q_363 ( // @[Decoupled.scala 361:21]
    .clock(q_363_clock),
    .reset(q_363_reset),
    .io_enq_ready(q_363_io_enq_ready),
    .io_enq_valid(q_363_io_enq_valid),
    .io_enq_bits(q_363_io_enq_bits),
    .io_deq_ready(q_363_io_deq_ready),
    .io_deq_valid(q_363_io_deq_valid),
    .io_deq_bits(q_363_io_deq_bits)
  );
  Queue q_364 ( // @[Decoupled.scala 361:21]
    .clock(q_364_clock),
    .reset(q_364_reset),
    .io_enq_ready(q_364_io_enq_ready),
    .io_enq_valid(q_364_io_enq_valid),
    .io_enq_bits(q_364_io_enq_bits),
    .io_deq_ready(q_364_io_deq_ready),
    .io_deq_valid(q_364_io_deq_valid),
    .io_deq_bits(q_364_io_deq_bits)
  );
  Queue q_365 ( // @[Decoupled.scala 361:21]
    .clock(q_365_clock),
    .reset(q_365_reset),
    .io_enq_ready(q_365_io_enq_ready),
    .io_enq_valid(q_365_io_enq_valid),
    .io_enq_bits(q_365_io_enq_bits),
    .io_deq_ready(q_365_io_deq_ready),
    .io_deq_valid(q_365_io_deq_valid),
    .io_deq_bits(q_365_io_deq_bits)
  );
  Queue q_366 ( // @[Decoupled.scala 361:21]
    .clock(q_366_clock),
    .reset(q_366_reset),
    .io_enq_ready(q_366_io_enq_ready),
    .io_enq_valid(q_366_io_enq_valid),
    .io_enq_bits(q_366_io_enq_bits),
    .io_deq_ready(q_366_io_deq_ready),
    .io_deq_valid(q_366_io_deq_valid),
    .io_deq_bits(q_366_io_deq_bits)
  );
  Queue q_367 ( // @[Decoupled.scala 361:21]
    .clock(q_367_clock),
    .reset(q_367_reset),
    .io_enq_ready(q_367_io_enq_ready),
    .io_enq_valid(q_367_io_enq_valid),
    .io_enq_bits(q_367_io_enq_bits),
    .io_deq_ready(q_367_io_deq_ready),
    .io_deq_valid(q_367_io_deq_valid),
    .io_deq_bits(q_367_io_deq_bits)
  );
  Queue q_368 ( // @[Decoupled.scala 361:21]
    .clock(q_368_clock),
    .reset(q_368_reset),
    .io_enq_ready(q_368_io_enq_ready),
    .io_enq_valid(q_368_io_enq_valid),
    .io_enq_bits(q_368_io_enq_bits),
    .io_deq_ready(q_368_io_deq_ready),
    .io_deq_valid(q_368_io_deq_valid),
    .io_deq_bits(q_368_io_deq_bits)
  );
  Queue q_369 ( // @[Decoupled.scala 361:21]
    .clock(q_369_clock),
    .reset(q_369_reset),
    .io_enq_ready(q_369_io_enq_ready),
    .io_enq_valid(q_369_io_enq_valid),
    .io_enq_bits(q_369_io_enq_bits),
    .io_deq_ready(q_369_io_deq_ready),
    .io_deq_valid(q_369_io_deq_valid),
    .io_deq_bits(q_369_io_deq_bits)
  );
  Queue q_370 ( // @[Decoupled.scala 361:21]
    .clock(q_370_clock),
    .reset(q_370_reset),
    .io_enq_ready(q_370_io_enq_ready),
    .io_enq_valid(q_370_io_enq_valid),
    .io_enq_bits(q_370_io_enq_bits),
    .io_deq_ready(q_370_io_deq_ready),
    .io_deq_valid(q_370_io_deq_valid),
    .io_deq_bits(q_370_io_deq_bits)
  );
  Queue q_371 ( // @[Decoupled.scala 361:21]
    .clock(q_371_clock),
    .reset(q_371_reset),
    .io_enq_ready(q_371_io_enq_ready),
    .io_enq_valid(q_371_io_enq_valid),
    .io_enq_bits(q_371_io_enq_bits),
    .io_deq_ready(q_371_io_deq_ready),
    .io_deq_valid(q_371_io_deq_valid),
    .io_deq_bits(q_371_io_deq_bits)
  );
  Queue q_372 ( // @[Decoupled.scala 361:21]
    .clock(q_372_clock),
    .reset(q_372_reset),
    .io_enq_ready(q_372_io_enq_ready),
    .io_enq_valid(q_372_io_enq_valid),
    .io_enq_bits(q_372_io_enq_bits),
    .io_deq_ready(q_372_io_deq_ready),
    .io_deq_valid(q_372_io_deq_valid),
    .io_deq_bits(q_372_io_deq_bits)
  );
  Queue q_373 ( // @[Decoupled.scala 361:21]
    .clock(q_373_clock),
    .reset(q_373_reset),
    .io_enq_ready(q_373_io_enq_ready),
    .io_enq_valid(q_373_io_enq_valid),
    .io_enq_bits(q_373_io_enq_bits),
    .io_deq_ready(q_373_io_deq_ready),
    .io_deq_valid(q_373_io_deq_valid),
    .io_deq_bits(q_373_io_deq_bits)
  );
  Queue q_374 ( // @[Decoupled.scala 361:21]
    .clock(q_374_clock),
    .reset(q_374_reset),
    .io_enq_ready(q_374_io_enq_ready),
    .io_enq_valid(q_374_io_enq_valid),
    .io_enq_bits(q_374_io_enq_bits),
    .io_deq_ready(q_374_io_deq_ready),
    .io_deq_valid(q_374_io_deq_valid),
    .io_deq_bits(q_374_io_deq_bits)
  );
  Queue q_375 ( // @[Decoupled.scala 361:21]
    .clock(q_375_clock),
    .reset(q_375_reset),
    .io_enq_ready(q_375_io_enq_ready),
    .io_enq_valid(q_375_io_enq_valid),
    .io_enq_bits(q_375_io_enq_bits),
    .io_deq_ready(q_375_io_deq_ready),
    .io_deq_valid(q_375_io_deq_valid),
    .io_deq_bits(q_375_io_deq_bits)
  );
  Queue q_376 ( // @[Decoupled.scala 361:21]
    .clock(q_376_clock),
    .reset(q_376_reset),
    .io_enq_ready(q_376_io_enq_ready),
    .io_enq_valid(q_376_io_enq_valid),
    .io_enq_bits(q_376_io_enq_bits),
    .io_deq_ready(q_376_io_deq_ready),
    .io_deq_valid(q_376_io_deq_valid),
    .io_deq_bits(q_376_io_deq_bits)
  );
  Queue q_377 ( // @[Decoupled.scala 361:21]
    .clock(q_377_clock),
    .reset(q_377_reset),
    .io_enq_ready(q_377_io_enq_ready),
    .io_enq_valid(q_377_io_enq_valid),
    .io_enq_bits(q_377_io_enq_bits),
    .io_deq_ready(q_377_io_deq_ready),
    .io_deq_valid(q_377_io_deq_valid),
    .io_deq_bits(q_377_io_deq_bits)
  );
  Queue q_378 ( // @[Decoupled.scala 361:21]
    .clock(q_378_clock),
    .reset(q_378_reset),
    .io_enq_ready(q_378_io_enq_ready),
    .io_enq_valid(q_378_io_enq_valid),
    .io_enq_bits(q_378_io_enq_bits),
    .io_deq_ready(q_378_io_deq_ready),
    .io_deq_valid(q_378_io_deq_valid),
    .io_deq_bits(q_378_io_deq_bits)
  );
  Queue q_379 ( // @[Decoupled.scala 361:21]
    .clock(q_379_clock),
    .reset(q_379_reset),
    .io_enq_ready(q_379_io_enq_ready),
    .io_enq_valid(q_379_io_enq_valid),
    .io_enq_bits(q_379_io_enq_bits),
    .io_deq_ready(q_379_io_deq_ready),
    .io_deq_valid(q_379_io_deq_valid),
    .io_deq_bits(q_379_io_deq_bits)
  );
  Queue q_380 ( // @[Decoupled.scala 361:21]
    .clock(q_380_clock),
    .reset(q_380_reset),
    .io_enq_ready(q_380_io_enq_ready),
    .io_enq_valid(q_380_io_enq_valid),
    .io_enq_bits(q_380_io_enq_bits),
    .io_deq_ready(q_380_io_deq_ready),
    .io_deq_valid(q_380_io_deq_valid),
    .io_deq_bits(q_380_io_deq_bits)
  );
  Queue q_381 ( // @[Decoupled.scala 361:21]
    .clock(q_381_clock),
    .reset(q_381_reset),
    .io_enq_ready(q_381_io_enq_ready),
    .io_enq_valid(q_381_io_enq_valid),
    .io_enq_bits(q_381_io_enq_bits),
    .io_deq_ready(q_381_io_deq_ready),
    .io_deq_valid(q_381_io_deq_valid),
    .io_deq_bits(q_381_io_deq_bits)
  );
  Queue q_382 ( // @[Decoupled.scala 361:21]
    .clock(q_382_clock),
    .reset(q_382_reset),
    .io_enq_ready(q_382_io_enq_ready),
    .io_enq_valid(q_382_io_enq_valid),
    .io_enq_bits(q_382_io_enq_bits),
    .io_deq_ready(q_382_io_deq_ready),
    .io_deq_valid(q_382_io_deq_valid),
    .io_deq_bits(q_382_io_deq_bits)
  );
  Queue q_383 ( // @[Decoupled.scala 361:21]
    .clock(q_383_clock),
    .reset(q_383_reset),
    .io_enq_ready(q_383_io_enq_ready),
    .io_enq_valid(q_383_io_enq_valid),
    .io_enq_bits(q_383_io_enq_bits),
    .io_deq_ready(q_383_io_deq_ready),
    .io_deq_valid(q_383_io_deq_valid),
    .io_deq_bits(q_383_io_deq_bits)
  );
  Queue q_384 ( // @[Decoupled.scala 361:21]
    .clock(q_384_clock),
    .reset(q_384_reset),
    .io_enq_ready(q_384_io_enq_ready),
    .io_enq_valid(q_384_io_enq_valid),
    .io_enq_bits(q_384_io_enq_bits),
    .io_deq_ready(q_384_io_deq_ready),
    .io_deq_valid(q_384_io_deq_valid),
    .io_deq_bits(q_384_io_deq_bits)
  );
  Queue q_385 ( // @[Decoupled.scala 361:21]
    .clock(q_385_clock),
    .reset(q_385_reset),
    .io_enq_ready(q_385_io_enq_ready),
    .io_enq_valid(q_385_io_enq_valid),
    .io_enq_bits(q_385_io_enq_bits),
    .io_deq_ready(q_385_io_deq_ready),
    .io_deq_valid(q_385_io_deq_valid),
    .io_deq_bits(q_385_io_deq_bits)
  );
  Queue q_386 ( // @[Decoupled.scala 361:21]
    .clock(q_386_clock),
    .reset(q_386_reset),
    .io_enq_ready(q_386_io_enq_ready),
    .io_enq_valid(q_386_io_enq_valid),
    .io_enq_bits(q_386_io_enq_bits),
    .io_deq_ready(q_386_io_deq_ready),
    .io_deq_valid(q_386_io_deq_valid),
    .io_deq_bits(q_386_io_deq_bits)
  );
  Queue q_387 ( // @[Decoupled.scala 361:21]
    .clock(q_387_clock),
    .reset(q_387_reset),
    .io_enq_ready(q_387_io_enq_ready),
    .io_enq_valid(q_387_io_enq_valid),
    .io_enq_bits(q_387_io_enq_bits),
    .io_deq_ready(q_387_io_deq_ready),
    .io_deq_valid(q_387_io_deq_valid),
    .io_deq_bits(q_387_io_deq_bits)
  );
  Queue q_388 ( // @[Decoupled.scala 361:21]
    .clock(q_388_clock),
    .reset(q_388_reset),
    .io_enq_ready(q_388_io_enq_ready),
    .io_enq_valid(q_388_io_enq_valid),
    .io_enq_bits(q_388_io_enq_bits),
    .io_deq_ready(q_388_io_deq_ready),
    .io_deq_valid(q_388_io_deq_valid),
    .io_deq_bits(q_388_io_deq_bits)
  );
  Queue q_389 ( // @[Decoupled.scala 361:21]
    .clock(q_389_clock),
    .reset(q_389_reset),
    .io_enq_ready(q_389_io_enq_ready),
    .io_enq_valid(q_389_io_enq_valid),
    .io_enq_bits(q_389_io_enq_bits),
    .io_deq_ready(q_389_io_deq_ready),
    .io_deq_valid(q_389_io_deq_valid),
    .io_deq_bits(q_389_io_deq_bits)
  );
  Queue q_390 ( // @[Decoupled.scala 361:21]
    .clock(q_390_clock),
    .reset(q_390_reset),
    .io_enq_ready(q_390_io_enq_ready),
    .io_enq_valid(q_390_io_enq_valid),
    .io_enq_bits(q_390_io_enq_bits),
    .io_deq_ready(q_390_io_deq_ready),
    .io_deq_valid(q_390_io_deq_valid),
    .io_deq_bits(q_390_io_deq_bits)
  );
  Queue q_391 ( // @[Decoupled.scala 361:21]
    .clock(q_391_clock),
    .reset(q_391_reset),
    .io_enq_ready(q_391_io_enq_ready),
    .io_enq_valid(q_391_io_enq_valid),
    .io_enq_bits(q_391_io_enq_bits),
    .io_deq_ready(q_391_io_deq_ready),
    .io_deq_valid(q_391_io_deq_valid),
    .io_deq_bits(q_391_io_deq_bits)
  );
  Queue q_392 ( // @[Decoupled.scala 361:21]
    .clock(q_392_clock),
    .reset(q_392_reset),
    .io_enq_ready(q_392_io_enq_ready),
    .io_enq_valid(q_392_io_enq_valid),
    .io_enq_bits(q_392_io_enq_bits),
    .io_deq_ready(q_392_io_deq_ready),
    .io_deq_valid(q_392_io_deq_valid),
    .io_deq_bits(q_392_io_deq_bits)
  );
  Queue q_393 ( // @[Decoupled.scala 361:21]
    .clock(q_393_clock),
    .reset(q_393_reset),
    .io_enq_ready(q_393_io_enq_ready),
    .io_enq_valid(q_393_io_enq_valid),
    .io_enq_bits(q_393_io_enq_bits),
    .io_deq_ready(q_393_io_deq_ready),
    .io_deq_valid(q_393_io_deq_valid),
    .io_deq_bits(q_393_io_deq_bits)
  );
  Queue q_394 ( // @[Decoupled.scala 361:21]
    .clock(q_394_clock),
    .reset(q_394_reset),
    .io_enq_ready(q_394_io_enq_ready),
    .io_enq_valid(q_394_io_enq_valid),
    .io_enq_bits(q_394_io_enq_bits),
    .io_deq_ready(q_394_io_deq_ready),
    .io_deq_valid(q_394_io_deq_valid),
    .io_deq_bits(q_394_io_deq_bits)
  );
  Queue q_395 ( // @[Decoupled.scala 361:21]
    .clock(q_395_clock),
    .reset(q_395_reset),
    .io_enq_ready(q_395_io_enq_ready),
    .io_enq_valid(q_395_io_enq_valid),
    .io_enq_bits(q_395_io_enq_bits),
    .io_deq_ready(q_395_io_deq_ready),
    .io_deq_valid(q_395_io_deq_valid),
    .io_deq_bits(q_395_io_deq_bits)
  );
  Queue q_396 ( // @[Decoupled.scala 361:21]
    .clock(q_396_clock),
    .reset(q_396_reset),
    .io_enq_ready(q_396_io_enq_ready),
    .io_enq_valid(q_396_io_enq_valid),
    .io_enq_bits(q_396_io_enq_bits),
    .io_deq_ready(q_396_io_deq_ready),
    .io_deq_valid(q_396_io_deq_valid),
    .io_deq_bits(q_396_io_deq_bits)
  );
  Queue q_397 ( // @[Decoupled.scala 361:21]
    .clock(q_397_clock),
    .reset(q_397_reset),
    .io_enq_ready(q_397_io_enq_ready),
    .io_enq_valid(q_397_io_enq_valid),
    .io_enq_bits(q_397_io_enq_bits),
    .io_deq_ready(q_397_io_deq_ready),
    .io_deq_valid(q_397_io_deq_valid),
    .io_deq_bits(q_397_io_deq_bits)
  );
  Queue q_398 ( // @[Decoupled.scala 361:21]
    .clock(q_398_clock),
    .reset(q_398_reset),
    .io_enq_ready(q_398_io_enq_ready),
    .io_enq_valid(q_398_io_enq_valid),
    .io_enq_bits(q_398_io_enq_bits),
    .io_deq_ready(q_398_io_deq_ready),
    .io_deq_valid(q_398_io_deq_valid),
    .io_deq_bits(q_398_io_deq_bits)
  );
  Queue q_399 ( // @[Decoupled.scala 361:21]
    .clock(q_399_clock),
    .reset(q_399_reset),
    .io_enq_ready(q_399_io_enq_ready),
    .io_enq_valid(q_399_io_enq_valid),
    .io_enq_bits(q_399_io_enq_bits),
    .io_deq_ready(q_399_io_deq_ready),
    .io_deq_valid(q_399_io_deq_valid),
    .io_deq_bits(q_399_io_deq_bits)
  );
  Queue q_400 ( // @[Decoupled.scala 361:21]
    .clock(q_400_clock),
    .reset(q_400_reset),
    .io_enq_ready(q_400_io_enq_ready),
    .io_enq_valid(q_400_io_enq_valid),
    .io_enq_bits(q_400_io_enq_bits),
    .io_deq_ready(q_400_io_deq_ready),
    .io_deq_valid(q_400_io_deq_valid),
    .io_deq_bits(q_400_io_deq_bits)
  );
  Queue q_401 ( // @[Decoupled.scala 361:21]
    .clock(q_401_clock),
    .reset(q_401_reset),
    .io_enq_ready(q_401_io_enq_ready),
    .io_enq_valid(q_401_io_enq_valid),
    .io_enq_bits(q_401_io_enq_bits),
    .io_deq_ready(q_401_io_deq_ready),
    .io_deq_valid(q_401_io_deq_valid),
    .io_deq_bits(q_401_io_deq_bits)
  );
  Queue q_402 ( // @[Decoupled.scala 361:21]
    .clock(q_402_clock),
    .reset(q_402_reset),
    .io_enq_ready(q_402_io_enq_ready),
    .io_enq_valid(q_402_io_enq_valid),
    .io_enq_bits(q_402_io_enq_bits),
    .io_deq_ready(q_402_io_deq_ready),
    .io_deq_valid(q_402_io_deq_valid),
    .io_deq_bits(q_402_io_deq_bits)
  );
  Queue q_403 ( // @[Decoupled.scala 361:21]
    .clock(q_403_clock),
    .reset(q_403_reset),
    .io_enq_ready(q_403_io_enq_ready),
    .io_enq_valid(q_403_io_enq_valid),
    .io_enq_bits(q_403_io_enq_bits),
    .io_deq_ready(q_403_io_deq_ready),
    .io_deq_valid(q_403_io_deq_valid),
    .io_deq_bits(q_403_io_deq_bits)
  );
  Queue q_404 ( // @[Decoupled.scala 361:21]
    .clock(q_404_clock),
    .reset(q_404_reset),
    .io_enq_ready(q_404_io_enq_ready),
    .io_enq_valid(q_404_io_enq_valid),
    .io_enq_bits(q_404_io_enq_bits),
    .io_deq_ready(q_404_io_deq_ready),
    .io_deq_valid(q_404_io_deq_valid),
    .io_deq_bits(q_404_io_deq_bits)
  );
  Queue q_405 ( // @[Decoupled.scala 361:21]
    .clock(q_405_clock),
    .reset(q_405_reset),
    .io_enq_ready(q_405_io_enq_ready),
    .io_enq_valid(q_405_io_enq_valid),
    .io_enq_bits(q_405_io_enq_bits),
    .io_deq_ready(q_405_io_deq_ready),
    .io_deq_valid(q_405_io_deq_valid),
    .io_deq_bits(q_405_io_deq_bits)
  );
  Queue q_406 ( // @[Decoupled.scala 361:21]
    .clock(q_406_clock),
    .reset(q_406_reset),
    .io_enq_ready(q_406_io_enq_ready),
    .io_enq_valid(q_406_io_enq_valid),
    .io_enq_bits(q_406_io_enq_bits),
    .io_deq_ready(q_406_io_deq_ready),
    .io_deq_valid(q_406_io_deq_valid),
    .io_deq_bits(q_406_io_deq_bits)
  );
  Queue q_407 ( // @[Decoupled.scala 361:21]
    .clock(q_407_clock),
    .reset(q_407_reset),
    .io_enq_ready(q_407_io_enq_ready),
    .io_enq_valid(q_407_io_enq_valid),
    .io_enq_bits(q_407_io_enq_bits),
    .io_deq_ready(q_407_io_deq_ready),
    .io_deq_valid(q_407_io_deq_valid),
    .io_deq_bits(q_407_io_deq_bits)
  );
  Queue q_408 ( // @[Decoupled.scala 361:21]
    .clock(q_408_clock),
    .reset(q_408_reset),
    .io_enq_ready(q_408_io_enq_ready),
    .io_enq_valid(q_408_io_enq_valid),
    .io_enq_bits(q_408_io_enq_bits),
    .io_deq_ready(q_408_io_deq_ready),
    .io_deq_valid(q_408_io_deq_valid),
    .io_deq_bits(q_408_io_deq_bits)
  );
  Queue q_409 ( // @[Decoupled.scala 361:21]
    .clock(q_409_clock),
    .reset(q_409_reset),
    .io_enq_ready(q_409_io_enq_ready),
    .io_enq_valid(q_409_io_enq_valid),
    .io_enq_bits(q_409_io_enq_bits),
    .io_deq_ready(q_409_io_deq_ready),
    .io_deq_valid(q_409_io_deq_valid),
    .io_deq_bits(q_409_io_deq_bits)
  );
  Queue q_410 ( // @[Decoupled.scala 361:21]
    .clock(q_410_clock),
    .reset(q_410_reset),
    .io_enq_ready(q_410_io_enq_ready),
    .io_enq_valid(q_410_io_enq_valid),
    .io_enq_bits(q_410_io_enq_bits),
    .io_deq_ready(q_410_io_deq_ready),
    .io_deq_valid(q_410_io_deq_valid),
    .io_deq_bits(q_410_io_deq_bits)
  );
  Queue q_411 ( // @[Decoupled.scala 361:21]
    .clock(q_411_clock),
    .reset(q_411_reset),
    .io_enq_ready(q_411_io_enq_ready),
    .io_enq_valid(q_411_io_enq_valid),
    .io_enq_bits(q_411_io_enq_bits),
    .io_deq_ready(q_411_io_deq_ready),
    .io_deq_valid(q_411_io_deq_valid),
    .io_deq_bits(q_411_io_deq_bits)
  );
  Queue q_412 ( // @[Decoupled.scala 361:21]
    .clock(q_412_clock),
    .reset(q_412_reset),
    .io_enq_ready(q_412_io_enq_ready),
    .io_enq_valid(q_412_io_enq_valid),
    .io_enq_bits(q_412_io_enq_bits),
    .io_deq_ready(q_412_io_deq_ready),
    .io_deq_valid(q_412_io_deq_valid),
    .io_deq_bits(q_412_io_deq_bits)
  );
  Queue q_413 ( // @[Decoupled.scala 361:21]
    .clock(q_413_clock),
    .reset(q_413_reset),
    .io_enq_ready(q_413_io_enq_ready),
    .io_enq_valid(q_413_io_enq_valid),
    .io_enq_bits(q_413_io_enq_bits),
    .io_deq_ready(q_413_io_deq_ready),
    .io_deq_valid(q_413_io_deq_valid),
    .io_deq_bits(q_413_io_deq_bits)
  );
  Queue q_414 ( // @[Decoupled.scala 361:21]
    .clock(q_414_clock),
    .reset(q_414_reset),
    .io_enq_ready(q_414_io_enq_ready),
    .io_enq_valid(q_414_io_enq_valid),
    .io_enq_bits(q_414_io_enq_bits),
    .io_deq_ready(q_414_io_deq_ready),
    .io_deq_valid(q_414_io_deq_valid),
    .io_deq_bits(q_414_io_deq_bits)
  );
  Queue q_415 ( // @[Decoupled.scala 361:21]
    .clock(q_415_clock),
    .reset(q_415_reset),
    .io_enq_ready(q_415_io_enq_ready),
    .io_enq_valid(q_415_io_enq_valid),
    .io_enq_bits(q_415_io_enq_bits),
    .io_deq_ready(q_415_io_deq_ready),
    .io_deq_valid(q_415_io_deq_valid),
    .io_deq_bits(q_415_io_deq_bits)
  );
  Queue q_416 ( // @[Decoupled.scala 361:21]
    .clock(q_416_clock),
    .reset(q_416_reset),
    .io_enq_ready(q_416_io_enq_ready),
    .io_enq_valid(q_416_io_enq_valid),
    .io_enq_bits(q_416_io_enq_bits),
    .io_deq_ready(q_416_io_deq_ready),
    .io_deq_valid(q_416_io_deq_valid),
    .io_deq_bits(q_416_io_deq_bits)
  );
  Queue q_417 ( // @[Decoupled.scala 361:21]
    .clock(q_417_clock),
    .reset(q_417_reset),
    .io_enq_ready(q_417_io_enq_ready),
    .io_enq_valid(q_417_io_enq_valid),
    .io_enq_bits(q_417_io_enq_bits),
    .io_deq_ready(q_417_io_deq_ready),
    .io_deq_valid(q_417_io_deq_valid),
    .io_deq_bits(q_417_io_deq_bits)
  );
  Queue q_418 ( // @[Decoupled.scala 361:21]
    .clock(q_418_clock),
    .reset(q_418_reset),
    .io_enq_ready(q_418_io_enq_ready),
    .io_enq_valid(q_418_io_enq_valid),
    .io_enq_bits(q_418_io_enq_bits),
    .io_deq_ready(q_418_io_deq_ready),
    .io_deq_valid(q_418_io_deq_valid),
    .io_deq_bits(q_418_io_deq_bits)
  );
  Queue q_419 ( // @[Decoupled.scala 361:21]
    .clock(q_419_clock),
    .reset(q_419_reset),
    .io_enq_ready(q_419_io_enq_ready),
    .io_enq_valid(q_419_io_enq_valid),
    .io_enq_bits(q_419_io_enq_bits),
    .io_deq_ready(q_419_io_deq_ready),
    .io_deq_valid(q_419_io_deq_valid),
    .io_deq_bits(q_419_io_deq_bits)
  );
  Queue q_420 ( // @[Decoupled.scala 361:21]
    .clock(q_420_clock),
    .reset(q_420_reset),
    .io_enq_ready(q_420_io_enq_ready),
    .io_enq_valid(q_420_io_enq_valid),
    .io_enq_bits(q_420_io_enq_bits),
    .io_deq_ready(q_420_io_deq_ready),
    .io_deq_valid(q_420_io_deq_valid),
    .io_deq_bits(q_420_io_deq_bits)
  );
  Queue q_421 ( // @[Decoupled.scala 361:21]
    .clock(q_421_clock),
    .reset(q_421_reset),
    .io_enq_ready(q_421_io_enq_ready),
    .io_enq_valid(q_421_io_enq_valid),
    .io_enq_bits(q_421_io_enq_bits),
    .io_deq_ready(q_421_io_deq_ready),
    .io_deq_valid(q_421_io_deq_valid),
    .io_deq_bits(q_421_io_deq_bits)
  );
  Queue q_422 ( // @[Decoupled.scala 361:21]
    .clock(q_422_clock),
    .reset(q_422_reset),
    .io_enq_ready(q_422_io_enq_ready),
    .io_enq_valid(q_422_io_enq_valid),
    .io_enq_bits(q_422_io_enq_bits),
    .io_deq_ready(q_422_io_deq_ready),
    .io_deq_valid(q_422_io_deq_valid),
    .io_deq_bits(q_422_io_deq_bits)
  );
  Queue q_423 ( // @[Decoupled.scala 361:21]
    .clock(q_423_clock),
    .reset(q_423_reset),
    .io_enq_ready(q_423_io_enq_ready),
    .io_enq_valid(q_423_io_enq_valid),
    .io_enq_bits(q_423_io_enq_bits),
    .io_deq_ready(q_423_io_deq_ready),
    .io_deq_valid(q_423_io_deq_valid),
    .io_deq_bits(q_423_io_deq_bits)
  );
  Queue q_424 ( // @[Decoupled.scala 361:21]
    .clock(q_424_clock),
    .reset(q_424_reset),
    .io_enq_ready(q_424_io_enq_ready),
    .io_enq_valid(q_424_io_enq_valid),
    .io_enq_bits(q_424_io_enq_bits),
    .io_deq_ready(q_424_io_deq_ready),
    .io_deq_valid(q_424_io_deq_valid),
    .io_deq_bits(q_424_io_deq_bits)
  );
  Queue q_425 ( // @[Decoupled.scala 361:21]
    .clock(q_425_clock),
    .reset(q_425_reset),
    .io_enq_ready(q_425_io_enq_ready),
    .io_enq_valid(q_425_io_enq_valid),
    .io_enq_bits(q_425_io_enq_bits),
    .io_deq_ready(q_425_io_deq_ready),
    .io_deq_valid(q_425_io_deq_valid),
    .io_deq_bits(q_425_io_deq_bits)
  );
  Queue q_426 ( // @[Decoupled.scala 361:21]
    .clock(q_426_clock),
    .reset(q_426_reset),
    .io_enq_ready(q_426_io_enq_ready),
    .io_enq_valid(q_426_io_enq_valid),
    .io_enq_bits(q_426_io_enq_bits),
    .io_deq_ready(q_426_io_deq_ready),
    .io_deq_valid(q_426_io_deq_valid),
    .io_deq_bits(q_426_io_deq_bits)
  );
  Queue q_427 ( // @[Decoupled.scala 361:21]
    .clock(q_427_clock),
    .reset(q_427_reset),
    .io_enq_ready(q_427_io_enq_ready),
    .io_enq_valid(q_427_io_enq_valid),
    .io_enq_bits(q_427_io_enq_bits),
    .io_deq_ready(q_427_io_deq_ready),
    .io_deq_valid(q_427_io_deq_valid),
    .io_deq_bits(q_427_io_deq_bits)
  );
  Queue q_428 ( // @[Decoupled.scala 361:21]
    .clock(q_428_clock),
    .reset(q_428_reset),
    .io_enq_ready(q_428_io_enq_ready),
    .io_enq_valid(q_428_io_enq_valid),
    .io_enq_bits(q_428_io_enq_bits),
    .io_deq_ready(q_428_io_deq_ready),
    .io_deq_valid(q_428_io_deq_valid),
    .io_deq_bits(q_428_io_deq_bits)
  );
  Queue q_429 ( // @[Decoupled.scala 361:21]
    .clock(q_429_clock),
    .reset(q_429_reset),
    .io_enq_ready(q_429_io_enq_ready),
    .io_enq_valid(q_429_io_enq_valid),
    .io_enq_bits(q_429_io_enq_bits),
    .io_deq_ready(q_429_io_deq_ready),
    .io_deq_valid(q_429_io_deq_valid),
    .io_deq_bits(q_429_io_deq_bits)
  );
  Queue q_430 ( // @[Decoupled.scala 361:21]
    .clock(q_430_clock),
    .reset(q_430_reset),
    .io_enq_ready(q_430_io_enq_ready),
    .io_enq_valid(q_430_io_enq_valid),
    .io_enq_bits(q_430_io_enq_bits),
    .io_deq_ready(q_430_io_deq_ready),
    .io_deq_valid(q_430_io_deq_valid),
    .io_deq_bits(q_430_io_deq_bits)
  );
  Queue q_431 ( // @[Decoupled.scala 361:21]
    .clock(q_431_clock),
    .reset(q_431_reset),
    .io_enq_ready(q_431_io_enq_ready),
    .io_enq_valid(q_431_io_enq_valid),
    .io_enq_bits(q_431_io_enq_bits),
    .io_deq_ready(q_431_io_deq_ready),
    .io_deq_valid(q_431_io_deq_valid),
    .io_deq_bits(q_431_io_deq_bits)
  );
  Queue q_432 ( // @[Decoupled.scala 361:21]
    .clock(q_432_clock),
    .reset(q_432_reset),
    .io_enq_ready(q_432_io_enq_ready),
    .io_enq_valid(q_432_io_enq_valid),
    .io_enq_bits(q_432_io_enq_bits),
    .io_deq_ready(q_432_io_deq_ready),
    .io_deq_valid(q_432_io_deq_valid),
    .io_deq_bits(q_432_io_deq_bits)
  );
  Queue q_433 ( // @[Decoupled.scala 361:21]
    .clock(q_433_clock),
    .reset(q_433_reset),
    .io_enq_ready(q_433_io_enq_ready),
    .io_enq_valid(q_433_io_enq_valid),
    .io_enq_bits(q_433_io_enq_bits),
    .io_deq_ready(q_433_io_deq_ready),
    .io_deq_valid(q_433_io_deq_valid),
    .io_deq_bits(q_433_io_deq_bits)
  );
  Queue q_434 ( // @[Decoupled.scala 361:21]
    .clock(q_434_clock),
    .reset(q_434_reset),
    .io_enq_ready(q_434_io_enq_ready),
    .io_enq_valid(q_434_io_enq_valid),
    .io_enq_bits(q_434_io_enq_bits),
    .io_deq_ready(q_434_io_deq_ready),
    .io_deq_valid(q_434_io_deq_valid),
    .io_deq_bits(q_434_io_deq_bits)
  );
  Queue q_435 ( // @[Decoupled.scala 361:21]
    .clock(q_435_clock),
    .reset(q_435_reset),
    .io_enq_ready(q_435_io_enq_ready),
    .io_enq_valid(q_435_io_enq_valid),
    .io_enq_bits(q_435_io_enq_bits),
    .io_deq_ready(q_435_io_deq_ready),
    .io_deq_valid(q_435_io_deq_valid),
    .io_deq_bits(q_435_io_deq_bits)
  );
  Queue q_436 ( // @[Decoupled.scala 361:21]
    .clock(q_436_clock),
    .reset(q_436_reset),
    .io_enq_ready(q_436_io_enq_ready),
    .io_enq_valid(q_436_io_enq_valid),
    .io_enq_bits(q_436_io_enq_bits),
    .io_deq_ready(q_436_io_deq_ready),
    .io_deq_valid(q_436_io_deq_valid),
    .io_deq_bits(q_436_io_deq_bits)
  );
  Queue q_437 ( // @[Decoupled.scala 361:21]
    .clock(q_437_clock),
    .reset(q_437_reset),
    .io_enq_ready(q_437_io_enq_ready),
    .io_enq_valid(q_437_io_enq_valid),
    .io_enq_bits(q_437_io_enq_bits),
    .io_deq_ready(q_437_io_deq_ready),
    .io_deq_valid(q_437_io_deq_valid),
    .io_deq_bits(q_437_io_deq_bits)
  );
  Queue q_438 ( // @[Decoupled.scala 361:21]
    .clock(q_438_clock),
    .reset(q_438_reset),
    .io_enq_ready(q_438_io_enq_ready),
    .io_enq_valid(q_438_io_enq_valid),
    .io_enq_bits(q_438_io_enq_bits),
    .io_deq_ready(q_438_io_deq_ready),
    .io_deq_valid(q_438_io_deq_valid),
    .io_deq_bits(q_438_io_deq_bits)
  );
  Queue q_439 ( // @[Decoupled.scala 361:21]
    .clock(q_439_clock),
    .reset(q_439_reset),
    .io_enq_ready(q_439_io_enq_ready),
    .io_enq_valid(q_439_io_enq_valid),
    .io_enq_bits(q_439_io_enq_bits),
    .io_deq_ready(q_439_io_deq_ready),
    .io_deq_valid(q_439_io_deq_valid),
    .io_deq_bits(q_439_io_deq_bits)
  );
  Queue q_440 ( // @[Decoupled.scala 361:21]
    .clock(q_440_clock),
    .reset(q_440_reset),
    .io_enq_ready(q_440_io_enq_ready),
    .io_enq_valid(q_440_io_enq_valid),
    .io_enq_bits(q_440_io_enq_bits),
    .io_deq_ready(q_440_io_deq_ready),
    .io_deq_valid(q_440_io_deq_valid),
    .io_deq_bits(q_440_io_deq_bits)
  );
  Queue q_441 ( // @[Decoupled.scala 361:21]
    .clock(q_441_clock),
    .reset(q_441_reset),
    .io_enq_ready(q_441_io_enq_ready),
    .io_enq_valid(q_441_io_enq_valid),
    .io_enq_bits(q_441_io_enq_bits),
    .io_deq_ready(q_441_io_deq_ready),
    .io_deq_valid(q_441_io_deq_valid),
    .io_deq_bits(q_441_io_deq_bits)
  );
  Queue q_442 ( // @[Decoupled.scala 361:21]
    .clock(q_442_clock),
    .reset(q_442_reset),
    .io_enq_ready(q_442_io_enq_ready),
    .io_enq_valid(q_442_io_enq_valid),
    .io_enq_bits(q_442_io_enq_bits),
    .io_deq_ready(q_442_io_deq_ready),
    .io_deq_valid(q_442_io_deq_valid),
    .io_deq_bits(q_442_io_deq_bits)
  );
  Queue q_443 ( // @[Decoupled.scala 361:21]
    .clock(q_443_clock),
    .reset(q_443_reset),
    .io_enq_ready(q_443_io_enq_ready),
    .io_enq_valid(q_443_io_enq_valid),
    .io_enq_bits(q_443_io_enq_bits),
    .io_deq_ready(q_443_io_deq_ready),
    .io_deq_valid(q_443_io_deq_valid),
    .io_deq_bits(q_443_io_deq_bits)
  );
  Queue q_444 ( // @[Decoupled.scala 361:21]
    .clock(q_444_clock),
    .reset(q_444_reset),
    .io_enq_ready(q_444_io_enq_ready),
    .io_enq_valid(q_444_io_enq_valid),
    .io_enq_bits(q_444_io_enq_bits),
    .io_deq_ready(q_444_io_deq_ready),
    .io_deq_valid(q_444_io_deq_valid),
    .io_deq_bits(q_444_io_deq_bits)
  );
  Queue q_445 ( // @[Decoupled.scala 361:21]
    .clock(q_445_clock),
    .reset(q_445_reset),
    .io_enq_ready(q_445_io_enq_ready),
    .io_enq_valid(q_445_io_enq_valid),
    .io_enq_bits(q_445_io_enq_bits),
    .io_deq_ready(q_445_io_deq_ready),
    .io_deq_valid(q_445_io_deq_valid),
    .io_deq_bits(q_445_io_deq_bits)
  );
  Queue q_446 ( // @[Decoupled.scala 361:21]
    .clock(q_446_clock),
    .reset(q_446_reset),
    .io_enq_ready(q_446_io_enq_ready),
    .io_enq_valid(q_446_io_enq_valid),
    .io_enq_bits(q_446_io_enq_bits),
    .io_deq_ready(q_446_io_deq_ready),
    .io_deq_valid(q_446_io_deq_valid),
    .io_deq_bits(q_446_io_deq_bits)
  );
  Queue q_447 ( // @[Decoupled.scala 361:21]
    .clock(q_447_clock),
    .reset(q_447_reset),
    .io_enq_ready(q_447_io_enq_ready),
    .io_enq_valid(q_447_io_enq_valid),
    .io_enq_bits(q_447_io_enq_bits),
    .io_deq_ready(q_447_io_deq_ready),
    .io_deq_valid(q_447_io_deq_valid),
    .io_deq_bits(q_447_io_deq_bits)
  );
  Queue q_448 ( // @[Decoupled.scala 361:21]
    .clock(q_448_clock),
    .reset(q_448_reset),
    .io_enq_ready(q_448_io_enq_ready),
    .io_enq_valid(q_448_io_enq_valid),
    .io_enq_bits(q_448_io_enq_bits),
    .io_deq_ready(q_448_io_deq_ready),
    .io_deq_valid(q_448_io_deq_valid),
    .io_deq_bits(q_448_io_deq_bits)
  );
  Queue q_449 ( // @[Decoupled.scala 361:21]
    .clock(q_449_clock),
    .reset(q_449_reset),
    .io_enq_ready(q_449_io_enq_ready),
    .io_enq_valid(q_449_io_enq_valid),
    .io_enq_bits(q_449_io_enq_bits),
    .io_deq_ready(q_449_io_deq_ready),
    .io_deq_valid(q_449_io_deq_valid),
    .io_deq_bits(q_449_io_deq_bits)
  );
  Queue q_450 ( // @[Decoupled.scala 361:21]
    .clock(q_450_clock),
    .reset(q_450_reset),
    .io_enq_ready(q_450_io_enq_ready),
    .io_enq_valid(q_450_io_enq_valid),
    .io_enq_bits(q_450_io_enq_bits),
    .io_deq_ready(q_450_io_deq_ready),
    .io_deq_valid(q_450_io_deq_valid),
    .io_deq_bits(q_450_io_deq_bits)
  );
  Queue q_451 ( // @[Decoupled.scala 361:21]
    .clock(q_451_clock),
    .reset(q_451_reset),
    .io_enq_ready(q_451_io_enq_ready),
    .io_enq_valid(q_451_io_enq_valid),
    .io_enq_bits(q_451_io_enq_bits),
    .io_deq_ready(q_451_io_deq_ready),
    .io_deq_valid(q_451_io_deq_valid),
    .io_deq_bits(q_451_io_deq_bits)
  );
  Queue q_452 ( // @[Decoupled.scala 361:21]
    .clock(q_452_clock),
    .reset(q_452_reset),
    .io_enq_ready(q_452_io_enq_ready),
    .io_enq_valid(q_452_io_enq_valid),
    .io_enq_bits(q_452_io_enq_bits),
    .io_deq_ready(q_452_io_deq_ready),
    .io_deq_valid(q_452_io_deq_valid),
    .io_deq_bits(q_452_io_deq_bits)
  );
  Queue q_453 ( // @[Decoupled.scala 361:21]
    .clock(q_453_clock),
    .reset(q_453_reset),
    .io_enq_ready(q_453_io_enq_ready),
    .io_enq_valid(q_453_io_enq_valid),
    .io_enq_bits(q_453_io_enq_bits),
    .io_deq_ready(q_453_io_deq_ready),
    .io_deq_valid(q_453_io_deq_valid),
    .io_deq_bits(q_453_io_deq_bits)
  );
  Queue q_454 ( // @[Decoupled.scala 361:21]
    .clock(q_454_clock),
    .reset(q_454_reset),
    .io_enq_ready(q_454_io_enq_ready),
    .io_enq_valid(q_454_io_enq_valid),
    .io_enq_bits(q_454_io_enq_bits),
    .io_deq_ready(q_454_io_deq_ready),
    .io_deq_valid(q_454_io_deq_valid),
    .io_deq_bits(q_454_io_deq_bits)
  );
  Queue q_455 ( // @[Decoupled.scala 361:21]
    .clock(q_455_clock),
    .reset(q_455_reset),
    .io_enq_ready(q_455_io_enq_ready),
    .io_enq_valid(q_455_io_enq_valid),
    .io_enq_bits(q_455_io_enq_bits),
    .io_deq_ready(q_455_io_deq_ready),
    .io_deq_valid(q_455_io_deq_valid),
    .io_deq_bits(q_455_io_deq_bits)
  );
  Queue q_456 ( // @[Decoupled.scala 361:21]
    .clock(q_456_clock),
    .reset(q_456_reset),
    .io_enq_ready(q_456_io_enq_ready),
    .io_enq_valid(q_456_io_enq_valid),
    .io_enq_bits(q_456_io_enq_bits),
    .io_deq_ready(q_456_io_deq_ready),
    .io_deq_valid(q_456_io_deq_valid),
    .io_deq_bits(q_456_io_deq_bits)
  );
  Queue q_457 ( // @[Decoupled.scala 361:21]
    .clock(q_457_clock),
    .reset(q_457_reset),
    .io_enq_ready(q_457_io_enq_ready),
    .io_enq_valid(q_457_io_enq_valid),
    .io_enq_bits(q_457_io_enq_bits),
    .io_deq_ready(q_457_io_deq_ready),
    .io_deq_valid(q_457_io_deq_valid),
    .io_deq_bits(q_457_io_deq_bits)
  );
  Queue q_458 ( // @[Decoupled.scala 361:21]
    .clock(q_458_clock),
    .reset(q_458_reset),
    .io_enq_ready(q_458_io_enq_ready),
    .io_enq_valid(q_458_io_enq_valid),
    .io_enq_bits(q_458_io_enq_bits),
    .io_deq_ready(q_458_io_deq_ready),
    .io_deq_valid(q_458_io_deq_valid),
    .io_deq_bits(q_458_io_deq_bits)
  );
  Queue q_459 ( // @[Decoupled.scala 361:21]
    .clock(q_459_clock),
    .reset(q_459_reset),
    .io_enq_ready(q_459_io_enq_ready),
    .io_enq_valid(q_459_io_enq_valid),
    .io_enq_bits(q_459_io_enq_bits),
    .io_deq_ready(q_459_io_deq_ready),
    .io_deq_valid(q_459_io_deq_valid),
    .io_deq_bits(q_459_io_deq_bits)
  );
  Queue q_460 ( // @[Decoupled.scala 361:21]
    .clock(q_460_clock),
    .reset(q_460_reset),
    .io_enq_ready(q_460_io_enq_ready),
    .io_enq_valid(q_460_io_enq_valid),
    .io_enq_bits(q_460_io_enq_bits),
    .io_deq_ready(q_460_io_deq_ready),
    .io_deq_valid(q_460_io_deq_valid),
    .io_deq_bits(q_460_io_deq_bits)
  );
  Queue q_461 ( // @[Decoupled.scala 361:21]
    .clock(q_461_clock),
    .reset(q_461_reset),
    .io_enq_ready(q_461_io_enq_ready),
    .io_enq_valid(q_461_io_enq_valid),
    .io_enq_bits(q_461_io_enq_bits),
    .io_deq_ready(q_461_io_deq_ready),
    .io_deq_valid(q_461_io_deq_valid),
    .io_deq_bits(q_461_io_deq_bits)
  );
  Queue q_462 ( // @[Decoupled.scala 361:21]
    .clock(q_462_clock),
    .reset(q_462_reset),
    .io_enq_ready(q_462_io_enq_ready),
    .io_enq_valid(q_462_io_enq_valid),
    .io_enq_bits(q_462_io_enq_bits),
    .io_deq_ready(q_462_io_deq_ready),
    .io_deq_valid(q_462_io_deq_valid),
    .io_deq_bits(q_462_io_deq_bits)
  );
  Queue q_463 ( // @[Decoupled.scala 361:21]
    .clock(q_463_clock),
    .reset(q_463_reset),
    .io_enq_ready(q_463_io_enq_ready),
    .io_enq_valid(q_463_io_enq_valid),
    .io_enq_bits(q_463_io_enq_bits),
    .io_deq_ready(q_463_io_deq_ready),
    .io_deq_valid(q_463_io_deq_valid),
    .io_deq_bits(q_463_io_deq_bits)
  );
  Queue q_464 ( // @[Decoupled.scala 361:21]
    .clock(q_464_clock),
    .reset(q_464_reset),
    .io_enq_ready(q_464_io_enq_ready),
    .io_enq_valid(q_464_io_enq_valid),
    .io_enq_bits(q_464_io_enq_bits),
    .io_deq_ready(q_464_io_deq_ready),
    .io_deq_valid(q_464_io_deq_valid),
    .io_deq_bits(q_464_io_deq_bits)
  );
  Queue q_465 ( // @[Decoupled.scala 361:21]
    .clock(q_465_clock),
    .reset(q_465_reset),
    .io_enq_ready(q_465_io_enq_ready),
    .io_enq_valid(q_465_io_enq_valid),
    .io_enq_bits(q_465_io_enq_bits),
    .io_deq_ready(q_465_io_deq_ready),
    .io_deq_valid(q_465_io_deq_valid),
    .io_deq_bits(q_465_io_deq_bits)
  );
  Queue q_466 ( // @[Decoupled.scala 361:21]
    .clock(q_466_clock),
    .reset(q_466_reset),
    .io_enq_ready(q_466_io_enq_ready),
    .io_enq_valid(q_466_io_enq_valid),
    .io_enq_bits(q_466_io_enq_bits),
    .io_deq_ready(q_466_io_deq_ready),
    .io_deq_valid(q_466_io_deq_valid),
    .io_deq_bits(q_466_io_deq_bits)
  );
  Queue q_467 ( // @[Decoupled.scala 361:21]
    .clock(q_467_clock),
    .reset(q_467_reset),
    .io_enq_ready(q_467_io_enq_ready),
    .io_enq_valid(q_467_io_enq_valid),
    .io_enq_bits(q_467_io_enq_bits),
    .io_deq_ready(q_467_io_deq_ready),
    .io_deq_valid(q_467_io_deq_valid),
    .io_deq_bits(q_467_io_deq_bits)
  );
  Queue q_468 ( // @[Decoupled.scala 361:21]
    .clock(q_468_clock),
    .reset(q_468_reset),
    .io_enq_ready(q_468_io_enq_ready),
    .io_enq_valid(q_468_io_enq_valid),
    .io_enq_bits(q_468_io_enq_bits),
    .io_deq_ready(q_468_io_deq_ready),
    .io_deq_valid(q_468_io_deq_valid),
    .io_deq_bits(q_468_io_deq_bits)
  );
  Queue q_469 ( // @[Decoupled.scala 361:21]
    .clock(q_469_clock),
    .reset(q_469_reset),
    .io_enq_ready(q_469_io_enq_ready),
    .io_enq_valid(q_469_io_enq_valid),
    .io_enq_bits(q_469_io_enq_bits),
    .io_deq_ready(q_469_io_deq_ready),
    .io_deq_valid(q_469_io_deq_valid),
    .io_deq_bits(q_469_io_deq_bits)
  );
  Queue q_470 ( // @[Decoupled.scala 361:21]
    .clock(q_470_clock),
    .reset(q_470_reset),
    .io_enq_ready(q_470_io_enq_ready),
    .io_enq_valid(q_470_io_enq_valid),
    .io_enq_bits(q_470_io_enq_bits),
    .io_deq_ready(q_470_io_deq_ready),
    .io_deq_valid(q_470_io_deq_valid),
    .io_deq_bits(q_470_io_deq_bits)
  );
  Queue q_471 ( // @[Decoupled.scala 361:21]
    .clock(q_471_clock),
    .reset(q_471_reset),
    .io_enq_ready(q_471_io_enq_ready),
    .io_enq_valid(q_471_io_enq_valid),
    .io_enq_bits(q_471_io_enq_bits),
    .io_deq_ready(q_471_io_deq_ready),
    .io_deq_valid(q_471_io_deq_valid),
    .io_deq_bits(q_471_io_deq_bits)
  );
  Queue q_472 ( // @[Decoupled.scala 361:21]
    .clock(q_472_clock),
    .reset(q_472_reset),
    .io_enq_ready(q_472_io_enq_ready),
    .io_enq_valid(q_472_io_enq_valid),
    .io_enq_bits(q_472_io_enq_bits),
    .io_deq_ready(q_472_io_deq_ready),
    .io_deq_valid(q_472_io_deq_valid),
    .io_deq_bits(q_472_io_deq_bits)
  );
  Queue q_473 ( // @[Decoupled.scala 361:21]
    .clock(q_473_clock),
    .reset(q_473_reset),
    .io_enq_ready(q_473_io_enq_ready),
    .io_enq_valid(q_473_io_enq_valid),
    .io_enq_bits(q_473_io_enq_bits),
    .io_deq_ready(q_473_io_deq_ready),
    .io_deq_valid(q_473_io_deq_valid),
    .io_deq_bits(q_473_io_deq_bits)
  );
  Queue q_474 ( // @[Decoupled.scala 361:21]
    .clock(q_474_clock),
    .reset(q_474_reset),
    .io_enq_ready(q_474_io_enq_ready),
    .io_enq_valid(q_474_io_enq_valid),
    .io_enq_bits(q_474_io_enq_bits),
    .io_deq_ready(q_474_io_deq_ready),
    .io_deq_valid(q_474_io_deq_valid),
    .io_deq_bits(q_474_io_deq_bits)
  );
  Queue q_475 ( // @[Decoupled.scala 361:21]
    .clock(q_475_clock),
    .reset(q_475_reset),
    .io_enq_ready(q_475_io_enq_ready),
    .io_enq_valid(q_475_io_enq_valid),
    .io_enq_bits(q_475_io_enq_bits),
    .io_deq_ready(q_475_io_deq_ready),
    .io_deq_valid(q_475_io_deq_valid),
    .io_deq_bits(q_475_io_deq_bits)
  );
  Queue q_476 ( // @[Decoupled.scala 361:21]
    .clock(q_476_clock),
    .reset(q_476_reset),
    .io_enq_ready(q_476_io_enq_ready),
    .io_enq_valid(q_476_io_enq_valid),
    .io_enq_bits(q_476_io_enq_bits),
    .io_deq_ready(q_476_io_deq_ready),
    .io_deq_valid(q_476_io_deq_valid),
    .io_deq_bits(q_476_io_deq_bits)
  );
  Queue q_477 ( // @[Decoupled.scala 361:21]
    .clock(q_477_clock),
    .reset(q_477_reset),
    .io_enq_ready(q_477_io_enq_ready),
    .io_enq_valid(q_477_io_enq_valid),
    .io_enq_bits(q_477_io_enq_bits),
    .io_deq_ready(q_477_io_deq_ready),
    .io_deq_valid(q_477_io_deq_valid),
    .io_deq_bits(q_477_io_deq_bits)
  );
  Queue q_478 ( // @[Decoupled.scala 361:21]
    .clock(q_478_clock),
    .reset(q_478_reset),
    .io_enq_ready(q_478_io_enq_ready),
    .io_enq_valid(q_478_io_enq_valid),
    .io_enq_bits(q_478_io_enq_bits),
    .io_deq_ready(q_478_io_deq_ready),
    .io_deq_valid(q_478_io_deq_valid),
    .io_deq_bits(q_478_io_deq_bits)
  );
  Queue q_479 ( // @[Decoupled.scala 361:21]
    .clock(q_479_clock),
    .reset(q_479_reset),
    .io_enq_ready(q_479_io_enq_ready),
    .io_enq_valid(q_479_io_enq_valid),
    .io_enq_bits(q_479_io_enq_bits),
    .io_deq_ready(q_479_io_deq_ready),
    .io_deq_valid(q_479_io_deq_valid),
    .io_deq_bits(q_479_io_deq_bits)
  );
  Queue q_480 ( // @[Decoupled.scala 361:21]
    .clock(q_480_clock),
    .reset(q_480_reset),
    .io_enq_ready(q_480_io_enq_ready),
    .io_enq_valid(q_480_io_enq_valid),
    .io_enq_bits(q_480_io_enq_bits),
    .io_deq_ready(q_480_io_deq_ready),
    .io_deq_valid(q_480_io_deq_valid),
    .io_deq_bits(q_480_io_deq_bits)
  );
  Queue q_481 ( // @[Decoupled.scala 361:21]
    .clock(q_481_clock),
    .reset(q_481_reset),
    .io_enq_ready(q_481_io_enq_ready),
    .io_enq_valid(q_481_io_enq_valid),
    .io_enq_bits(q_481_io_enq_bits),
    .io_deq_ready(q_481_io_deq_ready),
    .io_deq_valid(q_481_io_deq_valid),
    .io_deq_bits(q_481_io_deq_bits)
  );
  Queue q_482 ( // @[Decoupled.scala 361:21]
    .clock(q_482_clock),
    .reset(q_482_reset),
    .io_enq_ready(q_482_io_enq_ready),
    .io_enq_valid(q_482_io_enq_valid),
    .io_enq_bits(q_482_io_enq_bits),
    .io_deq_ready(q_482_io_deq_ready),
    .io_deq_valid(q_482_io_deq_valid),
    .io_deq_bits(q_482_io_deq_bits)
  );
  Queue q_483 ( // @[Decoupled.scala 361:21]
    .clock(q_483_clock),
    .reset(q_483_reset),
    .io_enq_ready(q_483_io_enq_ready),
    .io_enq_valid(q_483_io_enq_valid),
    .io_enq_bits(q_483_io_enq_bits),
    .io_deq_ready(q_483_io_deq_ready),
    .io_deq_valid(q_483_io_deq_valid),
    .io_deq_bits(q_483_io_deq_bits)
  );
  Queue q_484 ( // @[Decoupled.scala 361:21]
    .clock(q_484_clock),
    .reset(q_484_reset),
    .io_enq_ready(q_484_io_enq_ready),
    .io_enq_valid(q_484_io_enq_valid),
    .io_enq_bits(q_484_io_enq_bits),
    .io_deq_ready(q_484_io_deq_ready),
    .io_deq_valid(q_484_io_deq_valid),
    .io_deq_bits(q_484_io_deq_bits)
  );
  Queue q_485 ( // @[Decoupled.scala 361:21]
    .clock(q_485_clock),
    .reset(q_485_reset),
    .io_enq_ready(q_485_io_enq_ready),
    .io_enq_valid(q_485_io_enq_valid),
    .io_enq_bits(q_485_io_enq_bits),
    .io_deq_ready(q_485_io_deq_ready),
    .io_deq_valid(q_485_io_deq_valid),
    .io_deq_bits(q_485_io_deq_bits)
  );
  Queue q_486 ( // @[Decoupled.scala 361:21]
    .clock(q_486_clock),
    .reset(q_486_reset),
    .io_enq_ready(q_486_io_enq_ready),
    .io_enq_valid(q_486_io_enq_valid),
    .io_enq_bits(q_486_io_enq_bits),
    .io_deq_ready(q_486_io_deq_ready),
    .io_deq_valid(q_486_io_deq_valid),
    .io_deq_bits(q_486_io_deq_bits)
  );
  Queue q_487 ( // @[Decoupled.scala 361:21]
    .clock(q_487_clock),
    .reset(q_487_reset),
    .io_enq_ready(q_487_io_enq_ready),
    .io_enq_valid(q_487_io_enq_valid),
    .io_enq_bits(q_487_io_enq_bits),
    .io_deq_ready(q_487_io_deq_ready),
    .io_deq_valid(q_487_io_deq_valid),
    .io_deq_bits(q_487_io_deq_bits)
  );
  Queue q_488 ( // @[Decoupled.scala 361:21]
    .clock(q_488_clock),
    .reset(q_488_reset),
    .io_enq_ready(q_488_io_enq_ready),
    .io_enq_valid(q_488_io_enq_valid),
    .io_enq_bits(q_488_io_enq_bits),
    .io_deq_ready(q_488_io_deq_ready),
    .io_deq_valid(q_488_io_deq_valid),
    .io_deq_bits(q_488_io_deq_bits)
  );
  Queue q_489 ( // @[Decoupled.scala 361:21]
    .clock(q_489_clock),
    .reset(q_489_reset),
    .io_enq_ready(q_489_io_enq_ready),
    .io_enq_valid(q_489_io_enq_valid),
    .io_enq_bits(q_489_io_enq_bits),
    .io_deq_ready(q_489_io_deq_ready),
    .io_deq_valid(q_489_io_deq_valid),
    .io_deq_bits(q_489_io_deq_bits)
  );
  Queue q_490 ( // @[Decoupled.scala 361:21]
    .clock(q_490_clock),
    .reset(q_490_reset),
    .io_enq_ready(q_490_io_enq_ready),
    .io_enq_valid(q_490_io_enq_valid),
    .io_enq_bits(q_490_io_enq_bits),
    .io_deq_ready(q_490_io_deq_ready),
    .io_deq_valid(q_490_io_deq_valid),
    .io_deq_bits(q_490_io_deq_bits)
  );
  Queue q_491 ( // @[Decoupled.scala 361:21]
    .clock(q_491_clock),
    .reset(q_491_reset),
    .io_enq_ready(q_491_io_enq_ready),
    .io_enq_valid(q_491_io_enq_valid),
    .io_enq_bits(q_491_io_enq_bits),
    .io_deq_ready(q_491_io_deq_ready),
    .io_deq_valid(q_491_io_deq_valid),
    .io_deq_bits(q_491_io_deq_bits)
  );
  Queue q_492 ( // @[Decoupled.scala 361:21]
    .clock(q_492_clock),
    .reset(q_492_reset),
    .io_enq_ready(q_492_io_enq_ready),
    .io_enq_valid(q_492_io_enq_valid),
    .io_enq_bits(q_492_io_enq_bits),
    .io_deq_ready(q_492_io_deq_ready),
    .io_deq_valid(q_492_io_deq_valid),
    .io_deq_bits(q_492_io_deq_bits)
  );
  Queue q_493 ( // @[Decoupled.scala 361:21]
    .clock(q_493_clock),
    .reset(q_493_reset),
    .io_enq_ready(q_493_io_enq_ready),
    .io_enq_valid(q_493_io_enq_valid),
    .io_enq_bits(q_493_io_enq_bits),
    .io_deq_ready(q_493_io_deq_ready),
    .io_deq_valid(q_493_io_deq_valid),
    .io_deq_bits(q_493_io_deq_bits)
  );
  Queue q_494 ( // @[Decoupled.scala 361:21]
    .clock(q_494_clock),
    .reset(q_494_reset),
    .io_enq_ready(q_494_io_enq_ready),
    .io_enq_valid(q_494_io_enq_valid),
    .io_enq_bits(q_494_io_enq_bits),
    .io_deq_ready(q_494_io_deq_ready),
    .io_deq_valid(q_494_io_deq_valid),
    .io_deq_bits(q_494_io_deq_bits)
  );
  Queue q_495 ( // @[Decoupled.scala 361:21]
    .clock(q_495_clock),
    .reset(q_495_reset),
    .io_enq_ready(q_495_io_enq_ready),
    .io_enq_valid(q_495_io_enq_valid),
    .io_enq_bits(q_495_io_enq_bits),
    .io_deq_ready(q_495_io_deq_ready),
    .io_deq_valid(q_495_io_deq_valid),
    .io_deq_bits(q_495_io_deq_bits)
  );
  Queue q_496 ( // @[Decoupled.scala 361:21]
    .clock(q_496_clock),
    .reset(q_496_reset),
    .io_enq_ready(q_496_io_enq_ready),
    .io_enq_valid(q_496_io_enq_valid),
    .io_enq_bits(q_496_io_enq_bits),
    .io_deq_ready(q_496_io_deq_ready),
    .io_deq_valid(q_496_io_deq_valid),
    .io_deq_bits(q_496_io_deq_bits)
  );
  Queue q_497 ( // @[Decoupled.scala 361:21]
    .clock(q_497_clock),
    .reset(q_497_reset),
    .io_enq_ready(q_497_io_enq_ready),
    .io_enq_valid(q_497_io_enq_valid),
    .io_enq_bits(q_497_io_enq_bits),
    .io_deq_ready(q_497_io_deq_ready),
    .io_deq_valid(q_497_io_deq_valid),
    .io_deq_bits(q_497_io_deq_bits)
  );
  Queue q_498 ( // @[Decoupled.scala 361:21]
    .clock(q_498_clock),
    .reset(q_498_reset),
    .io_enq_ready(q_498_io_enq_ready),
    .io_enq_valid(q_498_io_enq_valid),
    .io_enq_bits(q_498_io_enq_bits),
    .io_deq_ready(q_498_io_deq_ready),
    .io_deq_valid(q_498_io_deq_valid),
    .io_deq_bits(q_498_io_deq_bits)
  );
  Queue q_499 ( // @[Decoupled.scala 361:21]
    .clock(q_499_clock),
    .reset(q_499_reset),
    .io_enq_ready(q_499_io_enq_ready),
    .io_enq_valid(q_499_io_enq_valid),
    .io_enq_bits(q_499_io_enq_bits),
    .io_deq_ready(q_499_io_deq_ready),
    .io_deq_valid(q_499_io_deq_valid),
    .io_deq_bits(q_499_io_deq_bits)
  );
  Queue q_500 ( // @[Decoupled.scala 361:21]
    .clock(q_500_clock),
    .reset(q_500_reset),
    .io_enq_ready(q_500_io_enq_ready),
    .io_enq_valid(q_500_io_enq_valid),
    .io_enq_bits(q_500_io_enq_bits),
    .io_deq_ready(q_500_io_deq_ready),
    .io_deq_valid(q_500_io_deq_valid),
    .io_deq_bits(q_500_io_deq_bits)
  );
  Queue q_501 ( // @[Decoupled.scala 361:21]
    .clock(q_501_clock),
    .reset(q_501_reset),
    .io_enq_ready(q_501_io_enq_ready),
    .io_enq_valid(q_501_io_enq_valid),
    .io_enq_bits(q_501_io_enq_bits),
    .io_deq_ready(q_501_io_deq_ready),
    .io_deq_valid(q_501_io_deq_valid),
    .io_deq_bits(q_501_io_deq_bits)
  );
  Queue q_502 ( // @[Decoupled.scala 361:21]
    .clock(q_502_clock),
    .reset(q_502_reset),
    .io_enq_ready(q_502_io_enq_ready),
    .io_enq_valid(q_502_io_enq_valid),
    .io_enq_bits(q_502_io_enq_bits),
    .io_deq_ready(q_502_io_deq_ready),
    .io_deq_valid(q_502_io_deq_valid),
    .io_deq_bits(q_502_io_deq_bits)
  );
  Queue q_503 ( // @[Decoupled.scala 361:21]
    .clock(q_503_clock),
    .reset(q_503_reset),
    .io_enq_ready(q_503_io_enq_ready),
    .io_enq_valid(q_503_io_enq_valid),
    .io_enq_bits(q_503_io_enq_bits),
    .io_deq_ready(q_503_io_deq_ready),
    .io_deq_valid(q_503_io_deq_valid),
    .io_deq_bits(q_503_io_deq_bits)
  );
  Queue q_504 ( // @[Decoupled.scala 361:21]
    .clock(q_504_clock),
    .reset(q_504_reset),
    .io_enq_ready(q_504_io_enq_ready),
    .io_enq_valid(q_504_io_enq_valid),
    .io_enq_bits(q_504_io_enq_bits),
    .io_deq_ready(q_504_io_deq_ready),
    .io_deq_valid(q_504_io_deq_valid),
    .io_deq_bits(q_504_io_deq_bits)
  );
  Queue q_505 ( // @[Decoupled.scala 361:21]
    .clock(q_505_clock),
    .reset(q_505_reset),
    .io_enq_ready(q_505_io_enq_ready),
    .io_enq_valid(q_505_io_enq_valid),
    .io_enq_bits(q_505_io_enq_bits),
    .io_deq_ready(q_505_io_deq_ready),
    .io_deq_valid(q_505_io_deq_valid),
    .io_deq_bits(q_505_io_deq_bits)
  );
  Queue q_506 ( // @[Decoupled.scala 361:21]
    .clock(q_506_clock),
    .reset(q_506_reset),
    .io_enq_ready(q_506_io_enq_ready),
    .io_enq_valid(q_506_io_enq_valid),
    .io_enq_bits(q_506_io_enq_bits),
    .io_deq_ready(q_506_io_deq_ready),
    .io_deq_valid(q_506_io_deq_valid),
    .io_deq_bits(q_506_io_deq_bits)
  );
  Queue q_507 ( // @[Decoupled.scala 361:21]
    .clock(q_507_clock),
    .reset(q_507_reset),
    .io_enq_ready(q_507_io_enq_ready),
    .io_enq_valid(q_507_io_enq_valid),
    .io_enq_bits(q_507_io_enq_bits),
    .io_deq_ready(q_507_io_deq_ready),
    .io_deq_valid(q_507_io_deq_valid),
    .io_deq_bits(q_507_io_deq_bits)
  );
  Queue q_508 ( // @[Decoupled.scala 361:21]
    .clock(q_508_clock),
    .reset(q_508_reset),
    .io_enq_ready(q_508_io_enq_ready),
    .io_enq_valid(q_508_io_enq_valid),
    .io_enq_bits(q_508_io_enq_bits),
    .io_deq_ready(q_508_io_deq_ready),
    .io_deq_valid(q_508_io_deq_valid),
    .io_deq_bits(q_508_io_deq_bits)
  );
  Queue q_509 ( // @[Decoupled.scala 361:21]
    .clock(q_509_clock),
    .reset(q_509_reset),
    .io_enq_ready(q_509_io_enq_ready),
    .io_enq_valid(q_509_io_enq_valid),
    .io_enq_bits(q_509_io_enq_bits),
    .io_deq_ready(q_509_io_deq_ready),
    .io_deq_valid(q_509_io_deq_valid),
    .io_deq_bits(q_509_io_deq_bits)
  );
  Queue q_510 ( // @[Decoupled.scala 361:21]
    .clock(q_510_clock),
    .reset(q_510_reset),
    .io_enq_ready(q_510_io_enq_ready),
    .io_enq_valid(q_510_io_enq_valid),
    .io_enq_bits(q_510_io_enq_bits),
    .io_deq_ready(q_510_io_deq_ready),
    .io_deq_valid(q_510_io_deq_valid),
    .io_deq_bits(q_510_io_deq_bits)
  );
  Queue q_511 ( // @[Decoupled.scala 361:21]
    .clock(q_511_clock),
    .reset(q_511_reset),
    .io_enq_ready(q_511_io_enq_ready),
    .io_enq_valid(q_511_io_enq_valid),
    .io_enq_bits(q_511_io_enq_bits),
    .io_deq_ready(q_511_io_deq_ready),
    .io_deq_valid(q_511_io_deq_valid),
    .io_deq_bits(q_511_io_deq_bits)
  );
  Queue q_512 ( // @[Decoupled.scala 361:21]
    .clock(q_512_clock),
    .reset(q_512_reset),
    .io_enq_ready(q_512_io_enq_ready),
    .io_enq_valid(q_512_io_enq_valid),
    .io_enq_bits(q_512_io_enq_bits),
    .io_deq_ready(q_512_io_deq_ready),
    .io_deq_valid(q_512_io_deq_valid),
    .io_deq_bits(q_512_io_deq_bits)
  );
  Queue q_513 ( // @[Decoupled.scala 361:21]
    .clock(q_513_clock),
    .reset(q_513_reset),
    .io_enq_ready(q_513_io_enq_ready),
    .io_enq_valid(q_513_io_enq_valid),
    .io_enq_bits(q_513_io_enq_bits),
    .io_deq_ready(q_513_io_deq_ready),
    .io_deq_valid(q_513_io_deq_valid),
    .io_deq_bits(q_513_io_deq_bits)
  );
  Queue q_514 ( // @[Decoupled.scala 361:21]
    .clock(q_514_clock),
    .reset(q_514_reset),
    .io_enq_ready(q_514_io_enq_ready),
    .io_enq_valid(q_514_io_enq_valid),
    .io_enq_bits(q_514_io_enq_bits),
    .io_deq_ready(q_514_io_deq_ready),
    .io_deq_valid(q_514_io_deq_valid),
    .io_deq_bits(q_514_io_deq_bits)
  );
  Queue q_515 ( // @[Decoupled.scala 361:21]
    .clock(q_515_clock),
    .reset(q_515_reset),
    .io_enq_ready(q_515_io_enq_ready),
    .io_enq_valid(q_515_io_enq_valid),
    .io_enq_bits(q_515_io_enq_bits),
    .io_deq_ready(q_515_io_deq_ready),
    .io_deq_valid(q_515_io_deq_valid),
    .io_deq_bits(q_515_io_deq_bits)
  );
  Queue q_516 ( // @[Decoupled.scala 361:21]
    .clock(q_516_clock),
    .reset(q_516_reset),
    .io_enq_ready(q_516_io_enq_ready),
    .io_enq_valid(q_516_io_enq_valid),
    .io_enq_bits(q_516_io_enq_bits),
    .io_deq_ready(q_516_io_deq_ready),
    .io_deq_valid(q_516_io_deq_valid),
    .io_deq_bits(q_516_io_deq_bits)
  );
  Queue q_517 ( // @[Decoupled.scala 361:21]
    .clock(q_517_clock),
    .reset(q_517_reset),
    .io_enq_ready(q_517_io_enq_ready),
    .io_enq_valid(q_517_io_enq_valid),
    .io_enq_bits(q_517_io_enq_bits),
    .io_deq_ready(q_517_io_deq_ready),
    .io_deq_valid(q_517_io_deq_valid),
    .io_deq_bits(q_517_io_deq_bits)
  );
  Queue q_518 ( // @[Decoupled.scala 361:21]
    .clock(q_518_clock),
    .reset(q_518_reset),
    .io_enq_ready(q_518_io_enq_ready),
    .io_enq_valid(q_518_io_enq_valid),
    .io_enq_bits(q_518_io_enq_bits),
    .io_deq_ready(q_518_io_deq_ready),
    .io_deq_valid(q_518_io_deq_valid),
    .io_deq_bits(q_518_io_deq_bits)
  );
  Queue q_519 ( // @[Decoupled.scala 361:21]
    .clock(q_519_clock),
    .reset(q_519_reset),
    .io_enq_ready(q_519_io_enq_ready),
    .io_enq_valid(q_519_io_enq_valid),
    .io_enq_bits(q_519_io_enq_bits),
    .io_deq_ready(q_519_io_deq_ready),
    .io_deq_valid(q_519_io_deq_valid),
    .io_deq_bits(q_519_io_deq_bits)
  );
  Queue q_520 ( // @[Decoupled.scala 361:21]
    .clock(q_520_clock),
    .reset(q_520_reset),
    .io_enq_ready(q_520_io_enq_ready),
    .io_enq_valid(q_520_io_enq_valid),
    .io_enq_bits(q_520_io_enq_bits),
    .io_deq_ready(q_520_io_deq_ready),
    .io_deq_valid(q_520_io_deq_valid),
    .io_deq_bits(q_520_io_deq_bits)
  );
  Queue q_521 ( // @[Decoupled.scala 361:21]
    .clock(q_521_clock),
    .reset(q_521_reset),
    .io_enq_ready(q_521_io_enq_ready),
    .io_enq_valid(q_521_io_enq_valid),
    .io_enq_bits(q_521_io_enq_bits),
    .io_deq_ready(q_521_io_deq_ready),
    .io_deq_valid(q_521_io_deq_valid),
    .io_deq_bits(q_521_io_deq_bits)
  );
  Queue q_522 ( // @[Decoupled.scala 361:21]
    .clock(q_522_clock),
    .reset(q_522_reset),
    .io_enq_ready(q_522_io_enq_ready),
    .io_enq_valid(q_522_io_enq_valid),
    .io_enq_bits(q_522_io_enq_bits),
    .io_deq_ready(q_522_io_deq_ready),
    .io_deq_valid(q_522_io_deq_valid),
    .io_deq_bits(q_522_io_deq_bits)
  );
  Queue q_523 ( // @[Decoupled.scala 361:21]
    .clock(q_523_clock),
    .reset(q_523_reset),
    .io_enq_ready(q_523_io_enq_ready),
    .io_enq_valid(q_523_io_enq_valid),
    .io_enq_bits(q_523_io_enq_bits),
    .io_deq_ready(q_523_io_deq_ready),
    .io_deq_valid(q_523_io_deq_valid),
    .io_deq_bits(q_523_io_deq_bits)
  );
  Queue q_524 ( // @[Decoupled.scala 361:21]
    .clock(q_524_clock),
    .reset(q_524_reset),
    .io_enq_ready(q_524_io_enq_ready),
    .io_enq_valid(q_524_io_enq_valid),
    .io_enq_bits(q_524_io_enq_bits),
    .io_deq_ready(q_524_io_deq_ready),
    .io_deq_valid(q_524_io_deq_valid),
    .io_deq_bits(q_524_io_deq_bits)
  );
  Queue q_525 ( // @[Decoupled.scala 361:21]
    .clock(q_525_clock),
    .reset(q_525_reset),
    .io_enq_ready(q_525_io_enq_ready),
    .io_enq_valid(q_525_io_enq_valid),
    .io_enq_bits(q_525_io_enq_bits),
    .io_deq_ready(q_525_io_deq_ready),
    .io_deq_valid(q_525_io_deq_valid),
    .io_deq_bits(q_525_io_deq_bits)
  );
  Queue q_526 ( // @[Decoupled.scala 361:21]
    .clock(q_526_clock),
    .reset(q_526_reset),
    .io_enq_ready(q_526_io_enq_ready),
    .io_enq_valid(q_526_io_enq_valid),
    .io_enq_bits(q_526_io_enq_bits),
    .io_deq_ready(q_526_io_deq_ready),
    .io_deq_valid(q_526_io_deq_valid),
    .io_deq_bits(q_526_io_deq_bits)
  );
  Queue q_527 ( // @[Decoupled.scala 361:21]
    .clock(q_527_clock),
    .reset(q_527_reset),
    .io_enq_ready(q_527_io_enq_ready),
    .io_enq_valid(q_527_io_enq_valid),
    .io_enq_bits(q_527_io_enq_bits),
    .io_deq_ready(q_527_io_deq_ready),
    .io_deq_valid(q_527_io_deq_valid),
    .io_deq_bits(q_527_io_deq_bits)
  );
  Queue q_528 ( // @[Decoupled.scala 361:21]
    .clock(q_528_clock),
    .reset(q_528_reset),
    .io_enq_ready(q_528_io_enq_ready),
    .io_enq_valid(q_528_io_enq_valid),
    .io_enq_bits(q_528_io_enq_bits),
    .io_deq_ready(q_528_io_deq_ready),
    .io_deq_valid(q_528_io_deq_valid),
    .io_deq_bits(q_528_io_deq_bits)
  );
  Queue q_529 ( // @[Decoupled.scala 361:21]
    .clock(q_529_clock),
    .reset(q_529_reset),
    .io_enq_ready(q_529_io_enq_ready),
    .io_enq_valid(q_529_io_enq_valid),
    .io_enq_bits(q_529_io_enq_bits),
    .io_deq_ready(q_529_io_deq_ready),
    .io_deq_valid(q_529_io_deq_valid),
    .io_deq_bits(q_529_io_deq_bits)
  );
  Queue q_530 ( // @[Decoupled.scala 361:21]
    .clock(q_530_clock),
    .reset(q_530_reset),
    .io_enq_ready(q_530_io_enq_ready),
    .io_enq_valid(q_530_io_enq_valid),
    .io_enq_bits(q_530_io_enq_bits),
    .io_deq_ready(q_530_io_deq_ready),
    .io_deq_valid(q_530_io_deq_valid),
    .io_deq_bits(q_530_io_deq_bits)
  );
  Queue q_531 ( // @[Decoupled.scala 361:21]
    .clock(q_531_clock),
    .reset(q_531_reset),
    .io_enq_ready(q_531_io_enq_ready),
    .io_enq_valid(q_531_io_enq_valid),
    .io_enq_bits(q_531_io_enq_bits),
    .io_deq_ready(q_531_io_deq_ready),
    .io_deq_valid(q_531_io_deq_valid),
    .io_deq_bits(q_531_io_deq_bits)
  );
  Queue q_532 ( // @[Decoupled.scala 361:21]
    .clock(q_532_clock),
    .reset(q_532_reset),
    .io_enq_ready(q_532_io_enq_ready),
    .io_enq_valid(q_532_io_enq_valid),
    .io_enq_bits(q_532_io_enq_bits),
    .io_deq_ready(q_532_io_deq_ready),
    .io_deq_valid(q_532_io_deq_valid),
    .io_deq_bits(q_532_io_deq_bits)
  );
  Queue q_533 ( // @[Decoupled.scala 361:21]
    .clock(q_533_clock),
    .reset(q_533_reset),
    .io_enq_ready(q_533_io_enq_ready),
    .io_enq_valid(q_533_io_enq_valid),
    .io_enq_bits(q_533_io_enq_bits),
    .io_deq_ready(q_533_io_deq_ready),
    .io_deq_valid(q_533_io_deq_valid),
    .io_deq_bits(q_533_io_deq_bits)
  );
  Queue q_534 ( // @[Decoupled.scala 361:21]
    .clock(q_534_clock),
    .reset(q_534_reset),
    .io_enq_ready(q_534_io_enq_ready),
    .io_enq_valid(q_534_io_enq_valid),
    .io_enq_bits(q_534_io_enq_bits),
    .io_deq_ready(q_534_io_deq_ready),
    .io_deq_valid(q_534_io_deq_valid),
    .io_deq_bits(q_534_io_deq_bits)
  );
  Queue q_535 ( // @[Decoupled.scala 361:21]
    .clock(q_535_clock),
    .reset(q_535_reset),
    .io_enq_ready(q_535_io_enq_ready),
    .io_enq_valid(q_535_io_enq_valid),
    .io_enq_bits(q_535_io_enq_bits),
    .io_deq_ready(q_535_io_deq_ready),
    .io_deq_valid(q_535_io_deq_valid),
    .io_deq_bits(q_535_io_deq_bits)
  );
  Queue q_536 ( // @[Decoupled.scala 361:21]
    .clock(q_536_clock),
    .reset(q_536_reset),
    .io_enq_ready(q_536_io_enq_ready),
    .io_enq_valid(q_536_io_enq_valid),
    .io_enq_bits(q_536_io_enq_bits),
    .io_deq_ready(q_536_io_deq_ready),
    .io_deq_valid(q_536_io_deq_valid),
    .io_deq_bits(q_536_io_deq_bits)
  );
  Queue q_537 ( // @[Decoupled.scala 361:21]
    .clock(q_537_clock),
    .reset(q_537_reset),
    .io_enq_ready(q_537_io_enq_ready),
    .io_enq_valid(q_537_io_enq_valid),
    .io_enq_bits(q_537_io_enq_bits),
    .io_deq_ready(q_537_io_deq_ready),
    .io_deq_valid(q_537_io_deq_valid),
    .io_deq_bits(q_537_io_deq_bits)
  );
  Queue q_538 ( // @[Decoupled.scala 361:21]
    .clock(q_538_clock),
    .reset(q_538_reset),
    .io_enq_ready(q_538_io_enq_ready),
    .io_enq_valid(q_538_io_enq_valid),
    .io_enq_bits(q_538_io_enq_bits),
    .io_deq_ready(q_538_io_deq_ready),
    .io_deq_valid(q_538_io_deq_valid),
    .io_deq_bits(q_538_io_deq_bits)
  );
  Queue q_539 ( // @[Decoupled.scala 361:21]
    .clock(q_539_clock),
    .reset(q_539_reset),
    .io_enq_ready(q_539_io_enq_ready),
    .io_enq_valid(q_539_io_enq_valid),
    .io_enq_bits(q_539_io_enq_bits),
    .io_deq_ready(q_539_io_deq_ready),
    .io_deq_valid(q_539_io_deq_valid),
    .io_deq_bits(q_539_io_deq_bits)
  );
  Queue q_540 ( // @[Decoupled.scala 361:21]
    .clock(q_540_clock),
    .reset(q_540_reset),
    .io_enq_ready(q_540_io_enq_ready),
    .io_enq_valid(q_540_io_enq_valid),
    .io_enq_bits(q_540_io_enq_bits),
    .io_deq_ready(q_540_io_deq_ready),
    .io_deq_valid(q_540_io_deq_valid),
    .io_deq_bits(q_540_io_deq_bits)
  );
  Queue q_541 ( // @[Decoupled.scala 361:21]
    .clock(q_541_clock),
    .reset(q_541_reset),
    .io_enq_ready(q_541_io_enq_ready),
    .io_enq_valid(q_541_io_enq_valid),
    .io_enq_bits(q_541_io_enq_bits),
    .io_deq_ready(q_541_io_deq_ready),
    .io_deq_valid(q_541_io_deq_valid),
    .io_deq_bits(q_541_io_deq_bits)
  );
  Queue q_542 ( // @[Decoupled.scala 361:21]
    .clock(q_542_clock),
    .reset(q_542_reset),
    .io_enq_ready(q_542_io_enq_ready),
    .io_enq_valid(q_542_io_enq_valid),
    .io_enq_bits(q_542_io_enq_bits),
    .io_deq_ready(q_542_io_deq_ready),
    .io_deq_valid(q_542_io_deq_valid),
    .io_deq_bits(q_542_io_deq_bits)
  );
  Queue q_543 ( // @[Decoupled.scala 361:21]
    .clock(q_543_clock),
    .reset(q_543_reset),
    .io_enq_ready(q_543_io_enq_ready),
    .io_enq_valid(q_543_io_enq_valid),
    .io_enq_bits(q_543_io_enq_bits),
    .io_deq_ready(q_543_io_deq_ready),
    .io_deq_valid(q_543_io_deq_valid),
    .io_deq_bits(q_543_io_deq_bits)
  );
  Queue q_544 ( // @[Decoupled.scala 361:21]
    .clock(q_544_clock),
    .reset(q_544_reset),
    .io_enq_ready(q_544_io_enq_ready),
    .io_enq_valid(q_544_io_enq_valid),
    .io_enq_bits(q_544_io_enq_bits),
    .io_deq_ready(q_544_io_deq_ready),
    .io_deq_valid(q_544_io_deq_valid),
    .io_deq_bits(q_544_io_deq_bits)
  );
  Queue q_545 ( // @[Decoupled.scala 361:21]
    .clock(q_545_clock),
    .reset(q_545_reset),
    .io_enq_ready(q_545_io_enq_ready),
    .io_enq_valid(q_545_io_enq_valid),
    .io_enq_bits(q_545_io_enq_bits),
    .io_deq_ready(q_545_io_deq_ready),
    .io_deq_valid(q_545_io_deq_valid),
    .io_deq_bits(q_545_io_deq_bits)
  );
  Queue q_546 ( // @[Decoupled.scala 361:21]
    .clock(q_546_clock),
    .reset(q_546_reset),
    .io_enq_ready(q_546_io_enq_ready),
    .io_enq_valid(q_546_io_enq_valid),
    .io_enq_bits(q_546_io_enq_bits),
    .io_deq_ready(q_546_io_deq_ready),
    .io_deq_valid(q_546_io_deq_valid),
    .io_deq_bits(q_546_io_deq_bits)
  );
  Queue q_547 ( // @[Decoupled.scala 361:21]
    .clock(q_547_clock),
    .reset(q_547_reset),
    .io_enq_ready(q_547_io_enq_ready),
    .io_enq_valid(q_547_io_enq_valid),
    .io_enq_bits(q_547_io_enq_bits),
    .io_deq_ready(q_547_io_deq_ready),
    .io_deq_valid(q_547_io_deq_valid),
    .io_deq_bits(q_547_io_deq_bits)
  );
  Queue q_548 ( // @[Decoupled.scala 361:21]
    .clock(q_548_clock),
    .reset(q_548_reset),
    .io_enq_ready(q_548_io_enq_ready),
    .io_enq_valid(q_548_io_enq_valid),
    .io_enq_bits(q_548_io_enq_bits),
    .io_deq_ready(q_548_io_deq_ready),
    .io_deq_valid(q_548_io_deq_valid),
    .io_deq_bits(q_548_io_deq_bits)
  );
  Queue q_549 ( // @[Decoupled.scala 361:21]
    .clock(q_549_clock),
    .reset(q_549_reset),
    .io_enq_ready(q_549_io_enq_ready),
    .io_enq_valid(q_549_io_enq_valid),
    .io_enq_bits(q_549_io_enq_bits),
    .io_deq_ready(q_549_io_deq_ready),
    .io_deq_valid(q_549_io_deq_valid),
    .io_deq_bits(q_549_io_deq_bits)
  );
  Queue q_550 ( // @[Decoupled.scala 361:21]
    .clock(q_550_clock),
    .reset(q_550_reset),
    .io_enq_ready(q_550_io_enq_ready),
    .io_enq_valid(q_550_io_enq_valid),
    .io_enq_bits(q_550_io_enq_bits),
    .io_deq_ready(q_550_io_deq_ready),
    .io_deq_valid(q_550_io_deq_valid),
    .io_deq_bits(q_550_io_deq_bits)
  );
  Queue q_551 ( // @[Decoupled.scala 361:21]
    .clock(q_551_clock),
    .reset(q_551_reset),
    .io_enq_ready(q_551_io_enq_ready),
    .io_enq_valid(q_551_io_enq_valid),
    .io_enq_bits(q_551_io_enq_bits),
    .io_deq_ready(q_551_io_deq_ready),
    .io_deq_valid(q_551_io_deq_valid),
    .io_deq_bits(q_551_io_deq_bits)
  );
  Queue q_552 ( // @[Decoupled.scala 361:21]
    .clock(q_552_clock),
    .reset(q_552_reset),
    .io_enq_ready(q_552_io_enq_ready),
    .io_enq_valid(q_552_io_enq_valid),
    .io_enq_bits(q_552_io_enq_bits),
    .io_deq_ready(q_552_io_deq_ready),
    .io_deq_valid(q_552_io_deq_valid),
    .io_deq_bits(q_552_io_deq_bits)
  );
  Queue q_553 ( // @[Decoupled.scala 361:21]
    .clock(q_553_clock),
    .reset(q_553_reset),
    .io_enq_ready(q_553_io_enq_ready),
    .io_enq_valid(q_553_io_enq_valid),
    .io_enq_bits(q_553_io_enq_bits),
    .io_deq_ready(q_553_io_deq_ready),
    .io_deq_valid(q_553_io_deq_valid),
    .io_deq_bits(q_553_io_deq_bits)
  );
  Queue q_554 ( // @[Decoupled.scala 361:21]
    .clock(q_554_clock),
    .reset(q_554_reset),
    .io_enq_ready(q_554_io_enq_ready),
    .io_enq_valid(q_554_io_enq_valid),
    .io_enq_bits(q_554_io_enq_bits),
    .io_deq_ready(q_554_io_deq_ready),
    .io_deq_valid(q_554_io_deq_valid),
    .io_deq_bits(q_554_io_deq_bits)
  );
  Queue q_555 ( // @[Decoupled.scala 361:21]
    .clock(q_555_clock),
    .reset(q_555_reset),
    .io_enq_ready(q_555_io_enq_ready),
    .io_enq_valid(q_555_io_enq_valid),
    .io_enq_bits(q_555_io_enq_bits),
    .io_deq_ready(q_555_io_deq_ready),
    .io_deq_valid(q_555_io_deq_valid),
    .io_deq_bits(q_555_io_deq_bits)
  );
  Queue q_556 ( // @[Decoupled.scala 361:21]
    .clock(q_556_clock),
    .reset(q_556_reset),
    .io_enq_ready(q_556_io_enq_ready),
    .io_enq_valid(q_556_io_enq_valid),
    .io_enq_bits(q_556_io_enq_bits),
    .io_deq_ready(q_556_io_deq_ready),
    .io_deq_valid(q_556_io_deq_valid),
    .io_deq_bits(q_556_io_deq_bits)
  );
  Queue q_557 ( // @[Decoupled.scala 361:21]
    .clock(q_557_clock),
    .reset(q_557_reset),
    .io_enq_ready(q_557_io_enq_ready),
    .io_enq_valid(q_557_io_enq_valid),
    .io_enq_bits(q_557_io_enq_bits),
    .io_deq_ready(q_557_io_deq_ready),
    .io_deq_valid(q_557_io_deq_valid),
    .io_deq_bits(q_557_io_deq_bits)
  );
  Queue q_558 ( // @[Decoupled.scala 361:21]
    .clock(q_558_clock),
    .reset(q_558_reset),
    .io_enq_ready(q_558_io_enq_ready),
    .io_enq_valid(q_558_io_enq_valid),
    .io_enq_bits(q_558_io_enq_bits),
    .io_deq_ready(q_558_io_deq_ready),
    .io_deq_valid(q_558_io_deq_valid),
    .io_deq_bits(q_558_io_deq_bits)
  );
  Queue q_559 ( // @[Decoupled.scala 361:21]
    .clock(q_559_clock),
    .reset(q_559_reset),
    .io_enq_ready(q_559_io_enq_ready),
    .io_enq_valid(q_559_io_enq_valid),
    .io_enq_bits(q_559_io_enq_bits),
    .io_deq_ready(q_559_io_deq_ready),
    .io_deq_valid(q_559_io_deq_valid),
    .io_deq_bits(q_559_io_deq_bits)
  );
  Queue q_560 ( // @[Decoupled.scala 361:21]
    .clock(q_560_clock),
    .reset(q_560_reset),
    .io_enq_ready(q_560_io_enq_ready),
    .io_enq_valid(q_560_io_enq_valid),
    .io_enq_bits(q_560_io_enq_bits),
    .io_deq_ready(q_560_io_deq_ready),
    .io_deq_valid(q_560_io_deq_valid),
    .io_deq_bits(q_560_io_deq_bits)
  );
  Queue q_561 ( // @[Decoupled.scala 361:21]
    .clock(q_561_clock),
    .reset(q_561_reset),
    .io_enq_ready(q_561_io_enq_ready),
    .io_enq_valid(q_561_io_enq_valid),
    .io_enq_bits(q_561_io_enq_bits),
    .io_deq_ready(q_561_io_deq_ready),
    .io_deq_valid(q_561_io_deq_valid),
    .io_deq_bits(q_561_io_deq_bits)
  );
  Queue q_562 ( // @[Decoupled.scala 361:21]
    .clock(q_562_clock),
    .reset(q_562_reset),
    .io_enq_ready(q_562_io_enq_ready),
    .io_enq_valid(q_562_io_enq_valid),
    .io_enq_bits(q_562_io_enq_bits),
    .io_deq_ready(q_562_io_deq_ready),
    .io_deq_valid(q_562_io_deq_valid),
    .io_deq_bits(q_562_io_deq_bits)
  );
  Queue q_563 ( // @[Decoupled.scala 361:21]
    .clock(q_563_clock),
    .reset(q_563_reset),
    .io_enq_ready(q_563_io_enq_ready),
    .io_enq_valid(q_563_io_enq_valid),
    .io_enq_bits(q_563_io_enq_bits),
    .io_deq_ready(q_563_io_deq_ready),
    .io_deq_valid(q_563_io_deq_valid),
    .io_deq_bits(q_563_io_deq_bits)
  );
  Queue q_564 ( // @[Decoupled.scala 361:21]
    .clock(q_564_clock),
    .reset(q_564_reset),
    .io_enq_ready(q_564_io_enq_ready),
    .io_enq_valid(q_564_io_enq_valid),
    .io_enq_bits(q_564_io_enq_bits),
    .io_deq_ready(q_564_io_deq_ready),
    .io_deq_valid(q_564_io_deq_valid),
    .io_deq_bits(q_564_io_deq_bits)
  );
  Queue q_565 ( // @[Decoupled.scala 361:21]
    .clock(q_565_clock),
    .reset(q_565_reset),
    .io_enq_ready(q_565_io_enq_ready),
    .io_enq_valid(q_565_io_enq_valid),
    .io_enq_bits(q_565_io_enq_bits),
    .io_deq_ready(q_565_io_deq_ready),
    .io_deq_valid(q_565_io_deq_valid),
    .io_deq_bits(q_565_io_deq_bits)
  );
  Queue q_566 ( // @[Decoupled.scala 361:21]
    .clock(q_566_clock),
    .reset(q_566_reset),
    .io_enq_ready(q_566_io_enq_ready),
    .io_enq_valid(q_566_io_enq_valid),
    .io_enq_bits(q_566_io_enq_bits),
    .io_deq_ready(q_566_io_deq_ready),
    .io_deq_valid(q_566_io_deq_valid),
    .io_deq_bits(q_566_io_deq_bits)
  );
  Queue q_567 ( // @[Decoupled.scala 361:21]
    .clock(q_567_clock),
    .reset(q_567_reset),
    .io_enq_ready(q_567_io_enq_ready),
    .io_enq_valid(q_567_io_enq_valid),
    .io_enq_bits(q_567_io_enq_bits),
    .io_deq_ready(q_567_io_deq_ready),
    .io_deq_valid(q_567_io_deq_valid),
    .io_deq_bits(q_567_io_deq_bits)
  );
  Queue q_568 ( // @[Decoupled.scala 361:21]
    .clock(q_568_clock),
    .reset(q_568_reset),
    .io_enq_ready(q_568_io_enq_ready),
    .io_enq_valid(q_568_io_enq_valid),
    .io_enq_bits(q_568_io_enq_bits),
    .io_deq_ready(q_568_io_deq_ready),
    .io_deq_valid(q_568_io_deq_valid),
    .io_deq_bits(q_568_io_deq_bits)
  );
  Queue q_569 ( // @[Decoupled.scala 361:21]
    .clock(q_569_clock),
    .reset(q_569_reset),
    .io_enq_ready(q_569_io_enq_ready),
    .io_enq_valid(q_569_io_enq_valid),
    .io_enq_bits(q_569_io_enq_bits),
    .io_deq_ready(q_569_io_deq_ready),
    .io_deq_valid(q_569_io_deq_valid),
    .io_deq_bits(q_569_io_deq_bits)
  );
  Queue q_570 ( // @[Decoupled.scala 361:21]
    .clock(q_570_clock),
    .reset(q_570_reset),
    .io_enq_ready(q_570_io_enq_ready),
    .io_enq_valid(q_570_io_enq_valid),
    .io_enq_bits(q_570_io_enq_bits),
    .io_deq_ready(q_570_io_deq_ready),
    .io_deq_valid(q_570_io_deq_valid),
    .io_deq_bits(q_570_io_deq_bits)
  );
  Queue q_571 ( // @[Decoupled.scala 361:21]
    .clock(q_571_clock),
    .reset(q_571_reset),
    .io_enq_ready(q_571_io_enq_ready),
    .io_enq_valid(q_571_io_enq_valid),
    .io_enq_bits(q_571_io_enq_bits),
    .io_deq_ready(q_571_io_deq_ready),
    .io_deq_valid(q_571_io_deq_valid),
    .io_deq_bits(q_571_io_deq_bits)
  );
  Queue q_572 ( // @[Decoupled.scala 361:21]
    .clock(q_572_clock),
    .reset(q_572_reset),
    .io_enq_ready(q_572_io_enq_ready),
    .io_enq_valid(q_572_io_enq_valid),
    .io_enq_bits(q_572_io_enq_bits),
    .io_deq_ready(q_572_io_deq_ready),
    .io_deq_valid(q_572_io_deq_valid),
    .io_deq_bits(q_572_io_deq_bits)
  );
  Queue q_573 ( // @[Decoupled.scala 361:21]
    .clock(q_573_clock),
    .reset(q_573_reset),
    .io_enq_ready(q_573_io_enq_ready),
    .io_enq_valid(q_573_io_enq_valid),
    .io_enq_bits(q_573_io_enq_bits),
    .io_deq_ready(q_573_io_deq_ready),
    .io_deq_valid(q_573_io_deq_valid),
    .io_deq_bits(q_573_io_deq_bits)
  );
  Queue q_574 ( // @[Decoupled.scala 361:21]
    .clock(q_574_clock),
    .reset(q_574_reset),
    .io_enq_ready(q_574_io_enq_ready),
    .io_enq_valid(q_574_io_enq_valid),
    .io_enq_bits(q_574_io_enq_bits),
    .io_deq_ready(q_574_io_deq_ready),
    .io_deq_valid(q_574_io_deq_valid),
    .io_deq_bits(q_574_io_deq_bits)
  );
  Queue q_575 ( // @[Decoupled.scala 361:21]
    .clock(q_575_clock),
    .reset(q_575_reset),
    .io_enq_ready(q_575_io_enq_ready),
    .io_enq_valid(q_575_io_enq_valid),
    .io_enq_bits(q_575_io_enq_bits),
    .io_deq_ready(q_575_io_deq_ready),
    .io_deq_valid(q_575_io_deq_valid),
    .io_deq_bits(q_575_io_deq_bits)
  );
  Queue q_576 ( // @[Decoupled.scala 361:21]
    .clock(q_576_clock),
    .reset(q_576_reset),
    .io_enq_ready(q_576_io_enq_ready),
    .io_enq_valid(q_576_io_enq_valid),
    .io_enq_bits(q_576_io_enq_bits),
    .io_deq_ready(q_576_io_deq_ready),
    .io_deq_valid(q_576_io_deq_valid),
    .io_deq_bits(q_576_io_deq_bits)
  );
  Queue q_577 ( // @[Decoupled.scala 361:21]
    .clock(q_577_clock),
    .reset(q_577_reset),
    .io_enq_ready(q_577_io_enq_ready),
    .io_enq_valid(q_577_io_enq_valid),
    .io_enq_bits(q_577_io_enq_bits),
    .io_deq_ready(q_577_io_deq_ready),
    .io_deq_valid(q_577_io_deq_valid),
    .io_deq_bits(q_577_io_deq_bits)
  );
  Queue q_578 ( // @[Decoupled.scala 361:21]
    .clock(q_578_clock),
    .reset(q_578_reset),
    .io_enq_ready(q_578_io_enq_ready),
    .io_enq_valid(q_578_io_enq_valid),
    .io_enq_bits(q_578_io_enq_bits),
    .io_deq_ready(q_578_io_deq_ready),
    .io_deq_valid(q_578_io_deq_valid),
    .io_deq_bits(q_578_io_deq_bits)
  );
  Queue q_579 ( // @[Decoupled.scala 361:21]
    .clock(q_579_clock),
    .reset(q_579_reset),
    .io_enq_ready(q_579_io_enq_ready),
    .io_enq_valid(q_579_io_enq_valid),
    .io_enq_bits(q_579_io_enq_bits),
    .io_deq_ready(q_579_io_deq_ready),
    .io_deq_valid(q_579_io_deq_valid),
    .io_deq_bits(q_579_io_deq_bits)
  );
  Queue q_580 ( // @[Decoupled.scala 361:21]
    .clock(q_580_clock),
    .reset(q_580_reset),
    .io_enq_ready(q_580_io_enq_ready),
    .io_enq_valid(q_580_io_enq_valid),
    .io_enq_bits(q_580_io_enq_bits),
    .io_deq_ready(q_580_io_deq_ready),
    .io_deq_valid(q_580_io_deq_valid),
    .io_deq_bits(q_580_io_deq_bits)
  );
  Queue q_581 ( // @[Decoupled.scala 361:21]
    .clock(q_581_clock),
    .reset(q_581_reset),
    .io_enq_ready(q_581_io_enq_ready),
    .io_enq_valid(q_581_io_enq_valid),
    .io_enq_bits(q_581_io_enq_bits),
    .io_deq_ready(q_581_io_deq_ready),
    .io_deq_valid(q_581_io_deq_valid),
    .io_deq_bits(q_581_io_deq_bits)
  );
  Queue q_582 ( // @[Decoupled.scala 361:21]
    .clock(q_582_clock),
    .reset(q_582_reset),
    .io_enq_ready(q_582_io_enq_ready),
    .io_enq_valid(q_582_io_enq_valid),
    .io_enq_bits(q_582_io_enq_bits),
    .io_deq_ready(q_582_io_deq_ready),
    .io_deq_valid(q_582_io_deq_valid),
    .io_deq_bits(q_582_io_deq_bits)
  );
  Queue q_583 ( // @[Decoupled.scala 361:21]
    .clock(q_583_clock),
    .reset(q_583_reset),
    .io_enq_ready(q_583_io_enq_ready),
    .io_enq_valid(q_583_io_enq_valid),
    .io_enq_bits(q_583_io_enq_bits),
    .io_deq_ready(q_583_io_deq_ready),
    .io_deq_valid(q_583_io_deq_valid),
    .io_deq_bits(q_583_io_deq_bits)
  );
  Queue q_584 ( // @[Decoupled.scala 361:21]
    .clock(q_584_clock),
    .reset(q_584_reset),
    .io_enq_ready(q_584_io_enq_ready),
    .io_enq_valid(q_584_io_enq_valid),
    .io_enq_bits(q_584_io_enq_bits),
    .io_deq_ready(q_584_io_deq_ready),
    .io_deq_valid(q_584_io_deq_valid),
    .io_deq_bits(q_584_io_deq_bits)
  );
  Queue q_585 ( // @[Decoupled.scala 361:21]
    .clock(q_585_clock),
    .reset(q_585_reset),
    .io_enq_ready(q_585_io_enq_ready),
    .io_enq_valid(q_585_io_enq_valid),
    .io_enq_bits(q_585_io_enq_bits),
    .io_deq_ready(q_585_io_deq_ready),
    .io_deq_valid(q_585_io_deq_valid),
    .io_deq_bits(q_585_io_deq_bits)
  );
  Queue q_586 ( // @[Decoupled.scala 361:21]
    .clock(q_586_clock),
    .reset(q_586_reset),
    .io_enq_ready(q_586_io_enq_ready),
    .io_enq_valid(q_586_io_enq_valid),
    .io_enq_bits(q_586_io_enq_bits),
    .io_deq_ready(q_586_io_deq_ready),
    .io_deq_valid(q_586_io_deq_valid),
    .io_deq_bits(q_586_io_deq_bits)
  );
  Queue q_587 ( // @[Decoupled.scala 361:21]
    .clock(q_587_clock),
    .reset(q_587_reset),
    .io_enq_ready(q_587_io_enq_ready),
    .io_enq_valid(q_587_io_enq_valid),
    .io_enq_bits(q_587_io_enq_bits),
    .io_deq_ready(q_587_io_deq_ready),
    .io_deq_valid(q_587_io_deq_valid),
    .io_deq_bits(q_587_io_deq_bits)
  );
  Queue q_588 ( // @[Decoupled.scala 361:21]
    .clock(q_588_clock),
    .reset(q_588_reset),
    .io_enq_ready(q_588_io_enq_ready),
    .io_enq_valid(q_588_io_enq_valid),
    .io_enq_bits(q_588_io_enq_bits),
    .io_deq_ready(q_588_io_deq_ready),
    .io_deq_valid(q_588_io_deq_valid),
    .io_deq_bits(q_588_io_deq_bits)
  );
  Queue q_589 ( // @[Decoupled.scala 361:21]
    .clock(q_589_clock),
    .reset(q_589_reset),
    .io_enq_ready(q_589_io_enq_ready),
    .io_enq_valid(q_589_io_enq_valid),
    .io_enq_bits(q_589_io_enq_bits),
    .io_deq_ready(q_589_io_deq_ready),
    .io_deq_valid(q_589_io_deq_valid),
    .io_deq_bits(q_589_io_deq_bits)
  );
  Queue q_590 ( // @[Decoupled.scala 361:21]
    .clock(q_590_clock),
    .reset(q_590_reset),
    .io_enq_ready(q_590_io_enq_ready),
    .io_enq_valid(q_590_io_enq_valid),
    .io_enq_bits(q_590_io_enq_bits),
    .io_deq_ready(q_590_io_deq_ready),
    .io_deq_valid(q_590_io_deq_valid),
    .io_deq_bits(q_590_io_deq_bits)
  );
  Queue q_591 ( // @[Decoupled.scala 361:21]
    .clock(q_591_clock),
    .reset(q_591_reset),
    .io_enq_ready(q_591_io_enq_ready),
    .io_enq_valid(q_591_io_enq_valid),
    .io_enq_bits(q_591_io_enq_bits),
    .io_deq_ready(q_591_io_deq_ready),
    .io_deq_valid(q_591_io_deq_valid),
    .io_deq_bits(q_591_io_deq_bits)
  );
  Queue q_592 ( // @[Decoupled.scala 361:21]
    .clock(q_592_clock),
    .reset(q_592_reset),
    .io_enq_ready(q_592_io_enq_ready),
    .io_enq_valid(q_592_io_enq_valid),
    .io_enq_bits(q_592_io_enq_bits),
    .io_deq_ready(q_592_io_deq_ready),
    .io_deq_valid(q_592_io_deq_valid),
    .io_deq_bits(q_592_io_deq_bits)
  );
  Queue q_593 ( // @[Decoupled.scala 361:21]
    .clock(q_593_clock),
    .reset(q_593_reset),
    .io_enq_ready(q_593_io_enq_ready),
    .io_enq_valid(q_593_io_enq_valid),
    .io_enq_bits(q_593_io_enq_bits),
    .io_deq_ready(q_593_io_deq_ready),
    .io_deq_valid(q_593_io_deq_valid),
    .io_deq_bits(q_593_io_deq_bits)
  );
  Queue q_594 ( // @[Decoupled.scala 361:21]
    .clock(q_594_clock),
    .reset(q_594_reset),
    .io_enq_ready(q_594_io_enq_ready),
    .io_enq_valid(q_594_io_enq_valid),
    .io_enq_bits(q_594_io_enq_bits),
    .io_deq_ready(q_594_io_deq_ready),
    .io_deq_valid(q_594_io_deq_valid),
    .io_deq_bits(q_594_io_deq_bits)
  );
  Queue q_595 ( // @[Decoupled.scala 361:21]
    .clock(q_595_clock),
    .reset(q_595_reset),
    .io_enq_ready(q_595_io_enq_ready),
    .io_enq_valid(q_595_io_enq_valid),
    .io_enq_bits(q_595_io_enq_bits),
    .io_deq_ready(q_595_io_deq_ready),
    .io_deq_valid(q_595_io_deq_valid),
    .io_deq_bits(q_595_io_deq_bits)
  );
  Queue q_596 ( // @[Decoupled.scala 361:21]
    .clock(q_596_clock),
    .reset(q_596_reset),
    .io_enq_ready(q_596_io_enq_ready),
    .io_enq_valid(q_596_io_enq_valid),
    .io_enq_bits(q_596_io_enq_bits),
    .io_deq_ready(q_596_io_deq_ready),
    .io_deq_valid(q_596_io_deq_valid),
    .io_deq_bits(q_596_io_deq_bits)
  );
  Queue q_597 ( // @[Decoupled.scala 361:21]
    .clock(q_597_clock),
    .reset(q_597_reset),
    .io_enq_ready(q_597_io_enq_ready),
    .io_enq_valid(q_597_io_enq_valid),
    .io_enq_bits(q_597_io_enq_bits),
    .io_deq_ready(q_597_io_deq_ready),
    .io_deq_valid(q_597_io_deq_valid),
    .io_deq_bits(q_597_io_deq_bits)
  );
  Queue q_598 ( // @[Decoupled.scala 361:21]
    .clock(q_598_clock),
    .reset(q_598_reset),
    .io_enq_ready(q_598_io_enq_ready),
    .io_enq_valid(q_598_io_enq_valid),
    .io_enq_bits(q_598_io_enq_bits),
    .io_deq_ready(q_598_io_deq_ready),
    .io_deq_valid(q_598_io_deq_valid),
    .io_deq_bits(q_598_io_deq_bits)
  );
  Queue q_599 ( // @[Decoupled.scala 361:21]
    .clock(q_599_clock),
    .reset(q_599_reset),
    .io_enq_ready(q_599_io_enq_ready),
    .io_enq_valid(q_599_io_enq_valid),
    .io_enq_bits(q_599_io_enq_bits),
    .io_deq_ready(q_599_io_deq_ready),
    .io_deq_valid(q_599_io_deq_valid),
    .io_deq_bits(q_599_io_deq_bits)
  );
  Queue q_600 ( // @[Decoupled.scala 361:21]
    .clock(q_600_clock),
    .reset(q_600_reset),
    .io_enq_ready(q_600_io_enq_ready),
    .io_enq_valid(q_600_io_enq_valid),
    .io_enq_bits(q_600_io_enq_bits),
    .io_deq_ready(q_600_io_deq_ready),
    .io_deq_valid(q_600_io_deq_valid),
    .io_deq_bits(q_600_io_deq_bits)
  );
  Queue q_601 ( // @[Decoupled.scala 361:21]
    .clock(q_601_clock),
    .reset(q_601_reset),
    .io_enq_ready(q_601_io_enq_ready),
    .io_enq_valid(q_601_io_enq_valid),
    .io_enq_bits(q_601_io_enq_bits),
    .io_deq_ready(q_601_io_deq_ready),
    .io_deq_valid(q_601_io_deq_valid),
    .io_deq_bits(q_601_io_deq_bits)
  );
  Queue q_602 ( // @[Decoupled.scala 361:21]
    .clock(q_602_clock),
    .reset(q_602_reset),
    .io_enq_ready(q_602_io_enq_ready),
    .io_enq_valid(q_602_io_enq_valid),
    .io_enq_bits(q_602_io_enq_bits),
    .io_deq_ready(q_602_io_deq_ready),
    .io_deq_valid(q_602_io_deq_valid),
    .io_deq_bits(q_602_io_deq_bits)
  );
  Queue q_603 ( // @[Decoupled.scala 361:21]
    .clock(q_603_clock),
    .reset(q_603_reset),
    .io_enq_ready(q_603_io_enq_ready),
    .io_enq_valid(q_603_io_enq_valid),
    .io_enq_bits(q_603_io_enq_bits),
    .io_deq_ready(q_603_io_deq_ready),
    .io_deq_valid(q_603_io_deq_valid),
    .io_deq_bits(q_603_io_deq_bits)
  );
  Queue q_604 ( // @[Decoupled.scala 361:21]
    .clock(q_604_clock),
    .reset(q_604_reset),
    .io_enq_ready(q_604_io_enq_ready),
    .io_enq_valid(q_604_io_enq_valid),
    .io_enq_bits(q_604_io_enq_bits),
    .io_deq_ready(q_604_io_deq_ready),
    .io_deq_valid(q_604_io_deq_valid),
    .io_deq_bits(q_604_io_deq_bits)
  );
  Queue q_605 ( // @[Decoupled.scala 361:21]
    .clock(q_605_clock),
    .reset(q_605_reset),
    .io_enq_ready(q_605_io_enq_ready),
    .io_enq_valid(q_605_io_enq_valid),
    .io_enq_bits(q_605_io_enq_bits),
    .io_deq_ready(q_605_io_deq_ready),
    .io_deq_valid(q_605_io_deq_valid),
    .io_deq_bits(q_605_io_deq_bits)
  );
  Queue q_606 ( // @[Decoupled.scala 361:21]
    .clock(q_606_clock),
    .reset(q_606_reset),
    .io_enq_ready(q_606_io_enq_ready),
    .io_enq_valid(q_606_io_enq_valid),
    .io_enq_bits(q_606_io_enq_bits),
    .io_deq_ready(q_606_io_deq_ready),
    .io_deq_valid(q_606_io_deq_valid),
    .io_deq_bits(q_606_io_deq_bits)
  );
  Queue q_607 ( // @[Decoupled.scala 361:21]
    .clock(q_607_clock),
    .reset(q_607_reset),
    .io_enq_ready(q_607_io_enq_ready),
    .io_enq_valid(q_607_io_enq_valid),
    .io_enq_bits(q_607_io_enq_bits),
    .io_deq_ready(q_607_io_deq_ready),
    .io_deq_valid(q_607_io_deq_valid),
    .io_deq_bits(q_607_io_deq_bits)
  );
  Queue q_608 ( // @[Decoupled.scala 361:21]
    .clock(q_608_clock),
    .reset(q_608_reset),
    .io_enq_ready(q_608_io_enq_ready),
    .io_enq_valid(q_608_io_enq_valid),
    .io_enq_bits(q_608_io_enq_bits),
    .io_deq_ready(q_608_io_deq_ready),
    .io_deq_valid(q_608_io_deq_valid),
    .io_deq_bits(q_608_io_deq_bits)
  );
  Queue q_609 ( // @[Decoupled.scala 361:21]
    .clock(q_609_clock),
    .reset(q_609_reset),
    .io_enq_ready(q_609_io_enq_ready),
    .io_enq_valid(q_609_io_enq_valid),
    .io_enq_bits(q_609_io_enq_bits),
    .io_deq_ready(q_609_io_deq_ready),
    .io_deq_valid(q_609_io_deq_valid),
    .io_deq_bits(q_609_io_deq_bits)
  );
  Queue q_610 ( // @[Decoupled.scala 361:21]
    .clock(q_610_clock),
    .reset(q_610_reset),
    .io_enq_ready(q_610_io_enq_ready),
    .io_enq_valid(q_610_io_enq_valid),
    .io_enq_bits(q_610_io_enq_bits),
    .io_deq_ready(q_610_io_deq_ready),
    .io_deq_valid(q_610_io_deq_valid),
    .io_deq_bits(q_610_io_deq_bits)
  );
  Queue q_611 ( // @[Decoupled.scala 361:21]
    .clock(q_611_clock),
    .reset(q_611_reset),
    .io_enq_ready(q_611_io_enq_ready),
    .io_enq_valid(q_611_io_enq_valid),
    .io_enq_bits(q_611_io_enq_bits),
    .io_deq_ready(q_611_io_deq_ready),
    .io_deq_valid(q_611_io_deq_valid),
    .io_deq_bits(q_611_io_deq_bits)
  );
  Queue q_612 ( // @[Decoupled.scala 361:21]
    .clock(q_612_clock),
    .reset(q_612_reset),
    .io_enq_ready(q_612_io_enq_ready),
    .io_enq_valid(q_612_io_enq_valid),
    .io_enq_bits(q_612_io_enq_bits),
    .io_deq_ready(q_612_io_deq_ready),
    .io_deq_valid(q_612_io_deq_valid),
    .io_deq_bits(q_612_io_deq_bits)
  );
  Queue q_613 ( // @[Decoupled.scala 361:21]
    .clock(q_613_clock),
    .reset(q_613_reset),
    .io_enq_ready(q_613_io_enq_ready),
    .io_enq_valid(q_613_io_enq_valid),
    .io_enq_bits(q_613_io_enq_bits),
    .io_deq_ready(q_613_io_deq_ready),
    .io_deq_valid(q_613_io_deq_valid),
    .io_deq_bits(q_613_io_deq_bits)
  );
  Queue q_614 ( // @[Decoupled.scala 361:21]
    .clock(q_614_clock),
    .reset(q_614_reset),
    .io_enq_ready(q_614_io_enq_ready),
    .io_enq_valid(q_614_io_enq_valid),
    .io_enq_bits(q_614_io_enq_bits),
    .io_deq_ready(q_614_io_deq_ready),
    .io_deq_valid(q_614_io_deq_valid),
    .io_deq_bits(q_614_io_deq_bits)
  );
  Queue q_615 ( // @[Decoupled.scala 361:21]
    .clock(q_615_clock),
    .reset(q_615_reset),
    .io_enq_ready(q_615_io_enq_ready),
    .io_enq_valid(q_615_io_enq_valid),
    .io_enq_bits(q_615_io_enq_bits),
    .io_deq_ready(q_615_io_deq_ready),
    .io_deq_valid(q_615_io_deq_valid),
    .io_deq_bits(q_615_io_deq_bits)
  );
  Queue q_616 ( // @[Decoupled.scala 361:21]
    .clock(q_616_clock),
    .reset(q_616_reset),
    .io_enq_ready(q_616_io_enq_ready),
    .io_enq_valid(q_616_io_enq_valid),
    .io_enq_bits(q_616_io_enq_bits),
    .io_deq_ready(q_616_io_deq_ready),
    .io_deq_valid(q_616_io_deq_valid),
    .io_deq_bits(q_616_io_deq_bits)
  );
  Queue q_617 ( // @[Decoupled.scala 361:21]
    .clock(q_617_clock),
    .reset(q_617_reset),
    .io_enq_ready(q_617_io_enq_ready),
    .io_enq_valid(q_617_io_enq_valid),
    .io_enq_bits(q_617_io_enq_bits),
    .io_deq_ready(q_617_io_deq_ready),
    .io_deq_valid(q_617_io_deq_valid),
    .io_deq_bits(q_617_io_deq_bits)
  );
  Queue q_618 ( // @[Decoupled.scala 361:21]
    .clock(q_618_clock),
    .reset(q_618_reset),
    .io_enq_ready(q_618_io_enq_ready),
    .io_enq_valid(q_618_io_enq_valid),
    .io_enq_bits(q_618_io_enq_bits),
    .io_deq_ready(q_618_io_deq_ready),
    .io_deq_valid(q_618_io_deq_valid),
    .io_deq_bits(q_618_io_deq_bits)
  );
  Queue q_619 ( // @[Decoupled.scala 361:21]
    .clock(q_619_clock),
    .reset(q_619_reset),
    .io_enq_ready(q_619_io_enq_ready),
    .io_enq_valid(q_619_io_enq_valid),
    .io_enq_bits(q_619_io_enq_bits),
    .io_deq_ready(q_619_io_deq_ready),
    .io_deq_valid(q_619_io_deq_valid),
    .io_deq_bits(q_619_io_deq_bits)
  );
  Queue q_620 ( // @[Decoupled.scala 361:21]
    .clock(q_620_clock),
    .reset(q_620_reset),
    .io_enq_ready(q_620_io_enq_ready),
    .io_enq_valid(q_620_io_enq_valid),
    .io_enq_bits(q_620_io_enq_bits),
    .io_deq_ready(q_620_io_deq_ready),
    .io_deq_valid(q_620_io_deq_valid),
    .io_deq_bits(q_620_io_deq_bits)
  );
  Queue q_621 ( // @[Decoupled.scala 361:21]
    .clock(q_621_clock),
    .reset(q_621_reset),
    .io_enq_ready(q_621_io_enq_ready),
    .io_enq_valid(q_621_io_enq_valid),
    .io_enq_bits(q_621_io_enq_bits),
    .io_deq_ready(q_621_io_deq_ready),
    .io_deq_valid(q_621_io_deq_valid),
    .io_deq_bits(q_621_io_deq_bits)
  );
  Queue q_622 ( // @[Decoupled.scala 361:21]
    .clock(q_622_clock),
    .reset(q_622_reset),
    .io_enq_ready(q_622_io_enq_ready),
    .io_enq_valid(q_622_io_enq_valid),
    .io_enq_bits(q_622_io_enq_bits),
    .io_deq_ready(q_622_io_deq_ready),
    .io_deq_valid(q_622_io_deq_valid),
    .io_deq_bits(q_622_io_deq_bits)
  );
  Queue q_623 ( // @[Decoupled.scala 361:21]
    .clock(q_623_clock),
    .reset(q_623_reset),
    .io_enq_ready(q_623_io_enq_ready),
    .io_enq_valid(q_623_io_enq_valid),
    .io_enq_bits(q_623_io_enq_bits),
    .io_deq_ready(q_623_io_deq_ready),
    .io_deq_valid(q_623_io_deq_valid),
    .io_deq_bits(q_623_io_deq_bits)
  );
  Queue q_624 ( // @[Decoupled.scala 361:21]
    .clock(q_624_clock),
    .reset(q_624_reset),
    .io_enq_ready(q_624_io_enq_ready),
    .io_enq_valid(q_624_io_enq_valid),
    .io_enq_bits(q_624_io_enq_bits),
    .io_deq_ready(q_624_io_deq_ready),
    .io_deq_valid(q_624_io_deq_valid),
    .io_deq_bits(q_624_io_deq_bits)
  );
  Queue q_625 ( // @[Decoupled.scala 361:21]
    .clock(q_625_clock),
    .reset(q_625_reset),
    .io_enq_ready(q_625_io_enq_ready),
    .io_enq_valid(q_625_io_enq_valid),
    .io_enq_bits(q_625_io_enq_bits),
    .io_deq_ready(q_625_io_deq_ready),
    .io_deq_valid(q_625_io_deq_valid),
    .io_deq_bits(q_625_io_deq_bits)
  );
  Queue q_626 ( // @[Decoupled.scala 361:21]
    .clock(q_626_clock),
    .reset(q_626_reset),
    .io_enq_ready(q_626_io_enq_ready),
    .io_enq_valid(q_626_io_enq_valid),
    .io_enq_bits(q_626_io_enq_bits),
    .io_deq_ready(q_626_io_deq_ready),
    .io_deq_valid(q_626_io_deq_valid),
    .io_deq_bits(q_626_io_deq_bits)
  );
  Queue q_627 ( // @[Decoupled.scala 361:21]
    .clock(q_627_clock),
    .reset(q_627_reset),
    .io_enq_ready(q_627_io_enq_ready),
    .io_enq_valid(q_627_io_enq_valid),
    .io_enq_bits(q_627_io_enq_bits),
    .io_deq_ready(q_627_io_deq_ready),
    .io_deq_valid(q_627_io_deq_valid),
    .io_deq_bits(q_627_io_deq_bits)
  );
  Queue q_628 ( // @[Decoupled.scala 361:21]
    .clock(q_628_clock),
    .reset(q_628_reset),
    .io_enq_ready(q_628_io_enq_ready),
    .io_enq_valid(q_628_io_enq_valid),
    .io_enq_bits(q_628_io_enq_bits),
    .io_deq_ready(q_628_io_deq_ready),
    .io_deq_valid(q_628_io_deq_valid),
    .io_deq_bits(q_628_io_deq_bits)
  );
  Queue q_629 ( // @[Decoupled.scala 361:21]
    .clock(q_629_clock),
    .reset(q_629_reset),
    .io_enq_ready(q_629_io_enq_ready),
    .io_enq_valid(q_629_io_enq_valid),
    .io_enq_bits(q_629_io_enq_bits),
    .io_deq_ready(q_629_io_deq_ready),
    .io_deq_valid(q_629_io_deq_valid),
    .io_deq_bits(q_629_io_deq_bits)
  );
  Queue q_630 ( // @[Decoupled.scala 361:21]
    .clock(q_630_clock),
    .reset(q_630_reset),
    .io_enq_ready(q_630_io_enq_ready),
    .io_enq_valid(q_630_io_enq_valid),
    .io_enq_bits(q_630_io_enq_bits),
    .io_deq_ready(q_630_io_deq_ready),
    .io_deq_valid(q_630_io_deq_valid),
    .io_deq_bits(q_630_io_deq_bits)
  );
  Queue q_631 ( // @[Decoupled.scala 361:21]
    .clock(q_631_clock),
    .reset(q_631_reset),
    .io_enq_ready(q_631_io_enq_ready),
    .io_enq_valid(q_631_io_enq_valid),
    .io_enq_bits(q_631_io_enq_bits),
    .io_deq_ready(q_631_io_deq_ready),
    .io_deq_valid(q_631_io_deq_valid),
    .io_deq_bits(q_631_io_deq_bits)
  );
  Queue q_632 ( // @[Decoupled.scala 361:21]
    .clock(q_632_clock),
    .reset(q_632_reset),
    .io_enq_ready(q_632_io_enq_ready),
    .io_enq_valid(q_632_io_enq_valid),
    .io_enq_bits(q_632_io_enq_bits),
    .io_deq_ready(q_632_io_deq_ready),
    .io_deq_valid(q_632_io_deq_valid),
    .io_deq_bits(q_632_io_deq_bits)
  );
  Queue q_633 ( // @[Decoupled.scala 361:21]
    .clock(q_633_clock),
    .reset(q_633_reset),
    .io_enq_ready(q_633_io_enq_ready),
    .io_enq_valid(q_633_io_enq_valid),
    .io_enq_bits(q_633_io_enq_bits),
    .io_deq_ready(q_633_io_deq_ready),
    .io_deq_valid(q_633_io_deq_valid),
    .io_deq_bits(q_633_io_deq_bits)
  );
  Queue q_634 ( // @[Decoupled.scala 361:21]
    .clock(q_634_clock),
    .reset(q_634_reset),
    .io_enq_ready(q_634_io_enq_ready),
    .io_enq_valid(q_634_io_enq_valid),
    .io_enq_bits(q_634_io_enq_bits),
    .io_deq_ready(q_634_io_deq_ready),
    .io_deq_valid(q_634_io_deq_valid),
    .io_deq_bits(q_634_io_deq_bits)
  );
  Queue q_635 ( // @[Decoupled.scala 361:21]
    .clock(q_635_clock),
    .reset(q_635_reset),
    .io_enq_ready(q_635_io_enq_ready),
    .io_enq_valid(q_635_io_enq_valid),
    .io_enq_bits(q_635_io_enq_bits),
    .io_deq_ready(q_635_io_deq_ready),
    .io_deq_valid(q_635_io_deq_valid),
    .io_deq_bits(q_635_io_deq_bits)
  );
  Queue q_636 ( // @[Decoupled.scala 361:21]
    .clock(q_636_clock),
    .reset(q_636_reset),
    .io_enq_ready(q_636_io_enq_ready),
    .io_enq_valid(q_636_io_enq_valid),
    .io_enq_bits(q_636_io_enq_bits),
    .io_deq_ready(q_636_io_deq_ready),
    .io_deq_valid(q_636_io_deq_valid),
    .io_deq_bits(q_636_io_deq_bits)
  );
  Queue q_637 ( // @[Decoupled.scala 361:21]
    .clock(q_637_clock),
    .reset(q_637_reset),
    .io_enq_ready(q_637_io_enq_ready),
    .io_enq_valid(q_637_io_enq_valid),
    .io_enq_bits(q_637_io_enq_bits),
    .io_deq_ready(q_637_io_deq_ready),
    .io_deq_valid(q_637_io_deq_valid),
    .io_deq_bits(q_637_io_deq_bits)
  );
  Queue q_638 ( // @[Decoupled.scala 361:21]
    .clock(q_638_clock),
    .reset(q_638_reset),
    .io_enq_ready(q_638_io_enq_ready),
    .io_enq_valid(q_638_io_enq_valid),
    .io_enq_bits(q_638_io_enq_bits),
    .io_deq_ready(q_638_io_deq_ready),
    .io_deq_valid(q_638_io_deq_valid),
    .io_deq_bits(q_638_io_deq_bits)
  );
  Queue q_639 ( // @[Decoupled.scala 361:21]
    .clock(q_639_clock),
    .reset(q_639_reset),
    .io_enq_ready(q_639_io_enq_ready),
    .io_enq_valid(q_639_io_enq_valid),
    .io_enq_bits(q_639_io_enq_bits),
    .io_deq_ready(q_639_io_deq_ready),
    .io_deq_valid(q_639_io_deq_valid),
    .io_deq_bits(q_639_io_deq_bits)
  );
  Queue q_640 ( // @[Decoupled.scala 361:21]
    .clock(q_640_clock),
    .reset(q_640_reset),
    .io_enq_ready(q_640_io_enq_ready),
    .io_enq_valid(q_640_io_enq_valid),
    .io_enq_bits(q_640_io_enq_bits),
    .io_deq_ready(q_640_io_deq_ready),
    .io_deq_valid(q_640_io_deq_valid),
    .io_deq_bits(q_640_io_deq_bits)
  );
  Queue q_641 ( // @[Decoupled.scala 361:21]
    .clock(q_641_clock),
    .reset(q_641_reset),
    .io_enq_ready(q_641_io_enq_ready),
    .io_enq_valid(q_641_io_enq_valid),
    .io_enq_bits(q_641_io_enq_bits),
    .io_deq_ready(q_641_io_deq_ready),
    .io_deq_valid(q_641_io_deq_valid),
    .io_deq_bits(q_641_io_deq_bits)
  );
  Queue q_642 ( // @[Decoupled.scala 361:21]
    .clock(q_642_clock),
    .reset(q_642_reset),
    .io_enq_ready(q_642_io_enq_ready),
    .io_enq_valid(q_642_io_enq_valid),
    .io_enq_bits(q_642_io_enq_bits),
    .io_deq_ready(q_642_io_deq_ready),
    .io_deq_valid(q_642_io_deq_valid),
    .io_deq_bits(q_642_io_deq_bits)
  );
  Queue q_643 ( // @[Decoupled.scala 361:21]
    .clock(q_643_clock),
    .reset(q_643_reset),
    .io_enq_ready(q_643_io_enq_ready),
    .io_enq_valid(q_643_io_enq_valid),
    .io_enq_bits(q_643_io_enq_bits),
    .io_deq_ready(q_643_io_deq_ready),
    .io_deq_valid(q_643_io_deq_valid),
    .io_deq_bits(q_643_io_deq_bits)
  );
  Queue q_644 ( // @[Decoupled.scala 361:21]
    .clock(q_644_clock),
    .reset(q_644_reset),
    .io_enq_ready(q_644_io_enq_ready),
    .io_enq_valid(q_644_io_enq_valid),
    .io_enq_bits(q_644_io_enq_bits),
    .io_deq_ready(q_644_io_deq_ready),
    .io_deq_valid(q_644_io_deq_valid),
    .io_deq_bits(q_644_io_deq_bits)
  );
  Queue q_645 ( // @[Decoupled.scala 361:21]
    .clock(q_645_clock),
    .reset(q_645_reset),
    .io_enq_ready(q_645_io_enq_ready),
    .io_enq_valid(q_645_io_enq_valid),
    .io_enq_bits(q_645_io_enq_bits),
    .io_deq_ready(q_645_io_deq_ready),
    .io_deq_valid(q_645_io_deq_valid),
    .io_deq_bits(q_645_io_deq_bits)
  );
  Queue q_646 ( // @[Decoupled.scala 361:21]
    .clock(q_646_clock),
    .reset(q_646_reset),
    .io_enq_ready(q_646_io_enq_ready),
    .io_enq_valid(q_646_io_enq_valid),
    .io_enq_bits(q_646_io_enq_bits),
    .io_deq_ready(q_646_io_deq_ready),
    .io_deq_valid(q_646_io_deq_valid),
    .io_deq_bits(q_646_io_deq_bits)
  );
  Queue q_647 ( // @[Decoupled.scala 361:21]
    .clock(q_647_clock),
    .reset(q_647_reset),
    .io_enq_ready(q_647_io_enq_ready),
    .io_enq_valid(q_647_io_enq_valid),
    .io_enq_bits(q_647_io_enq_bits),
    .io_deq_ready(q_647_io_deq_ready),
    .io_deq_valid(q_647_io_deq_valid),
    .io_deq_bits(q_647_io_deq_bits)
  );
  Queue q_648 ( // @[Decoupled.scala 361:21]
    .clock(q_648_clock),
    .reset(q_648_reset),
    .io_enq_ready(q_648_io_enq_ready),
    .io_enq_valid(q_648_io_enq_valid),
    .io_enq_bits(q_648_io_enq_bits),
    .io_deq_ready(q_648_io_deq_ready),
    .io_deq_valid(q_648_io_deq_valid),
    .io_deq_bits(q_648_io_deq_bits)
  );
  Queue q_649 ( // @[Decoupled.scala 361:21]
    .clock(q_649_clock),
    .reset(q_649_reset),
    .io_enq_ready(q_649_io_enq_ready),
    .io_enq_valid(q_649_io_enq_valid),
    .io_enq_bits(q_649_io_enq_bits),
    .io_deq_ready(q_649_io_deq_ready),
    .io_deq_valid(q_649_io_deq_valid),
    .io_deq_bits(q_649_io_deq_bits)
  );
  Queue q_650 ( // @[Decoupled.scala 361:21]
    .clock(q_650_clock),
    .reset(q_650_reset),
    .io_enq_ready(q_650_io_enq_ready),
    .io_enq_valid(q_650_io_enq_valid),
    .io_enq_bits(q_650_io_enq_bits),
    .io_deq_ready(q_650_io_deq_ready),
    .io_deq_valid(q_650_io_deq_valid),
    .io_deq_bits(q_650_io_deq_bits)
  );
  Queue q_651 ( // @[Decoupled.scala 361:21]
    .clock(q_651_clock),
    .reset(q_651_reset),
    .io_enq_ready(q_651_io_enq_ready),
    .io_enq_valid(q_651_io_enq_valid),
    .io_enq_bits(q_651_io_enq_bits),
    .io_deq_ready(q_651_io_deq_ready),
    .io_deq_valid(q_651_io_deq_valid),
    .io_deq_bits(q_651_io_deq_bits)
  );
  Queue q_652 ( // @[Decoupled.scala 361:21]
    .clock(q_652_clock),
    .reset(q_652_reset),
    .io_enq_ready(q_652_io_enq_ready),
    .io_enq_valid(q_652_io_enq_valid),
    .io_enq_bits(q_652_io_enq_bits),
    .io_deq_ready(q_652_io_deq_ready),
    .io_deq_valid(q_652_io_deq_valid),
    .io_deq_bits(q_652_io_deq_bits)
  );
  Queue q_653 ( // @[Decoupled.scala 361:21]
    .clock(q_653_clock),
    .reset(q_653_reset),
    .io_enq_ready(q_653_io_enq_ready),
    .io_enq_valid(q_653_io_enq_valid),
    .io_enq_bits(q_653_io_enq_bits),
    .io_deq_ready(q_653_io_deq_ready),
    .io_deq_valid(q_653_io_deq_valid),
    .io_deq_bits(q_653_io_deq_bits)
  );
  Queue q_654 ( // @[Decoupled.scala 361:21]
    .clock(q_654_clock),
    .reset(q_654_reset),
    .io_enq_ready(q_654_io_enq_ready),
    .io_enq_valid(q_654_io_enq_valid),
    .io_enq_bits(q_654_io_enq_bits),
    .io_deq_ready(q_654_io_deq_ready),
    .io_deq_valid(q_654_io_deq_valid),
    .io_deq_bits(q_654_io_deq_bits)
  );
  Queue q_655 ( // @[Decoupled.scala 361:21]
    .clock(q_655_clock),
    .reset(q_655_reset),
    .io_enq_ready(q_655_io_enq_ready),
    .io_enq_valid(q_655_io_enq_valid),
    .io_enq_bits(q_655_io_enq_bits),
    .io_deq_ready(q_655_io_deq_ready),
    .io_deq_valid(q_655_io_deq_valid),
    .io_deq_bits(q_655_io_deq_bits)
  );
  Queue q_656 ( // @[Decoupled.scala 361:21]
    .clock(q_656_clock),
    .reset(q_656_reset),
    .io_enq_ready(q_656_io_enq_ready),
    .io_enq_valid(q_656_io_enq_valid),
    .io_enq_bits(q_656_io_enq_bits),
    .io_deq_ready(q_656_io_deq_ready),
    .io_deq_valid(q_656_io_deq_valid),
    .io_deq_bits(q_656_io_deq_bits)
  );
  Queue q_657 ( // @[Decoupled.scala 361:21]
    .clock(q_657_clock),
    .reset(q_657_reset),
    .io_enq_ready(q_657_io_enq_ready),
    .io_enq_valid(q_657_io_enq_valid),
    .io_enq_bits(q_657_io_enq_bits),
    .io_deq_ready(q_657_io_deq_ready),
    .io_deq_valid(q_657_io_deq_valid),
    .io_deq_bits(q_657_io_deq_bits)
  );
  Queue q_658 ( // @[Decoupled.scala 361:21]
    .clock(q_658_clock),
    .reset(q_658_reset),
    .io_enq_ready(q_658_io_enq_ready),
    .io_enq_valid(q_658_io_enq_valid),
    .io_enq_bits(q_658_io_enq_bits),
    .io_deq_ready(q_658_io_deq_ready),
    .io_deq_valid(q_658_io_deq_valid),
    .io_deq_bits(q_658_io_deq_bits)
  );
  Queue q_659 ( // @[Decoupled.scala 361:21]
    .clock(q_659_clock),
    .reset(q_659_reset),
    .io_enq_ready(q_659_io_enq_ready),
    .io_enq_valid(q_659_io_enq_valid),
    .io_enq_bits(q_659_io_enq_bits),
    .io_deq_ready(q_659_io_deq_ready),
    .io_deq_valid(q_659_io_deq_valid),
    .io_deq_bits(q_659_io_deq_bits)
  );
  Queue q_660 ( // @[Decoupled.scala 361:21]
    .clock(q_660_clock),
    .reset(q_660_reset),
    .io_enq_ready(q_660_io_enq_ready),
    .io_enq_valid(q_660_io_enq_valid),
    .io_enq_bits(q_660_io_enq_bits),
    .io_deq_ready(q_660_io_deq_ready),
    .io_deq_valid(q_660_io_deq_valid),
    .io_deq_bits(q_660_io_deq_bits)
  );
  Queue q_661 ( // @[Decoupled.scala 361:21]
    .clock(q_661_clock),
    .reset(q_661_reset),
    .io_enq_ready(q_661_io_enq_ready),
    .io_enq_valid(q_661_io_enq_valid),
    .io_enq_bits(q_661_io_enq_bits),
    .io_deq_ready(q_661_io_deq_ready),
    .io_deq_valid(q_661_io_deq_valid),
    .io_deq_bits(q_661_io_deq_bits)
  );
  Queue q_662 ( // @[Decoupled.scala 361:21]
    .clock(q_662_clock),
    .reset(q_662_reset),
    .io_enq_ready(q_662_io_enq_ready),
    .io_enq_valid(q_662_io_enq_valid),
    .io_enq_bits(q_662_io_enq_bits),
    .io_deq_ready(q_662_io_deq_ready),
    .io_deq_valid(q_662_io_deq_valid),
    .io_deq_bits(q_662_io_deq_bits)
  );
  Queue q_663 ( // @[Decoupled.scala 361:21]
    .clock(q_663_clock),
    .reset(q_663_reset),
    .io_enq_ready(q_663_io_enq_ready),
    .io_enq_valid(q_663_io_enq_valid),
    .io_enq_bits(q_663_io_enq_bits),
    .io_deq_ready(q_663_io_deq_ready),
    .io_deq_valid(q_663_io_deq_valid),
    .io_deq_bits(q_663_io_deq_bits)
  );
  Queue q_664 ( // @[Decoupled.scala 361:21]
    .clock(q_664_clock),
    .reset(q_664_reset),
    .io_enq_ready(q_664_io_enq_ready),
    .io_enq_valid(q_664_io_enq_valid),
    .io_enq_bits(q_664_io_enq_bits),
    .io_deq_ready(q_664_io_deq_ready),
    .io_deq_valid(q_664_io_deq_valid),
    .io_deq_bits(q_664_io_deq_bits)
  );
  Queue q_665 ( // @[Decoupled.scala 361:21]
    .clock(q_665_clock),
    .reset(q_665_reset),
    .io_enq_ready(q_665_io_enq_ready),
    .io_enq_valid(q_665_io_enq_valid),
    .io_enq_bits(q_665_io_enq_bits),
    .io_deq_ready(q_665_io_deq_ready),
    .io_deq_valid(q_665_io_deq_valid),
    .io_deq_bits(q_665_io_deq_bits)
  );
  Queue q_666 ( // @[Decoupled.scala 361:21]
    .clock(q_666_clock),
    .reset(q_666_reset),
    .io_enq_ready(q_666_io_enq_ready),
    .io_enq_valid(q_666_io_enq_valid),
    .io_enq_bits(q_666_io_enq_bits),
    .io_deq_ready(q_666_io_deq_ready),
    .io_deq_valid(q_666_io_deq_valid),
    .io_deq_bits(q_666_io_deq_bits)
  );
  Queue q_667 ( // @[Decoupled.scala 361:21]
    .clock(q_667_clock),
    .reset(q_667_reset),
    .io_enq_ready(q_667_io_enq_ready),
    .io_enq_valid(q_667_io_enq_valid),
    .io_enq_bits(q_667_io_enq_bits),
    .io_deq_ready(q_667_io_deq_ready),
    .io_deq_valid(q_667_io_deq_valid),
    .io_deq_bits(q_667_io_deq_bits)
  );
  Queue q_668 ( // @[Decoupled.scala 361:21]
    .clock(q_668_clock),
    .reset(q_668_reset),
    .io_enq_ready(q_668_io_enq_ready),
    .io_enq_valid(q_668_io_enq_valid),
    .io_enq_bits(q_668_io_enq_bits),
    .io_deq_ready(q_668_io_deq_ready),
    .io_deq_valid(q_668_io_deq_valid),
    .io_deq_bits(q_668_io_deq_bits)
  );
  Queue q_669 ( // @[Decoupled.scala 361:21]
    .clock(q_669_clock),
    .reset(q_669_reset),
    .io_enq_ready(q_669_io_enq_ready),
    .io_enq_valid(q_669_io_enq_valid),
    .io_enq_bits(q_669_io_enq_bits),
    .io_deq_ready(q_669_io_deq_ready),
    .io_deq_valid(q_669_io_deq_valid),
    .io_deq_bits(q_669_io_deq_bits)
  );
  Queue q_670 ( // @[Decoupled.scala 361:21]
    .clock(q_670_clock),
    .reset(q_670_reset),
    .io_enq_ready(q_670_io_enq_ready),
    .io_enq_valid(q_670_io_enq_valid),
    .io_enq_bits(q_670_io_enq_bits),
    .io_deq_ready(q_670_io_deq_ready),
    .io_deq_valid(q_670_io_deq_valid),
    .io_deq_bits(q_670_io_deq_bits)
  );
  Queue q_671 ( // @[Decoupled.scala 361:21]
    .clock(q_671_clock),
    .reset(q_671_reset),
    .io_enq_ready(q_671_io_enq_ready),
    .io_enq_valid(q_671_io_enq_valid),
    .io_enq_bits(q_671_io_enq_bits),
    .io_deq_ready(q_671_io_deq_ready),
    .io_deq_valid(q_671_io_deq_valid),
    .io_deq_bits(q_671_io_deq_bits)
  );
  Queue q_672 ( // @[Decoupled.scala 361:21]
    .clock(q_672_clock),
    .reset(q_672_reset),
    .io_enq_ready(q_672_io_enq_ready),
    .io_enq_valid(q_672_io_enq_valid),
    .io_enq_bits(q_672_io_enq_bits),
    .io_deq_ready(q_672_io_deq_ready),
    .io_deq_valid(q_672_io_deq_valid),
    .io_deq_bits(q_672_io_deq_bits)
  );
  Queue q_673 ( // @[Decoupled.scala 361:21]
    .clock(q_673_clock),
    .reset(q_673_reset),
    .io_enq_ready(q_673_io_enq_ready),
    .io_enq_valid(q_673_io_enq_valid),
    .io_enq_bits(q_673_io_enq_bits),
    .io_deq_ready(q_673_io_deq_ready),
    .io_deq_valid(q_673_io_deq_valid),
    .io_deq_bits(q_673_io_deq_bits)
  );
  Queue q_674 ( // @[Decoupled.scala 361:21]
    .clock(q_674_clock),
    .reset(q_674_reset),
    .io_enq_ready(q_674_io_enq_ready),
    .io_enq_valid(q_674_io_enq_valid),
    .io_enq_bits(q_674_io_enq_bits),
    .io_deq_ready(q_674_io_deq_ready),
    .io_deq_valid(q_674_io_deq_valid),
    .io_deq_bits(q_674_io_deq_bits)
  );
  Queue q_675 ( // @[Decoupled.scala 361:21]
    .clock(q_675_clock),
    .reset(q_675_reset),
    .io_enq_ready(q_675_io_enq_ready),
    .io_enq_valid(q_675_io_enq_valid),
    .io_enq_bits(q_675_io_enq_bits),
    .io_deq_ready(q_675_io_deq_ready),
    .io_deq_valid(q_675_io_deq_valid),
    .io_deq_bits(q_675_io_deq_bits)
  );
  Queue q_676 ( // @[Decoupled.scala 361:21]
    .clock(q_676_clock),
    .reset(q_676_reset),
    .io_enq_ready(q_676_io_enq_ready),
    .io_enq_valid(q_676_io_enq_valid),
    .io_enq_bits(q_676_io_enq_bits),
    .io_deq_ready(q_676_io_deq_ready),
    .io_deq_valid(q_676_io_deq_valid),
    .io_deq_bits(q_676_io_deq_bits)
  );
  Queue q_677 ( // @[Decoupled.scala 361:21]
    .clock(q_677_clock),
    .reset(q_677_reset),
    .io_enq_ready(q_677_io_enq_ready),
    .io_enq_valid(q_677_io_enq_valid),
    .io_enq_bits(q_677_io_enq_bits),
    .io_deq_ready(q_677_io_deq_ready),
    .io_deq_valid(q_677_io_deq_valid),
    .io_deq_bits(q_677_io_deq_bits)
  );
  Queue q_678 ( // @[Decoupled.scala 361:21]
    .clock(q_678_clock),
    .reset(q_678_reset),
    .io_enq_ready(q_678_io_enq_ready),
    .io_enq_valid(q_678_io_enq_valid),
    .io_enq_bits(q_678_io_enq_bits),
    .io_deq_ready(q_678_io_deq_ready),
    .io_deq_valid(q_678_io_deq_valid),
    .io_deq_bits(q_678_io_deq_bits)
  );
  Queue q_679 ( // @[Decoupled.scala 361:21]
    .clock(q_679_clock),
    .reset(q_679_reset),
    .io_enq_ready(q_679_io_enq_ready),
    .io_enq_valid(q_679_io_enq_valid),
    .io_enq_bits(q_679_io_enq_bits),
    .io_deq_ready(q_679_io_deq_ready),
    .io_deq_valid(q_679_io_deq_valid),
    .io_deq_bits(q_679_io_deq_bits)
  );
  Queue q_680 ( // @[Decoupled.scala 361:21]
    .clock(q_680_clock),
    .reset(q_680_reset),
    .io_enq_ready(q_680_io_enq_ready),
    .io_enq_valid(q_680_io_enq_valid),
    .io_enq_bits(q_680_io_enq_bits),
    .io_deq_ready(q_680_io_deq_ready),
    .io_deq_valid(q_680_io_deq_valid),
    .io_deq_bits(q_680_io_deq_bits)
  );
  Queue q_681 ( // @[Decoupled.scala 361:21]
    .clock(q_681_clock),
    .reset(q_681_reset),
    .io_enq_ready(q_681_io_enq_ready),
    .io_enq_valid(q_681_io_enq_valid),
    .io_enq_bits(q_681_io_enq_bits),
    .io_deq_ready(q_681_io_deq_ready),
    .io_deq_valid(q_681_io_deq_valid),
    .io_deq_bits(q_681_io_deq_bits)
  );
  Queue q_682 ( // @[Decoupled.scala 361:21]
    .clock(q_682_clock),
    .reset(q_682_reset),
    .io_enq_ready(q_682_io_enq_ready),
    .io_enq_valid(q_682_io_enq_valid),
    .io_enq_bits(q_682_io_enq_bits),
    .io_deq_ready(q_682_io_deq_ready),
    .io_deq_valid(q_682_io_deq_valid),
    .io_deq_bits(q_682_io_deq_bits)
  );
  Queue q_683 ( // @[Decoupled.scala 361:21]
    .clock(q_683_clock),
    .reset(q_683_reset),
    .io_enq_ready(q_683_io_enq_ready),
    .io_enq_valid(q_683_io_enq_valid),
    .io_enq_bits(q_683_io_enq_bits),
    .io_deq_ready(q_683_io_deq_ready),
    .io_deq_valid(q_683_io_deq_valid),
    .io_deq_bits(q_683_io_deq_bits)
  );
  Queue q_684 ( // @[Decoupled.scala 361:21]
    .clock(q_684_clock),
    .reset(q_684_reset),
    .io_enq_ready(q_684_io_enq_ready),
    .io_enq_valid(q_684_io_enq_valid),
    .io_enq_bits(q_684_io_enq_bits),
    .io_deq_ready(q_684_io_deq_ready),
    .io_deq_valid(q_684_io_deq_valid),
    .io_deq_bits(q_684_io_deq_bits)
  );
  Queue q_685 ( // @[Decoupled.scala 361:21]
    .clock(q_685_clock),
    .reset(q_685_reset),
    .io_enq_ready(q_685_io_enq_ready),
    .io_enq_valid(q_685_io_enq_valid),
    .io_enq_bits(q_685_io_enq_bits),
    .io_deq_ready(q_685_io_deq_ready),
    .io_deq_valid(q_685_io_deq_valid),
    .io_deq_bits(q_685_io_deq_bits)
  );
  Queue q_686 ( // @[Decoupled.scala 361:21]
    .clock(q_686_clock),
    .reset(q_686_reset),
    .io_enq_ready(q_686_io_enq_ready),
    .io_enq_valid(q_686_io_enq_valid),
    .io_enq_bits(q_686_io_enq_bits),
    .io_deq_ready(q_686_io_deq_ready),
    .io_deq_valid(q_686_io_deq_valid),
    .io_deq_bits(q_686_io_deq_bits)
  );
  Queue q_687 ( // @[Decoupled.scala 361:21]
    .clock(q_687_clock),
    .reset(q_687_reset),
    .io_enq_ready(q_687_io_enq_ready),
    .io_enq_valid(q_687_io_enq_valid),
    .io_enq_bits(q_687_io_enq_bits),
    .io_deq_ready(q_687_io_deq_ready),
    .io_deq_valid(q_687_io_deq_valid),
    .io_deq_bits(q_687_io_deq_bits)
  );
  Queue q_688 ( // @[Decoupled.scala 361:21]
    .clock(q_688_clock),
    .reset(q_688_reset),
    .io_enq_ready(q_688_io_enq_ready),
    .io_enq_valid(q_688_io_enq_valid),
    .io_enq_bits(q_688_io_enq_bits),
    .io_deq_ready(q_688_io_deq_ready),
    .io_deq_valid(q_688_io_deq_valid),
    .io_deq_bits(q_688_io_deq_bits)
  );
  Queue q_689 ( // @[Decoupled.scala 361:21]
    .clock(q_689_clock),
    .reset(q_689_reset),
    .io_enq_ready(q_689_io_enq_ready),
    .io_enq_valid(q_689_io_enq_valid),
    .io_enq_bits(q_689_io_enq_bits),
    .io_deq_ready(q_689_io_deq_ready),
    .io_deq_valid(q_689_io_deq_valid),
    .io_deq_bits(q_689_io_deq_bits)
  );
  Queue q_690 ( // @[Decoupled.scala 361:21]
    .clock(q_690_clock),
    .reset(q_690_reset),
    .io_enq_ready(q_690_io_enq_ready),
    .io_enq_valid(q_690_io_enq_valid),
    .io_enq_bits(q_690_io_enq_bits),
    .io_deq_ready(q_690_io_deq_ready),
    .io_deq_valid(q_690_io_deq_valid),
    .io_deq_bits(q_690_io_deq_bits)
  );
  Queue q_691 ( // @[Decoupled.scala 361:21]
    .clock(q_691_clock),
    .reset(q_691_reset),
    .io_enq_ready(q_691_io_enq_ready),
    .io_enq_valid(q_691_io_enq_valid),
    .io_enq_bits(q_691_io_enq_bits),
    .io_deq_ready(q_691_io_deq_ready),
    .io_deq_valid(q_691_io_deq_valid),
    .io_deq_bits(q_691_io_deq_bits)
  );
  Queue q_692 ( // @[Decoupled.scala 361:21]
    .clock(q_692_clock),
    .reset(q_692_reset),
    .io_enq_ready(q_692_io_enq_ready),
    .io_enq_valid(q_692_io_enq_valid),
    .io_enq_bits(q_692_io_enq_bits),
    .io_deq_ready(q_692_io_deq_ready),
    .io_deq_valid(q_692_io_deq_valid),
    .io_deq_bits(q_692_io_deq_bits)
  );
  Queue q_693 ( // @[Decoupled.scala 361:21]
    .clock(q_693_clock),
    .reset(q_693_reset),
    .io_enq_ready(q_693_io_enq_ready),
    .io_enq_valid(q_693_io_enq_valid),
    .io_enq_bits(q_693_io_enq_bits),
    .io_deq_ready(q_693_io_deq_ready),
    .io_deq_valid(q_693_io_deq_valid),
    .io_deq_bits(q_693_io_deq_bits)
  );
  Queue q_694 ( // @[Decoupled.scala 361:21]
    .clock(q_694_clock),
    .reset(q_694_reset),
    .io_enq_ready(q_694_io_enq_ready),
    .io_enq_valid(q_694_io_enq_valid),
    .io_enq_bits(q_694_io_enq_bits),
    .io_deq_ready(q_694_io_deq_ready),
    .io_deq_valid(q_694_io_deq_valid),
    .io_deq_bits(q_694_io_deq_bits)
  );
  Queue q_695 ( // @[Decoupled.scala 361:21]
    .clock(q_695_clock),
    .reset(q_695_reset),
    .io_enq_ready(q_695_io_enq_ready),
    .io_enq_valid(q_695_io_enq_valid),
    .io_enq_bits(q_695_io_enq_bits),
    .io_deq_ready(q_695_io_deq_ready),
    .io_deq_valid(q_695_io_deq_valid),
    .io_deq_bits(q_695_io_deq_bits)
  );
  Queue q_696 ( // @[Decoupled.scala 361:21]
    .clock(q_696_clock),
    .reset(q_696_reset),
    .io_enq_ready(q_696_io_enq_ready),
    .io_enq_valid(q_696_io_enq_valid),
    .io_enq_bits(q_696_io_enq_bits),
    .io_deq_ready(q_696_io_deq_ready),
    .io_deq_valid(q_696_io_deq_valid),
    .io_deq_bits(q_696_io_deq_bits)
  );
  Queue q_697 ( // @[Decoupled.scala 361:21]
    .clock(q_697_clock),
    .reset(q_697_reset),
    .io_enq_ready(q_697_io_enq_ready),
    .io_enq_valid(q_697_io_enq_valid),
    .io_enq_bits(q_697_io_enq_bits),
    .io_deq_ready(q_697_io_deq_ready),
    .io_deq_valid(q_697_io_deq_valid),
    .io_deq_bits(q_697_io_deq_bits)
  );
  Queue q_698 ( // @[Decoupled.scala 361:21]
    .clock(q_698_clock),
    .reset(q_698_reset),
    .io_enq_ready(q_698_io_enq_ready),
    .io_enq_valid(q_698_io_enq_valid),
    .io_enq_bits(q_698_io_enq_bits),
    .io_deq_ready(q_698_io_deq_ready),
    .io_deq_valid(q_698_io_deq_valid),
    .io_deq_bits(q_698_io_deq_bits)
  );
  Queue q_699 ( // @[Decoupled.scala 361:21]
    .clock(q_699_clock),
    .reset(q_699_reset),
    .io_enq_ready(q_699_io_enq_ready),
    .io_enq_valid(q_699_io_enq_valid),
    .io_enq_bits(q_699_io_enq_bits),
    .io_deq_ready(q_699_io_deq_ready),
    .io_deq_valid(q_699_io_deq_valid),
    .io_deq_bits(q_699_io_deq_bits)
  );
  Queue q_700 ( // @[Decoupled.scala 361:21]
    .clock(q_700_clock),
    .reset(q_700_reset),
    .io_enq_ready(q_700_io_enq_ready),
    .io_enq_valid(q_700_io_enq_valid),
    .io_enq_bits(q_700_io_enq_bits),
    .io_deq_ready(q_700_io_deq_ready),
    .io_deq_valid(q_700_io_deq_valid),
    .io_deq_bits(q_700_io_deq_bits)
  );
  Queue q_701 ( // @[Decoupled.scala 361:21]
    .clock(q_701_clock),
    .reset(q_701_reset),
    .io_enq_ready(q_701_io_enq_ready),
    .io_enq_valid(q_701_io_enq_valid),
    .io_enq_bits(q_701_io_enq_bits),
    .io_deq_ready(q_701_io_deq_ready),
    .io_deq_valid(q_701_io_deq_valid),
    .io_deq_bits(q_701_io_deq_bits)
  );
  Queue q_702 ( // @[Decoupled.scala 361:21]
    .clock(q_702_clock),
    .reset(q_702_reset),
    .io_enq_ready(q_702_io_enq_ready),
    .io_enq_valid(q_702_io_enq_valid),
    .io_enq_bits(q_702_io_enq_bits),
    .io_deq_ready(q_702_io_deq_ready),
    .io_deq_valid(q_702_io_deq_valid),
    .io_deq_bits(q_702_io_deq_bits)
  );
  Queue q_703 ( // @[Decoupled.scala 361:21]
    .clock(q_703_clock),
    .reset(q_703_reset),
    .io_enq_ready(q_703_io_enq_ready),
    .io_enq_valid(q_703_io_enq_valid),
    .io_enq_bits(q_703_io_enq_bits),
    .io_deq_ready(q_703_io_deq_ready),
    .io_deq_valid(q_703_io_deq_valid),
    .io_deq_bits(q_703_io_deq_bits)
  );
  Queue q_704 ( // @[Decoupled.scala 361:21]
    .clock(q_704_clock),
    .reset(q_704_reset),
    .io_enq_ready(q_704_io_enq_ready),
    .io_enq_valid(q_704_io_enq_valid),
    .io_enq_bits(q_704_io_enq_bits),
    .io_deq_ready(q_704_io_deq_ready),
    .io_deq_valid(q_704_io_deq_valid),
    .io_deq_bits(q_704_io_deq_bits)
  );
  Queue q_705 ( // @[Decoupled.scala 361:21]
    .clock(q_705_clock),
    .reset(q_705_reset),
    .io_enq_ready(q_705_io_enq_ready),
    .io_enq_valid(q_705_io_enq_valid),
    .io_enq_bits(q_705_io_enq_bits),
    .io_deq_ready(q_705_io_deq_ready),
    .io_deq_valid(q_705_io_deq_valid),
    .io_deq_bits(q_705_io_deq_bits)
  );
  Queue q_706 ( // @[Decoupled.scala 361:21]
    .clock(q_706_clock),
    .reset(q_706_reset),
    .io_enq_ready(q_706_io_enq_ready),
    .io_enq_valid(q_706_io_enq_valid),
    .io_enq_bits(q_706_io_enq_bits),
    .io_deq_ready(q_706_io_deq_ready),
    .io_deq_valid(q_706_io_deq_valid),
    .io_deq_bits(q_706_io_deq_bits)
  );
  Queue q_707 ( // @[Decoupled.scala 361:21]
    .clock(q_707_clock),
    .reset(q_707_reset),
    .io_enq_ready(q_707_io_enq_ready),
    .io_enq_valid(q_707_io_enq_valid),
    .io_enq_bits(q_707_io_enq_bits),
    .io_deq_ready(q_707_io_deq_ready),
    .io_deq_valid(q_707_io_deq_valid),
    .io_deq_bits(q_707_io_deq_bits)
  );
  Queue q_708 ( // @[Decoupled.scala 361:21]
    .clock(q_708_clock),
    .reset(q_708_reset),
    .io_enq_ready(q_708_io_enq_ready),
    .io_enq_valid(q_708_io_enq_valid),
    .io_enq_bits(q_708_io_enq_bits),
    .io_deq_ready(q_708_io_deq_ready),
    .io_deq_valid(q_708_io_deq_valid),
    .io_deq_bits(q_708_io_deq_bits)
  );
  Queue q_709 ( // @[Decoupled.scala 361:21]
    .clock(q_709_clock),
    .reset(q_709_reset),
    .io_enq_ready(q_709_io_enq_ready),
    .io_enq_valid(q_709_io_enq_valid),
    .io_enq_bits(q_709_io_enq_bits),
    .io_deq_ready(q_709_io_deq_ready),
    .io_deq_valid(q_709_io_deq_valid),
    .io_deq_bits(q_709_io_deq_bits)
  );
  Queue q_710 ( // @[Decoupled.scala 361:21]
    .clock(q_710_clock),
    .reset(q_710_reset),
    .io_enq_ready(q_710_io_enq_ready),
    .io_enq_valid(q_710_io_enq_valid),
    .io_enq_bits(q_710_io_enq_bits),
    .io_deq_ready(q_710_io_deq_ready),
    .io_deq_valid(q_710_io_deq_valid),
    .io_deq_bits(q_710_io_deq_bits)
  );
  Queue q_711 ( // @[Decoupled.scala 361:21]
    .clock(q_711_clock),
    .reset(q_711_reset),
    .io_enq_ready(q_711_io_enq_ready),
    .io_enq_valid(q_711_io_enq_valid),
    .io_enq_bits(q_711_io_enq_bits),
    .io_deq_ready(q_711_io_deq_ready),
    .io_deq_valid(q_711_io_deq_valid),
    .io_deq_bits(q_711_io_deq_bits)
  );
  Queue q_712 ( // @[Decoupled.scala 361:21]
    .clock(q_712_clock),
    .reset(q_712_reset),
    .io_enq_ready(q_712_io_enq_ready),
    .io_enq_valid(q_712_io_enq_valid),
    .io_enq_bits(q_712_io_enq_bits),
    .io_deq_ready(q_712_io_deq_ready),
    .io_deq_valid(q_712_io_deq_valid),
    .io_deq_bits(q_712_io_deq_bits)
  );
  Queue q_713 ( // @[Decoupled.scala 361:21]
    .clock(q_713_clock),
    .reset(q_713_reset),
    .io_enq_ready(q_713_io_enq_ready),
    .io_enq_valid(q_713_io_enq_valid),
    .io_enq_bits(q_713_io_enq_bits),
    .io_deq_ready(q_713_io_deq_ready),
    .io_deq_valid(q_713_io_deq_valid),
    .io_deq_bits(q_713_io_deq_bits)
  );
  Queue q_714 ( // @[Decoupled.scala 361:21]
    .clock(q_714_clock),
    .reset(q_714_reset),
    .io_enq_ready(q_714_io_enq_ready),
    .io_enq_valid(q_714_io_enq_valid),
    .io_enq_bits(q_714_io_enq_bits),
    .io_deq_ready(q_714_io_deq_ready),
    .io_deq_valid(q_714_io_deq_valid),
    .io_deq_bits(q_714_io_deq_bits)
  );
  Queue q_715 ( // @[Decoupled.scala 361:21]
    .clock(q_715_clock),
    .reset(q_715_reset),
    .io_enq_ready(q_715_io_enq_ready),
    .io_enq_valid(q_715_io_enq_valid),
    .io_enq_bits(q_715_io_enq_bits),
    .io_deq_ready(q_715_io_deq_ready),
    .io_deq_valid(q_715_io_deq_valid),
    .io_deq_bits(q_715_io_deq_bits)
  );
  Queue q_716 ( // @[Decoupled.scala 361:21]
    .clock(q_716_clock),
    .reset(q_716_reset),
    .io_enq_ready(q_716_io_enq_ready),
    .io_enq_valid(q_716_io_enq_valid),
    .io_enq_bits(q_716_io_enq_bits),
    .io_deq_ready(q_716_io_deq_ready),
    .io_deq_valid(q_716_io_deq_valid),
    .io_deq_bits(q_716_io_deq_bits)
  );
  Queue q_717 ( // @[Decoupled.scala 361:21]
    .clock(q_717_clock),
    .reset(q_717_reset),
    .io_enq_ready(q_717_io_enq_ready),
    .io_enq_valid(q_717_io_enq_valid),
    .io_enq_bits(q_717_io_enq_bits),
    .io_deq_ready(q_717_io_deq_ready),
    .io_deq_valid(q_717_io_deq_valid),
    .io_deq_bits(q_717_io_deq_bits)
  );
  Queue q_718 ( // @[Decoupled.scala 361:21]
    .clock(q_718_clock),
    .reset(q_718_reset),
    .io_enq_ready(q_718_io_enq_ready),
    .io_enq_valid(q_718_io_enq_valid),
    .io_enq_bits(q_718_io_enq_bits),
    .io_deq_ready(q_718_io_deq_ready),
    .io_deq_valid(q_718_io_deq_valid),
    .io_deq_bits(q_718_io_deq_bits)
  );
  Queue q_719 ( // @[Decoupled.scala 361:21]
    .clock(q_719_clock),
    .reset(q_719_reset),
    .io_enq_ready(q_719_io_enq_ready),
    .io_enq_valid(q_719_io_enq_valid),
    .io_enq_bits(q_719_io_enq_bits),
    .io_deq_ready(q_719_io_deq_ready),
    .io_deq_valid(q_719_io_deq_valid),
    .io_deq_bits(q_719_io_deq_bits)
  );
  Queue q_720 ( // @[Decoupled.scala 361:21]
    .clock(q_720_clock),
    .reset(q_720_reset),
    .io_enq_ready(q_720_io_enq_ready),
    .io_enq_valid(q_720_io_enq_valid),
    .io_enq_bits(q_720_io_enq_bits),
    .io_deq_ready(q_720_io_deq_ready),
    .io_deq_valid(q_720_io_deq_valid),
    .io_deq_bits(q_720_io_deq_bits)
  );
  Queue q_721 ( // @[Decoupled.scala 361:21]
    .clock(q_721_clock),
    .reset(q_721_reset),
    .io_enq_ready(q_721_io_enq_ready),
    .io_enq_valid(q_721_io_enq_valid),
    .io_enq_bits(q_721_io_enq_bits),
    .io_deq_ready(q_721_io_deq_ready),
    .io_deq_valid(q_721_io_deq_valid),
    .io_deq_bits(q_721_io_deq_bits)
  );
  Queue q_722 ( // @[Decoupled.scala 361:21]
    .clock(q_722_clock),
    .reset(q_722_reset),
    .io_enq_ready(q_722_io_enq_ready),
    .io_enq_valid(q_722_io_enq_valid),
    .io_enq_bits(q_722_io_enq_bits),
    .io_deq_ready(q_722_io_deq_ready),
    .io_deq_valid(q_722_io_deq_valid),
    .io_deq_bits(q_722_io_deq_bits)
  );
  Queue q_723 ( // @[Decoupled.scala 361:21]
    .clock(q_723_clock),
    .reset(q_723_reset),
    .io_enq_ready(q_723_io_enq_ready),
    .io_enq_valid(q_723_io_enq_valid),
    .io_enq_bits(q_723_io_enq_bits),
    .io_deq_ready(q_723_io_deq_ready),
    .io_deq_valid(q_723_io_deq_valid),
    .io_deq_bits(q_723_io_deq_bits)
  );
  Queue q_724 ( // @[Decoupled.scala 361:21]
    .clock(q_724_clock),
    .reset(q_724_reset),
    .io_enq_ready(q_724_io_enq_ready),
    .io_enq_valid(q_724_io_enq_valid),
    .io_enq_bits(q_724_io_enq_bits),
    .io_deq_ready(q_724_io_deq_ready),
    .io_deq_valid(q_724_io_deq_valid),
    .io_deq_bits(q_724_io_deq_bits)
  );
  Queue q_725 ( // @[Decoupled.scala 361:21]
    .clock(q_725_clock),
    .reset(q_725_reset),
    .io_enq_ready(q_725_io_enq_ready),
    .io_enq_valid(q_725_io_enq_valid),
    .io_enq_bits(q_725_io_enq_bits),
    .io_deq_ready(q_725_io_deq_ready),
    .io_deq_valid(q_725_io_deq_valid),
    .io_deq_bits(q_725_io_deq_bits)
  );
  Queue q_726 ( // @[Decoupled.scala 361:21]
    .clock(q_726_clock),
    .reset(q_726_reset),
    .io_enq_ready(q_726_io_enq_ready),
    .io_enq_valid(q_726_io_enq_valid),
    .io_enq_bits(q_726_io_enq_bits),
    .io_deq_ready(q_726_io_deq_ready),
    .io_deq_valid(q_726_io_deq_valid),
    .io_deq_bits(q_726_io_deq_bits)
  );
  Queue q_727 ( // @[Decoupled.scala 361:21]
    .clock(q_727_clock),
    .reset(q_727_reset),
    .io_enq_ready(q_727_io_enq_ready),
    .io_enq_valid(q_727_io_enq_valid),
    .io_enq_bits(q_727_io_enq_bits),
    .io_deq_ready(q_727_io_deq_ready),
    .io_deq_valid(q_727_io_deq_valid),
    .io_deq_bits(q_727_io_deq_bits)
  );
  Queue q_728 ( // @[Decoupled.scala 361:21]
    .clock(q_728_clock),
    .reset(q_728_reset),
    .io_enq_ready(q_728_io_enq_ready),
    .io_enq_valid(q_728_io_enq_valid),
    .io_enq_bits(q_728_io_enq_bits),
    .io_deq_ready(q_728_io_deq_ready),
    .io_deq_valid(q_728_io_deq_valid),
    .io_deq_bits(q_728_io_deq_bits)
  );
  Queue q_729 ( // @[Decoupled.scala 361:21]
    .clock(q_729_clock),
    .reset(q_729_reset),
    .io_enq_ready(q_729_io_enq_ready),
    .io_enq_valid(q_729_io_enq_valid),
    .io_enq_bits(q_729_io_enq_bits),
    .io_deq_ready(q_729_io_deq_ready),
    .io_deq_valid(q_729_io_deq_valid),
    .io_deq_bits(q_729_io_deq_bits)
  );
  Queue q_730 ( // @[Decoupled.scala 361:21]
    .clock(q_730_clock),
    .reset(q_730_reset),
    .io_enq_ready(q_730_io_enq_ready),
    .io_enq_valid(q_730_io_enq_valid),
    .io_enq_bits(q_730_io_enq_bits),
    .io_deq_ready(q_730_io_deq_ready),
    .io_deq_valid(q_730_io_deq_valid),
    .io_deq_bits(q_730_io_deq_bits)
  );
  Queue q_731 ( // @[Decoupled.scala 361:21]
    .clock(q_731_clock),
    .reset(q_731_reset),
    .io_enq_ready(q_731_io_enq_ready),
    .io_enq_valid(q_731_io_enq_valid),
    .io_enq_bits(q_731_io_enq_bits),
    .io_deq_ready(q_731_io_deq_ready),
    .io_deq_valid(q_731_io_deq_valid),
    .io_deq_bits(q_731_io_deq_bits)
  );
  Queue q_732 ( // @[Decoupled.scala 361:21]
    .clock(q_732_clock),
    .reset(q_732_reset),
    .io_enq_ready(q_732_io_enq_ready),
    .io_enq_valid(q_732_io_enq_valid),
    .io_enq_bits(q_732_io_enq_bits),
    .io_deq_ready(q_732_io_deq_ready),
    .io_deq_valid(q_732_io_deq_valid),
    .io_deq_bits(q_732_io_deq_bits)
  );
  Queue q_733 ( // @[Decoupled.scala 361:21]
    .clock(q_733_clock),
    .reset(q_733_reset),
    .io_enq_ready(q_733_io_enq_ready),
    .io_enq_valid(q_733_io_enq_valid),
    .io_enq_bits(q_733_io_enq_bits),
    .io_deq_ready(q_733_io_deq_ready),
    .io_deq_valid(q_733_io_deq_valid),
    .io_deq_bits(q_733_io_deq_bits)
  );
  Queue q_734 ( // @[Decoupled.scala 361:21]
    .clock(q_734_clock),
    .reset(q_734_reset),
    .io_enq_ready(q_734_io_enq_ready),
    .io_enq_valid(q_734_io_enq_valid),
    .io_enq_bits(q_734_io_enq_bits),
    .io_deq_ready(q_734_io_deq_ready),
    .io_deq_valid(q_734_io_deq_valid),
    .io_deq_bits(q_734_io_deq_bits)
  );
  Queue q_735 ( // @[Decoupled.scala 361:21]
    .clock(q_735_clock),
    .reset(q_735_reset),
    .io_enq_ready(q_735_io_enq_ready),
    .io_enq_valid(q_735_io_enq_valid),
    .io_enq_bits(q_735_io_enq_bits),
    .io_deq_ready(q_735_io_deq_ready),
    .io_deq_valid(q_735_io_deq_valid),
    .io_deq_bits(q_735_io_deq_bits)
  );
  Queue q_736 ( // @[Decoupled.scala 361:21]
    .clock(q_736_clock),
    .reset(q_736_reset),
    .io_enq_ready(q_736_io_enq_ready),
    .io_enq_valid(q_736_io_enq_valid),
    .io_enq_bits(q_736_io_enq_bits),
    .io_deq_ready(q_736_io_deq_ready),
    .io_deq_valid(q_736_io_deq_valid),
    .io_deq_bits(q_736_io_deq_bits)
  );
  Queue q_737 ( // @[Decoupled.scala 361:21]
    .clock(q_737_clock),
    .reset(q_737_reset),
    .io_enq_ready(q_737_io_enq_ready),
    .io_enq_valid(q_737_io_enq_valid),
    .io_enq_bits(q_737_io_enq_bits),
    .io_deq_ready(q_737_io_deq_ready),
    .io_deq_valid(q_737_io_deq_valid),
    .io_deq_bits(q_737_io_deq_bits)
  );
  Queue q_738 ( // @[Decoupled.scala 361:21]
    .clock(q_738_clock),
    .reset(q_738_reset),
    .io_enq_ready(q_738_io_enq_ready),
    .io_enq_valid(q_738_io_enq_valid),
    .io_enq_bits(q_738_io_enq_bits),
    .io_deq_ready(q_738_io_deq_ready),
    .io_deq_valid(q_738_io_deq_valid),
    .io_deq_bits(q_738_io_deq_bits)
  );
  Queue q_739 ( // @[Decoupled.scala 361:21]
    .clock(q_739_clock),
    .reset(q_739_reset),
    .io_enq_ready(q_739_io_enq_ready),
    .io_enq_valid(q_739_io_enq_valid),
    .io_enq_bits(q_739_io_enq_bits),
    .io_deq_ready(q_739_io_deq_ready),
    .io_deq_valid(q_739_io_deq_valid),
    .io_deq_bits(q_739_io_deq_bits)
  );
  Queue q_740 ( // @[Decoupled.scala 361:21]
    .clock(q_740_clock),
    .reset(q_740_reset),
    .io_enq_ready(q_740_io_enq_ready),
    .io_enq_valid(q_740_io_enq_valid),
    .io_enq_bits(q_740_io_enq_bits),
    .io_deq_ready(q_740_io_deq_ready),
    .io_deq_valid(q_740_io_deq_valid),
    .io_deq_bits(q_740_io_deq_bits)
  );
  Queue q_741 ( // @[Decoupled.scala 361:21]
    .clock(q_741_clock),
    .reset(q_741_reset),
    .io_enq_ready(q_741_io_enq_ready),
    .io_enq_valid(q_741_io_enq_valid),
    .io_enq_bits(q_741_io_enq_bits),
    .io_deq_ready(q_741_io_deq_ready),
    .io_deq_valid(q_741_io_deq_valid),
    .io_deq_bits(q_741_io_deq_bits)
  );
  Queue q_742 ( // @[Decoupled.scala 361:21]
    .clock(q_742_clock),
    .reset(q_742_reset),
    .io_enq_ready(q_742_io_enq_ready),
    .io_enq_valid(q_742_io_enq_valid),
    .io_enq_bits(q_742_io_enq_bits),
    .io_deq_ready(q_742_io_deq_ready),
    .io_deq_valid(q_742_io_deq_valid),
    .io_deq_bits(q_742_io_deq_bits)
  );
  Queue q_743 ( // @[Decoupled.scala 361:21]
    .clock(q_743_clock),
    .reset(q_743_reset),
    .io_enq_ready(q_743_io_enq_ready),
    .io_enq_valid(q_743_io_enq_valid),
    .io_enq_bits(q_743_io_enq_bits),
    .io_deq_ready(q_743_io_deq_ready),
    .io_deq_valid(q_743_io_deq_valid),
    .io_deq_bits(q_743_io_deq_bits)
  );
  Queue q_744 ( // @[Decoupled.scala 361:21]
    .clock(q_744_clock),
    .reset(q_744_reset),
    .io_enq_ready(q_744_io_enq_ready),
    .io_enq_valid(q_744_io_enq_valid),
    .io_enq_bits(q_744_io_enq_bits),
    .io_deq_ready(q_744_io_deq_ready),
    .io_deq_valid(q_744_io_deq_valid),
    .io_deq_bits(q_744_io_deq_bits)
  );
  Queue q_745 ( // @[Decoupled.scala 361:21]
    .clock(q_745_clock),
    .reset(q_745_reset),
    .io_enq_ready(q_745_io_enq_ready),
    .io_enq_valid(q_745_io_enq_valid),
    .io_enq_bits(q_745_io_enq_bits),
    .io_deq_ready(q_745_io_deq_ready),
    .io_deq_valid(q_745_io_deq_valid),
    .io_deq_bits(q_745_io_deq_bits)
  );
  Queue q_746 ( // @[Decoupled.scala 361:21]
    .clock(q_746_clock),
    .reset(q_746_reset),
    .io_enq_ready(q_746_io_enq_ready),
    .io_enq_valid(q_746_io_enq_valid),
    .io_enq_bits(q_746_io_enq_bits),
    .io_deq_ready(q_746_io_deq_ready),
    .io_deq_valid(q_746_io_deq_valid),
    .io_deq_bits(q_746_io_deq_bits)
  );
  Queue q_747 ( // @[Decoupled.scala 361:21]
    .clock(q_747_clock),
    .reset(q_747_reset),
    .io_enq_ready(q_747_io_enq_ready),
    .io_enq_valid(q_747_io_enq_valid),
    .io_enq_bits(q_747_io_enq_bits),
    .io_deq_ready(q_747_io_deq_ready),
    .io_deq_valid(q_747_io_deq_valid),
    .io_deq_bits(q_747_io_deq_bits)
  );
  Queue q_748 ( // @[Decoupled.scala 361:21]
    .clock(q_748_clock),
    .reset(q_748_reset),
    .io_enq_ready(q_748_io_enq_ready),
    .io_enq_valid(q_748_io_enq_valid),
    .io_enq_bits(q_748_io_enq_bits),
    .io_deq_ready(q_748_io_deq_ready),
    .io_deq_valid(q_748_io_deq_valid),
    .io_deq_bits(q_748_io_deq_bits)
  );
  Queue q_749 ( // @[Decoupled.scala 361:21]
    .clock(q_749_clock),
    .reset(q_749_reset),
    .io_enq_ready(q_749_io_enq_ready),
    .io_enq_valid(q_749_io_enq_valid),
    .io_enq_bits(q_749_io_enq_bits),
    .io_deq_ready(q_749_io_deq_ready),
    .io_deq_valid(q_749_io_deq_valid),
    .io_deq_bits(q_749_io_deq_bits)
  );
  Queue q_750 ( // @[Decoupled.scala 361:21]
    .clock(q_750_clock),
    .reset(q_750_reset),
    .io_enq_ready(q_750_io_enq_ready),
    .io_enq_valid(q_750_io_enq_valid),
    .io_enq_bits(q_750_io_enq_bits),
    .io_deq_ready(q_750_io_deq_ready),
    .io_deq_valid(q_750_io_deq_valid),
    .io_deq_bits(q_750_io_deq_bits)
  );
  Queue q_751 ( // @[Decoupled.scala 361:21]
    .clock(q_751_clock),
    .reset(q_751_reset),
    .io_enq_ready(q_751_io_enq_ready),
    .io_enq_valid(q_751_io_enq_valid),
    .io_enq_bits(q_751_io_enq_bits),
    .io_deq_ready(q_751_io_deq_ready),
    .io_deq_valid(q_751_io_deq_valid),
    .io_deq_bits(q_751_io_deq_bits)
  );
  Queue q_752 ( // @[Decoupled.scala 361:21]
    .clock(q_752_clock),
    .reset(q_752_reset),
    .io_enq_ready(q_752_io_enq_ready),
    .io_enq_valid(q_752_io_enq_valid),
    .io_enq_bits(q_752_io_enq_bits),
    .io_deq_ready(q_752_io_deq_ready),
    .io_deq_valid(q_752_io_deq_valid),
    .io_deq_bits(q_752_io_deq_bits)
  );
  Queue q_753 ( // @[Decoupled.scala 361:21]
    .clock(q_753_clock),
    .reset(q_753_reset),
    .io_enq_ready(q_753_io_enq_ready),
    .io_enq_valid(q_753_io_enq_valid),
    .io_enq_bits(q_753_io_enq_bits),
    .io_deq_ready(q_753_io_deq_ready),
    .io_deq_valid(q_753_io_deq_valid),
    .io_deq_bits(q_753_io_deq_bits)
  );
  Queue q_754 ( // @[Decoupled.scala 361:21]
    .clock(q_754_clock),
    .reset(q_754_reset),
    .io_enq_ready(q_754_io_enq_ready),
    .io_enq_valid(q_754_io_enq_valid),
    .io_enq_bits(q_754_io_enq_bits),
    .io_deq_ready(q_754_io_deq_ready),
    .io_deq_valid(q_754_io_deq_valid),
    .io_deq_bits(q_754_io_deq_bits)
  );
  Queue q_755 ( // @[Decoupled.scala 361:21]
    .clock(q_755_clock),
    .reset(q_755_reset),
    .io_enq_ready(q_755_io_enq_ready),
    .io_enq_valid(q_755_io_enq_valid),
    .io_enq_bits(q_755_io_enq_bits),
    .io_deq_ready(q_755_io_deq_ready),
    .io_deq_valid(q_755_io_deq_valid),
    .io_deq_bits(q_755_io_deq_bits)
  );
  Queue q_756 ( // @[Decoupled.scala 361:21]
    .clock(q_756_clock),
    .reset(q_756_reset),
    .io_enq_ready(q_756_io_enq_ready),
    .io_enq_valid(q_756_io_enq_valid),
    .io_enq_bits(q_756_io_enq_bits),
    .io_deq_ready(q_756_io_deq_ready),
    .io_deq_valid(q_756_io_deq_valid),
    .io_deq_bits(q_756_io_deq_bits)
  );
  Queue q_757 ( // @[Decoupled.scala 361:21]
    .clock(q_757_clock),
    .reset(q_757_reset),
    .io_enq_ready(q_757_io_enq_ready),
    .io_enq_valid(q_757_io_enq_valid),
    .io_enq_bits(q_757_io_enq_bits),
    .io_deq_ready(q_757_io_deq_ready),
    .io_deq_valid(q_757_io_deq_valid),
    .io_deq_bits(q_757_io_deq_bits)
  );
  Queue q_758 ( // @[Decoupled.scala 361:21]
    .clock(q_758_clock),
    .reset(q_758_reset),
    .io_enq_ready(q_758_io_enq_ready),
    .io_enq_valid(q_758_io_enq_valid),
    .io_enq_bits(q_758_io_enq_bits),
    .io_deq_ready(q_758_io_deq_ready),
    .io_deq_valid(q_758_io_deq_valid),
    .io_deq_bits(q_758_io_deq_bits)
  );
  Queue q_759 ( // @[Decoupled.scala 361:21]
    .clock(q_759_clock),
    .reset(q_759_reset),
    .io_enq_ready(q_759_io_enq_ready),
    .io_enq_valid(q_759_io_enq_valid),
    .io_enq_bits(q_759_io_enq_bits),
    .io_deq_ready(q_759_io_deq_ready),
    .io_deq_valid(q_759_io_deq_valid),
    .io_deq_bits(q_759_io_deq_bits)
  );
  Queue q_760 ( // @[Decoupled.scala 361:21]
    .clock(q_760_clock),
    .reset(q_760_reset),
    .io_enq_ready(q_760_io_enq_ready),
    .io_enq_valid(q_760_io_enq_valid),
    .io_enq_bits(q_760_io_enq_bits),
    .io_deq_ready(q_760_io_deq_ready),
    .io_deq_valid(q_760_io_deq_valid),
    .io_deq_bits(q_760_io_deq_bits)
  );
  Queue q_761 ( // @[Decoupled.scala 361:21]
    .clock(q_761_clock),
    .reset(q_761_reset),
    .io_enq_ready(q_761_io_enq_ready),
    .io_enq_valid(q_761_io_enq_valid),
    .io_enq_bits(q_761_io_enq_bits),
    .io_deq_ready(q_761_io_deq_ready),
    .io_deq_valid(q_761_io_deq_valid),
    .io_deq_bits(q_761_io_deq_bits)
  );
  Queue q_762 ( // @[Decoupled.scala 361:21]
    .clock(q_762_clock),
    .reset(q_762_reset),
    .io_enq_ready(q_762_io_enq_ready),
    .io_enq_valid(q_762_io_enq_valid),
    .io_enq_bits(q_762_io_enq_bits),
    .io_deq_ready(q_762_io_deq_ready),
    .io_deq_valid(q_762_io_deq_valid),
    .io_deq_bits(q_762_io_deq_bits)
  );
  Queue q_763 ( // @[Decoupled.scala 361:21]
    .clock(q_763_clock),
    .reset(q_763_reset),
    .io_enq_ready(q_763_io_enq_ready),
    .io_enq_valid(q_763_io_enq_valid),
    .io_enq_bits(q_763_io_enq_bits),
    .io_deq_ready(q_763_io_deq_ready),
    .io_deq_valid(q_763_io_deq_valid),
    .io_deq_bits(q_763_io_deq_bits)
  );
  Queue q_764 ( // @[Decoupled.scala 361:21]
    .clock(q_764_clock),
    .reset(q_764_reset),
    .io_enq_ready(q_764_io_enq_ready),
    .io_enq_valid(q_764_io_enq_valid),
    .io_enq_bits(q_764_io_enq_bits),
    .io_deq_ready(q_764_io_deq_ready),
    .io_deq_valid(q_764_io_deq_valid),
    .io_deq_bits(q_764_io_deq_bits)
  );
  Queue q_765 ( // @[Decoupled.scala 361:21]
    .clock(q_765_clock),
    .reset(q_765_reset),
    .io_enq_ready(q_765_io_enq_ready),
    .io_enq_valid(q_765_io_enq_valid),
    .io_enq_bits(q_765_io_enq_bits),
    .io_deq_ready(q_765_io_deq_ready),
    .io_deq_valid(q_765_io_deq_valid),
    .io_deq_bits(q_765_io_deq_bits)
  );
  Queue q_766 ( // @[Decoupled.scala 361:21]
    .clock(q_766_clock),
    .reset(q_766_reset),
    .io_enq_ready(q_766_io_enq_ready),
    .io_enq_valid(q_766_io_enq_valid),
    .io_enq_bits(q_766_io_enq_bits),
    .io_deq_ready(q_766_io_deq_ready),
    .io_deq_valid(q_766_io_deq_valid),
    .io_deq_bits(q_766_io_deq_bits)
  );
  Queue q_767 ( // @[Decoupled.scala 361:21]
    .clock(q_767_clock),
    .reset(q_767_reset),
    .io_enq_ready(q_767_io_enq_ready),
    .io_enq_valid(q_767_io_enq_valid),
    .io_enq_bits(q_767_io_enq_bits),
    .io_deq_ready(q_767_io_deq_ready),
    .io_deq_valid(q_767_io_deq_valid),
    .io_deq_bits(q_767_io_deq_bits)
  );
  assign io_weight_in_0_ready = q_240_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_weight_in_1_ready = q_241_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_weight_in_2_ready = q_242_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_weight_in_3_ready = q_243_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_weight_in_4_ready = q_244_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_weight_in_5_ready = q_245_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_weight_in_6_ready = q_246_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_weight_in_7_ready = q_247_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_weight_in_8_ready = q_248_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_weight_in_9_ready = q_249_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_weight_in_10_ready = q_250_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_weight_in_11_ready = q_251_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_weight_in_12_ready = q_252_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_weight_in_13_ready = q_253_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_weight_in_14_ready = q_254_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_weight_in_15_ready = q_255_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_in_0_ready = q_496_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_in_1_ready = q_497_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_in_2_ready = q_498_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_in_3_ready = q_499_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_in_4_ready = q_500_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_in_5_ready = q_501_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_in_6_ready = q_502_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_in_7_ready = q_503_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_in_8_ready = q_504_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_in_9_ready = q_505_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_in_10_ready = q_506_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_in_11_ready = q_507_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_in_12_ready = q_508_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_in_13_ready = q_509_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_in_14_ready = q_510_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_in_15_ready = q_511_io_enq_ready; // @[Decoupled.scala 365:17]
  assign io_value_out_0_0_valid = q_512_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_0_0_bits = q_512_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_0_1_valid = q_513_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_0_1_bits = q_513_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_0_2_valid = q_514_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_0_2_bits = q_514_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_0_3_valid = q_515_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_0_3_bits = q_515_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_0_4_valid = q_516_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_0_4_bits = q_516_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_0_5_valid = q_517_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_0_5_bits = q_517_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_0_6_valid = q_518_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_0_6_bits = q_518_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_0_7_valid = q_519_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_0_7_bits = q_519_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_0_8_valid = q_520_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_0_8_bits = q_520_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_0_9_valid = q_521_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_0_9_bits = q_521_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_0_10_valid = q_522_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_0_10_bits = q_522_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_0_11_valid = q_523_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_0_11_bits = q_523_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_0_12_valid = q_524_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_0_12_bits = q_524_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_0_13_valid = q_525_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_0_13_bits = q_525_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_0_14_valid = q_526_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_0_14_bits = q_526_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_0_15_valid = q_527_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_0_15_bits = q_527_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_1_0_valid = q_528_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_1_0_bits = q_528_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_1_1_valid = q_529_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_1_1_bits = q_529_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_1_2_valid = q_530_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_1_2_bits = q_530_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_1_3_valid = q_531_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_1_3_bits = q_531_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_1_4_valid = q_532_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_1_4_bits = q_532_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_1_5_valid = q_533_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_1_5_bits = q_533_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_1_6_valid = q_534_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_1_6_bits = q_534_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_1_7_valid = q_535_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_1_7_bits = q_535_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_1_8_valid = q_536_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_1_8_bits = q_536_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_1_9_valid = q_537_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_1_9_bits = q_537_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_1_10_valid = q_538_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_1_10_bits = q_538_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_1_11_valid = q_539_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_1_11_bits = q_539_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_1_12_valid = q_540_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_1_12_bits = q_540_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_1_13_valid = q_541_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_1_13_bits = q_541_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_1_14_valid = q_542_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_1_14_bits = q_542_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_1_15_valid = q_543_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_1_15_bits = q_543_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_2_0_valid = q_544_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_2_0_bits = q_544_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_2_1_valid = q_545_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_2_1_bits = q_545_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_2_2_valid = q_546_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_2_2_bits = q_546_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_2_3_valid = q_547_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_2_3_bits = q_547_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_2_4_valid = q_548_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_2_4_bits = q_548_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_2_5_valid = q_549_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_2_5_bits = q_549_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_2_6_valid = q_550_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_2_6_bits = q_550_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_2_7_valid = q_551_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_2_7_bits = q_551_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_2_8_valid = q_552_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_2_8_bits = q_552_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_2_9_valid = q_553_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_2_9_bits = q_553_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_2_10_valid = q_554_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_2_10_bits = q_554_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_2_11_valid = q_555_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_2_11_bits = q_555_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_2_12_valid = q_556_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_2_12_bits = q_556_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_2_13_valid = q_557_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_2_13_bits = q_557_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_2_14_valid = q_558_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_2_14_bits = q_558_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_2_15_valid = q_559_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_2_15_bits = q_559_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_3_0_valid = q_560_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_3_0_bits = q_560_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_3_1_valid = q_561_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_3_1_bits = q_561_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_3_2_valid = q_562_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_3_2_bits = q_562_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_3_3_valid = q_563_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_3_3_bits = q_563_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_3_4_valid = q_564_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_3_4_bits = q_564_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_3_5_valid = q_565_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_3_5_bits = q_565_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_3_6_valid = q_566_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_3_6_bits = q_566_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_3_7_valid = q_567_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_3_7_bits = q_567_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_3_8_valid = q_568_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_3_8_bits = q_568_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_3_9_valid = q_569_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_3_9_bits = q_569_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_3_10_valid = q_570_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_3_10_bits = q_570_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_3_11_valid = q_571_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_3_11_bits = q_571_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_3_12_valid = q_572_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_3_12_bits = q_572_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_3_13_valid = q_573_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_3_13_bits = q_573_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_3_14_valid = q_574_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_3_14_bits = q_574_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_3_15_valid = q_575_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_3_15_bits = q_575_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_4_0_valid = q_576_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_4_0_bits = q_576_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_4_1_valid = q_577_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_4_1_bits = q_577_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_4_2_valid = q_578_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_4_2_bits = q_578_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_4_3_valid = q_579_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_4_3_bits = q_579_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_4_4_valid = q_580_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_4_4_bits = q_580_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_4_5_valid = q_581_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_4_5_bits = q_581_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_4_6_valid = q_582_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_4_6_bits = q_582_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_4_7_valid = q_583_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_4_7_bits = q_583_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_4_8_valid = q_584_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_4_8_bits = q_584_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_4_9_valid = q_585_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_4_9_bits = q_585_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_4_10_valid = q_586_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_4_10_bits = q_586_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_4_11_valid = q_587_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_4_11_bits = q_587_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_4_12_valid = q_588_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_4_12_bits = q_588_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_4_13_valid = q_589_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_4_13_bits = q_589_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_4_14_valid = q_590_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_4_14_bits = q_590_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_4_15_valid = q_591_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_4_15_bits = q_591_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_5_0_valid = q_592_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_5_0_bits = q_592_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_5_1_valid = q_593_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_5_1_bits = q_593_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_5_2_valid = q_594_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_5_2_bits = q_594_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_5_3_valid = q_595_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_5_3_bits = q_595_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_5_4_valid = q_596_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_5_4_bits = q_596_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_5_5_valid = q_597_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_5_5_bits = q_597_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_5_6_valid = q_598_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_5_6_bits = q_598_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_5_7_valid = q_599_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_5_7_bits = q_599_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_5_8_valid = q_600_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_5_8_bits = q_600_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_5_9_valid = q_601_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_5_9_bits = q_601_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_5_10_valid = q_602_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_5_10_bits = q_602_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_5_11_valid = q_603_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_5_11_bits = q_603_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_5_12_valid = q_604_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_5_12_bits = q_604_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_5_13_valid = q_605_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_5_13_bits = q_605_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_5_14_valid = q_606_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_5_14_bits = q_606_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_5_15_valid = q_607_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_5_15_bits = q_607_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_6_0_valid = q_608_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_6_0_bits = q_608_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_6_1_valid = q_609_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_6_1_bits = q_609_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_6_2_valid = q_610_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_6_2_bits = q_610_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_6_3_valid = q_611_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_6_3_bits = q_611_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_6_4_valid = q_612_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_6_4_bits = q_612_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_6_5_valid = q_613_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_6_5_bits = q_613_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_6_6_valid = q_614_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_6_6_bits = q_614_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_6_7_valid = q_615_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_6_7_bits = q_615_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_6_8_valid = q_616_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_6_8_bits = q_616_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_6_9_valid = q_617_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_6_9_bits = q_617_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_6_10_valid = q_618_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_6_10_bits = q_618_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_6_11_valid = q_619_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_6_11_bits = q_619_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_6_12_valid = q_620_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_6_12_bits = q_620_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_6_13_valid = q_621_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_6_13_bits = q_621_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_6_14_valid = q_622_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_6_14_bits = q_622_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_6_15_valid = q_623_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_6_15_bits = q_623_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_7_0_valid = q_624_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_7_0_bits = q_624_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_7_1_valid = q_625_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_7_1_bits = q_625_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_7_2_valid = q_626_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_7_2_bits = q_626_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_7_3_valid = q_627_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_7_3_bits = q_627_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_7_4_valid = q_628_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_7_4_bits = q_628_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_7_5_valid = q_629_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_7_5_bits = q_629_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_7_6_valid = q_630_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_7_6_bits = q_630_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_7_7_valid = q_631_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_7_7_bits = q_631_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_7_8_valid = q_632_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_7_8_bits = q_632_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_7_9_valid = q_633_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_7_9_bits = q_633_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_7_10_valid = q_634_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_7_10_bits = q_634_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_7_11_valid = q_635_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_7_11_bits = q_635_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_7_12_valid = q_636_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_7_12_bits = q_636_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_7_13_valid = q_637_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_7_13_bits = q_637_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_7_14_valid = q_638_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_7_14_bits = q_638_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_7_15_valid = q_639_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_7_15_bits = q_639_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_8_0_valid = q_640_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_8_0_bits = q_640_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_8_1_valid = q_641_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_8_1_bits = q_641_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_8_2_valid = q_642_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_8_2_bits = q_642_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_8_3_valid = q_643_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_8_3_bits = q_643_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_8_4_valid = q_644_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_8_4_bits = q_644_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_8_5_valid = q_645_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_8_5_bits = q_645_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_8_6_valid = q_646_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_8_6_bits = q_646_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_8_7_valid = q_647_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_8_7_bits = q_647_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_8_8_valid = q_648_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_8_8_bits = q_648_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_8_9_valid = q_649_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_8_9_bits = q_649_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_8_10_valid = q_650_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_8_10_bits = q_650_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_8_11_valid = q_651_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_8_11_bits = q_651_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_8_12_valid = q_652_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_8_12_bits = q_652_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_8_13_valid = q_653_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_8_13_bits = q_653_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_8_14_valid = q_654_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_8_14_bits = q_654_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_8_15_valid = q_655_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_8_15_bits = q_655_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_9_0_valid = q_656_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_9_0_bits = q_656_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_9_1_valid = q_657_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_9_1_bits = q_657_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_9_2_valid = q_658_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_9_2_bits = q_658_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_9_3_valid = q_659_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_9_3_bits = q_659_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_9_4_valid = q_660_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_9_4_bits = q_660_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_9_5_valid = q_661_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_9_5_bits = q_661_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_9_6_valid = q_662_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_9_6_bits = q_662_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_9_7_valid = q_663_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_9_7_bits = q_663_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_9_8_valid = q_664_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_9_8_bits = q_664_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_9_9_valid = q_665_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_9_9_bits = q_665_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_9_10_valid = q_666_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_9_10_bits = q_666_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_9_11_valid = q_667_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_9_11_bits = q_667_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_9_12_valid = q_668_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_9_12_bits = q_668_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_9_13_valid = q_669_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_9_13_bits = q_669_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_9_14_valid = q_670_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_9_14_bits = q_670_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_9_15_valid = q_671_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_9_15_bits = q_671_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_10_0_valid = q_672_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_10_0_bits = q_672_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_10_1_valid = q_673_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_10_1_bits = q_673_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_10_2_valid = q_674_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_10_2_bits = q_674_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_10_3_valid = q_675_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_10_3_bits = q_675_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_10_4_valid = q_676_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_10_4_bits = q_676_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_10_5_valid = q_677_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_10_5_bits = q_677_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_10_6_valid = q_678_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_10_6_bits = q_678_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_10_7_valid = q_679_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_10_7_bits = q_679_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_10_8_valid = q_680_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_10_8_bits = q_680_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_10_9_valid = q_681_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_10_9_bits = q_681_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_10_10_valid = q_682_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_10_10_bits = q_682_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_10_11_valid = q_683_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_10_11_bits = q_683_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_10_12_valid = q_684_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_10_12_bits = q_684_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_10_13_valid = q_685_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_10_13_bits = q_685_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_10_14_valid = q_686_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_10_14_bits = q_686_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_10_15_valid = q_687_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_10_15_bits = q_687_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_11_0_valid = q_688_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_11_0_bits = q_688_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_11_1_valid = q_689_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_11_1_bits = q_689_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_11_2_valid = q_690_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_11_2_bits = q_690_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_11_3_valid = q_691_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_11_3_bits = q_691_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_11_4_valid = q_692_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_11_4_bits = q_692_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_11_5_valid = q_693_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_11_5_bits = q_693_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_11_6_valid = q_694_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_11_6_bits = q_694_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_11_7_valid = q_695_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_11_7_bits = q_695_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_11_8_valid = q_696_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_11_8_bits = q_696_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_11_9_valid = q_697_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_11_9_bits = q_697_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_11_10_valid = q_698_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_11_10_bits = q_698_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_11_11_valid = q_699_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_11_11_bits = q_699_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_11_12_valid = q_700_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_11_12_bits = q_700_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_11_13_valid = q_701_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_11_13_bits = q_701_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_11_14_valid = q_702_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_11_14_bits = q_702_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_11_15_valid = q_703_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_11_15_bits = q_703_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_12_0_valid = q_704_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_12_0_bits = q_704_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_12_1_valid = q_705_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_12_1_bits = q_705_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_12_2_valid = q_706_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_12_2_bits = q_706_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_12_3_valid = q_707_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_12_3_bits = q_707_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_12_4_valid = q_708_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_12_4_bits = q_708_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_12_5_valid = q_709_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_12_5_bits = q_709_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_12_6_valid = q_710_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_12_6_bits = q_710_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_12_7_valid = q_711_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_12_7_bits = q_711_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_12_8_valid = q_712_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_12_8_bits = q_712_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_12_9_valid = q_713_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_12_9_bits = q_713_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_12_10_valid = q_714_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_12_10_bits = q_714_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_12_11_valid = q_715_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_12_11_bits = q_715_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_12_12_valid = q_716_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_12_12_bits = q_716_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_12_13_valid = q_717_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_12_13_bits = q_717_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_12_14_valid = q_718_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_12_14_bits = q_718_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_12_15_valid = q_719_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_12_15_bits = q_719_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_13_0_valid = q_720_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_13_0_bits = q_720_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_13_1_valid = q_721_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_13_1_bits = q_721_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_13_2_valid = q_722_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_13_2_bits = q_722_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_13_3_valid = q_723_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_13_3_bits = q_723_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_13_4_valid = q_724_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_13_4_bits = q_724_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_13_5_valid = q_725_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_13_5_bits = q_725_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_13_6_valid = q_726_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_13_6_bits = q_726_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_13_7_valid = q_727_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_13_7_bits = q_727_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_13_8_valid = q_728_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_13_8_bits = q_728_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_13_9_valid = q_729_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_13_9_bits = q_729_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_13_10_valid = q_730_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_13_10_bits = q_730_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_13_11_valid = q_731_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_13_11_bits = q_731_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_13_12_valid = q_732_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_13_12_bits = q_732_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_13_13_valid = q_733_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_13_13_bits = q_733_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_13_14_valid = q_734_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_13_14_bits = q_734_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_13_15_valid = q_735_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_13_15_bits = q_735_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_14_0_valid = q_736_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_14_0_bits = q_736_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_14_1_valid = q_737_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_14_1_bits = q_737_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_14_2_valid = q_738_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_14_2_bits = q_738_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_14_3_valid = q_739_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_14_3_bits = q_739_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_14_4_valid = q_740_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_14_4_bits = q_740_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_14_5_valid = q_741_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_14_5_bits = q_741_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_14_6_valid = q_742_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_14_6_bits = q_742_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_14_7_valid = q_743_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_14_7_bits = q_743_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_14_8_valid = q_744_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_14_8_bits = q_744_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_14_9_valid = q_745_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_14_9_bits = q_745_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_14_10_valid = q_746_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_14_10_bits = q_746_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_14_11_valid = q_747_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_14_11_bits = q_747_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_14_12_valid = q_748_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_14_12_bits = q_748_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_14_13_valid = q_749_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_14_13_bits = q_749_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_14_14_valid = q_750_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_14_14_bits = q_750_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_14_15_valid = q_751_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_14_15_bits = q_751_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_15_0_valid = q_752_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_15_0_bits = q_752_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_15_1_valid = q_753_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_15_1_bits = q_753_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_15_2_valid = q_754_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_15_2_bits = q_754_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_15_3_valid = q_755_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_15_3_bits = q_755_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_15_4_valid = q_756_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_15_4_bits = q_756_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_15_5_valid = q_757_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_15_5_bits = q_757_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_15_6_valid = q_758_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_15_6_bits = q_758_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_15_7_valid = q_759_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_15_7_bits = q_759_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_15_8_valid = q_760_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_15_8_bits = q_760_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_15_9_valid = q_761_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_15_9_bits = q_761_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_15_10_valid = q_762_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_15_10_bits = q_762_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_15_11_valid = q_763_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_15_11_bits = q_763_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_15_12_valid = q_764_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_15_12_bits = q_764_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_15_13_valid = q_765_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_15_13_bits = q_765_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_15_14_valid = q_766_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_15_14_bits = q_766_io_deq_bits; // @[Stab.scala 104:101]
  assign io_value_out_15_15_valid = q_767_io_deq_valid; // @[Stab.scala 104:101]
  assign io_value_out_15_15_bits = q_767_io_deq_bits; // @[Stab.scala 104:101]
  assign cols_0_0_clock = clock;
  assign cols_0_0_reset = reset;
  assign cols_0_0_io_left_in_valid = q_496_io_deq_valid; // @[Stab.scala 100:101]
  assign cols_0_0_io_left_in_bits = q_496_io_deq_bits; // @[Stab.scala 100:101]
  assign cols_0_0_io_top_in_valid = q_240_io_deq_valid; // @[Stab.scala 93:102]
  assign cols_0_0_io_top_in_bits = q_240_io_deq_bits; // @[Stab.scala 93:102]
  assign cols_0_0_io_sum_ready = q_512_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_0_io_right_out_ready = q_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_0_io_bottom_out_ready = q_256_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_0_clock = clock;
  assign cols_1_0_reset = reset;
  assign cols_1_0_io_left_in_valid = q_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_1_0_io_left_in_bits = q_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_1_0_io_top_in_valid = q_241_io_deq_valid; // @[Stab.scala 93:102]
  assign cols_1_0_io_top_in_bits = q_241_io_deq_bits; // @[Stab.scala 93:102]
  assign cols_1_0_io_sum_ready = q_513_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_0_io_right_out_ready = q_1_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_0_io_bottom_out_ready = q_271_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_0_clock = clock;
  assign cols_2_0_reset = reset;
  assign cols_2_0_io_left_in_valid = q_1_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_2_0_io_left_in_bits = q_1_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_2_0_io_top_in_valid = q_242_io_deq_valid; // @[Stab.scala 93:102]
  assign cols_2_0_io_top_in_bits = q_242_io_deq_bits; // @[Stab.scala 93:102]
  assign cols_2_0_io_sum_ready = q_514_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_0_io_right_out_ready = q_2_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_0_io_bottom_out_ready = q_286_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_0_clock = clock;
  assign cols_3_0_reset = reset;
  assign cols_3_0_io_left_in_valid = q_2_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_3_0_io_left_in_bits = q_2_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_3_0_io_top_in_valid = q_243_io_deq_valid; // @[Stab.scala 93:102]
  assign cols_3_0_io_top_in_bits = q_243_io_deq_bits; // @[Stab.scala 93:102]
  assign cols_3_0_io_sum_ready = q_515_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_0_io_right_out_ready = q_3_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_0_io_bottom_out_ready = q_301_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_0_clock = clock;
  assign cols_4_0_reset = reset;
  assign cols_4_0_io_left_in_valid = q_3_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_4_0_io_left_in_bits = q_3_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_4_0_io_top_in_valid = q_244_io_deq_valid; // @[Stab.scala 93:102]
  assign cols_4_0_io_top_in_bits = q_244_io_deq_bits; // @[Stab.scala 93:102]
  assign cols_4_0_io_sum_ready = q_516_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_0_io_right_out_ready = q_4_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_0_io_bottom_out_ready = q_316_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_0_clock = clock;
  assign cols_5_0_reset = reset;
  assign cols_5_0_io_left_in_valid = q_4_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_5_0_io_left_in_bits = q_4_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_5_0_io_top_in_valid = q_245_io_deq_valid; // @[Stab.scala 93:102]
  assign cols_5_0_io_top_in_bits = q_245_io_deq_bits; // @[Stab.scala 93:102]
  assign cols_5_0_io_sum_ready = q_517_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_0_io_right_out_ready = q_5_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_0_io_bottom_out_ready = q_331_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_0_clock = clock;
  assign cols_6_0_reset = reset;
  assign cols_6_0_io_left_in_valid = q_5_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_6_0_io_left_in_bits = q_5_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_6_0_io_top_in_valid = q_246_io_deq_valid; // @[Stab.scala 93:102]
  assign cols_6_0_io_top_in_bits = q_246_io_deq_bits; // @[Stab.scala 93:102]
  assign cols_6_0_io_sum_ready = q_518_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_0_io_right_out_ready = q_6_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_0_io_bottom_out_ready = q_346_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_0_clock = clock;
  assign cols_7_0_reset = reset;
  assign cols_7_0_io_left_in_valid = q_6_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_7_0_io_left_in_bits = q_6_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_7_0_io_top_in_valid = q_247_io_deq_valid; // @[Stab.scala 93:102]
  assign cols_7_0_io_top_in_bits = q_247_io_deq_bits; // @[Stab.scala 93:102]
  assign cols_7_0_io_sum_ready = q_519_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_0_io_right_out_ready = q_7_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_0_io_bottom_out_ready = q_361_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_0_clock = clock;
  assign cols_8_0_reset = reset;
  assign cols_8_0_io_left_in_valid = q_7_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_8_0_io_left_in_bits = q_7_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_8_0_io_top_in_valid = q_248_io_deq_valid; // @[Stab.scala 93:102]
  assign cols_8_0_io_top_in_bits = q_248_io_deq_bits; // @[Stab.scala 93:102]
  assign cols_8_0_io_sum_ready = q_520_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_0_io_right_out_ready = q_8_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_0_io_bottom_out_ready = q_376_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_0_clock = clock;
  assign cols_9_0_reset = reset;
  assign cols_9_0_io_left_in_valid = q_8_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_9_0_io_left_in_bits = q_8_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_9_0_io_top_in_valid = q_249_io_deq_valid; // @[Stab.scala 93:102]
  assign cols_9_0_io_top_in_bits = q_249_io_deq_bits; // @[Stab.scala 93:102]
  assign cols_9_0_io_sum_ready = q_521_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_0_io_right_out_ready = q_9_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_0_io_bottom_out_ready = q_391_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_0_clock = clock;
  assign cols_10_0_reset = reset;
  assign cols_10_0_io_left_in_valid = q_9_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_10_0_io_left_in_bits = q_9_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_10_0_io_top_in_valid = q_250_io_deq_valid; // @[Stab.scala 93:102]
  assign cols_10_0_io_top_in_bits = q_250_io_deq_bits; // @[Stab.scala 93:102]
  assign cols_10_0_io_sum_ready = q_522_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_0_io_right_out_ready = q_10_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_0_io_bottom_out_ready = q_406_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_0_clock = clock;
  assign cols_11_0_reset = reset;
  assign cols_11_0_io_left_in_valid = q_10_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_11_0_io_left_in_bits = q_10_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_11_0_io_top_in_valid = q_251_io_deq_valid; // @[Stab.scala 93:102]
  assign cols_11_0_io_top_in_bits = q_251_io_deq_bits; // @[Stab.scala 93:102]
  assign cols_11_0_io_sum_ready = q_523_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_0_io_right_out_ready = q_11_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_0_io_bottom_out_ready = q_421_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_0_clock = clock;
  assign cols_12_0_reset = reset;
  assign cols_12_0_io_left_in_valid = q_11_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_12_0_io_left_in_bits = q_11_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_12_0_io_top_in_valid = q_252_io_deq_valid; // @[Stab.scala 93:102]
  assign cols_12_0_io_top_in_bits = q_252_io_deq_bits; // @[Stab.scala 93:102]
  assign cols_12_0_io_sum_ready = q_524_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_0_io_right_out_ready = q_12_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_0_io_bottom_out_ready = q_436_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_0_clock = clock;
  assign cols_13_0_reset = reset;
  assign cols_13_0_io_left_in_valid = q_12_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_13_0_io_left_in_bits = q_12_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_13_0_io_top_in_valid = q_253_io_deq_valid; // @[Stab.scala 93:102]
  assign cols_13_0_io_top_in_bits = q_253_io_deq_bits; // @[Stab.scala 93:102]
  assign cols_13_0_io_sum_ready = q_525_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_0_io_right_out_ready = q_13_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_0_io_bottom_out_ready = q_451_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_0_clock = clock;
  assign cols_14_0_reset = reset;
  assign cols_14_0_io_left_in_valid = q_13_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_14_0_io_left_in_bits = q_13_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_14_0_io_top_in_valid = q_254_io_deq_valid; // @[Stab.scala 93:102]
  assign cols_14_0_io_top_in_bits = q_254_io_deq_bits; // @[Stab.scala 93:102]
  assign cols_14_0_io_sum_ready = q_526_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_0_io_right_out_ready = q_14_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_0_io_bottom_out_ready = q_466_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_0_clock = clock;
  assign cols_15_0_reset = reset;
  assign cols_15_0_io_left_in_valid = q_14_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_15_0_io_left_in_bits = q_14_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_15_0_io_top_in_valid = q_255_io_deq_valid; // @[Stab.scala 93:102]
  assign cols_15_0_io_top_in_bits = q_255_io_deq_bits; // @[Stab.scala 93:102]
  assign cols_15_0_io_sum_ready = q_527_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_0_io_right_out_ready = 1'h1; // @[Stab.scala 102:51]
  assign cols_15_0_io_bottom_out_ready = q_481_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_1_clock = clock;
  assign cols_0_1_reset = reset;
  assign cols_0_1_io_left_in_valid = q_497_io_deq_valid; // @[Stab.scala 100:101]
  assign cols_0_1_io_left_in_bits = q_497_io_deq_bits; // @[Stab.scala 100:101]
  assign cols_0_1_io_top_in_valid = q_256_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_0_1_io_top_in_bits = q_256_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_0_1_io_sum_ready = q_528_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_1_io_right_out_ready = q_15_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_1_io_bottom_out_ready = q_257_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_1_clock = clock;
  assign cols_1_1_reset = reset;
  assign cols_1_1_io_left_in_valid = q_15_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_1_1_io_left_in_bits = q_15_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_1_1_io_top_in_valid = q_271_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_1_1_io_top_in_bits = q_271_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_1_1_io_sum_ready = q_529_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_1_io_right_out_ready = q_16_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_1_io_bottom_out_ready = q_272_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_1_clock = clock;
  assign cols_2_1_reset = reset;
  assign cols_2_1_io_left_in_valid = q_16_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_2_1_io_left_in_bits = q_16_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_2_1_io_top_in_valid = q_286_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_2_1_io_top_in_bits = q_286_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_2_1_io_sum_ready = q_530_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_1_io_right_out_ready = q_17_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_1_io_bottom_out_ready = q_287_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_1_clock = clock;
  assign cols_3_1_reset = reset;
  assign cols_3_1_io_left_in_valid = q_17_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_3_1_io_left_in_bits = q_17_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_3_1_io_top_in_valid = q_301_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_3_1_io_top_in_bits = q_301_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_3_1_io_sum_ready = q_531_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_1_io_right_out_ready = q_18_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_1_io_bottom_out_ready = q_302_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_1_clock = clock;
  assign cols_4_1_reset = reset;
  assign cols_4_1_io_left_in_valid = q_18_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_4_1_io_left_in_bits = q_18_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_4_1_io_top_in_valid = q_316_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_4_1_io_top_in_bits = q_316_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_4_1_io_sum_ready = q_532_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_1_io_right_out_ready = q_19_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_1_io_bottom_out_ready = q_317_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_1_clock = clock;
  assign cols_5_1_reset = reset;
  assign cols_5_1_io_left_in_valid = q_19_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_5_1_io_left_in_bits = q_19_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_5_1_io_top_in_valid = q_331_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_5_1_io_top_in_bits = q_331_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_5_1_io_sum_ready = q_533_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_1_io_right_out_ready = q_20_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_1_io_bottom_out_ready = q_332_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_1_clock = clock;
  assign cols_6_1_reset = reset;
  assign cols_6_1_io_left_in_valid = q_20_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_6_1_io_left_in_bits = q_20_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_6_1_io_top_in_valid = q_346_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_6_1_io_top_in_bits = q_346_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_6_1_io_sum_ready = q_534_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_1_io_right_out_ready = q_21_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_1_io_bottom_out_ready = q_347_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_1_clock = clock;
  assign cols_7_1_reset = reset;
  assign cols_7_1_io_left_in_valid = q_21_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_7_1_io_left_in_bits = q_21_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_7_1_io_top_in_valid = q_361_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_7_1_io_top_in_bits = q_361_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_7_1_io_sum_ready = q_535_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_1_io_right_out_ready = q_22_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_1_io_bottom_out_ready = q_362_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_1_clock = clock;
  assign cols_8_1_reset = reset;
  assign cols_8_1_io_left_in_valid = q_22_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_8_1_io_left_in_bits = q_22_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_8_1_io_top_in_valid = q_376_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_8_1_io_top_in_bits = q_376_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_8_1_io_sum_ready = q_536_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_1_io_right_out_ready = q_23_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_1_io_bottom_out_ready = q_377_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_1_clock = clock;
  assign cols_9_1_reset = reset;
  assign cols_9_1_io_left_in_valid = q_23_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_9_1_io_left_in_bits = q_23_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_9_1_io_top_in_valid = q_391_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_9_1_io_top_in_bits = q_391_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_9_1_io_sum_ready = q_537_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_1_io_right_out_ready = q_24_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_1_io_bottom_out_ready = q_392_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_1_clock = clock;
  assign cols_10_1_reset = reset;
  assign cols_10_1_io_left_in_valid = q_24_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_10_1_io_left_in_bits = q_24_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_10_1_io_top_in_valid = q_406_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_10_1_io_top_in_bits = q_406_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_10_1_io_sum_ready = q_538_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_1_io_right_out_ready = q_25_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_1_io_bottom_out_ready = q_407_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_1_clock = clock;
  assign cols_11_1_reset = reset;
  assign cols_11_1_io_left_in_valid = q_25_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_11_1_io_left_in_bits = q_25_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_11_1_io_top_in_valid = q_421_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_11_1_io_top_in_bits = q_421_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_11_1_io_sum_ready = q_539_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_1_io_right_out_ready = q_26_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_1_io_bottom_out_ready = q_422_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_1_clock = clock;
  assign cols_12_1_reset = reset;
  assign cols_12_1_io_left_in_valid = q_26_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_12_1_io_left_in_bits = q_26_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_12_1_io_top_in_valid = q_436_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_12_1_io_top_in_bits = q_436_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_12_1_io_sum_ready = q_540_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_1_io_right_out_ready = q_27_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_1_io_bottom_out_ready = q_437_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_1_clock = clock;
  assign cols_13_1_reset = reset;
  assign cols_13_1_io_left_in_valid = q_27_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_13_1_io_left_in_bits = q_27_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_13_1_io_top_in_valid = q_451_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_13_1_io_top_in_bits = q_451_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_13_1_io_sum_ready = q_541_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_1_io_right_out_ready = q_28_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_1_io_bottom_out_ready = q_452_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_1_clock = clock;
  assign cols_14_1_reset = reset;
  assign cols_14_1_io_left_in_valid = q_28_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_14_1_io_left_in_bits = q_28_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_14_1_io_top_in_valid = q_466_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_14_1_io_top_in_bits = q_466_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_14_1_io_sum_ready = q_542_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_1_io_right_out_ready = q_29_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_1_io_bottom_out_ready = q_467_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_1_clock = clock;
  assign cols_15_1_reset = reset;
  assign cols_15_1_io_left_in_valid = q_29_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_15_1_io_left_in_bits = q_29_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_15_1_io_top_in_valid = q_481_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_15_1_io_top_in_bits = q_481_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_15_1_io_sum_ready = q_543_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_1_io_right_out_ready = 1'h1; // @[Stab.scala 102:51]
  assign cols_15_1_io_bottom_out_ready = q_482_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_2_clock = clock;
  assign cols_0_2_reset = reset;
  assign cols_0_2_io_left_in_valid = q_498_io_deq_valid; // @[Stab.scala 100:101]
  assign cols_0_2_io_left_in_bits = q_498_io_deq_bits; // @[Stab.scala 100:101]
  assign cols_0_2_io_top_in_valid = q_257_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_0_2_io_top_in_bits = q_257_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_0_2_io_sum_ready = q_544_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_2_io_right_out_ready = q_30_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_2_io_bottom_out_ready = q_258_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_2_clock = clock;
  assign cols_1_2_reset = reset;
  assign cols_1_2_io_left_in_valid = q_30_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_1_2_io_left_in_bits = q_30_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_1_2_io_top_in_valid = q_272_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_1_2_io_top_in_bits = q_272_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_1_2_io_sum_ready = q_545_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_2_io_right_out_ready = q_31_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_2_io_bottom_out_ready = q_273_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_2_clock = clock;
  assign cols_2_2_reset = reset;
  assign cols_2_2_io_left_in_valid = q_31_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_2_2_io_left_in_bits = q_31_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_2_2_io_top_in_valid = q_287_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_2_2_io_top_in_bits = q_287_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_2_2_io_sum_ready = q_546_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_2_io_right_out_ready = q_32_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_2_io_bottom_out_ready = q_288_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_2_clock = clock;
  assign cols_3_2_reset = reset;
  assign cols_3_2_io_left_in_valid = q_32_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_3_2_io_left_in_bits = q_32_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_3_2_io_top_in_valid = q_302_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_3_2_io_top_in_bits = q_302_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_3_2_io_sum_ready = q_547_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_2_io_right_out_ready = q_33_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_2_io_bottom_out_ready = q_303_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_2_clock = clock;
  assign cols_4_2_reset = reset;
  assign cols_4_2_io_left_in_valid = q_33_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_4_2_io_left_in_bits = q_33_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_4_2_io_top_in_valid = q_317_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_4_2_io_top_in_bits = q_317_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_4_2_io_sum_ready = q_548_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_2_io_right_out_ready = q_34_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_2_io_bottom_out_ready = q_318_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_2_clock = clock;
  assign cols_5_2_reset = reset;
  assign cols_5_2_io_left_in_valid = q_34_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_5_2_io_left_in_bits = q_34_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_5_2_io_top_in_valid = q_332_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_5_2_io_top_in_bits = q_332_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_5_2_io_sum_ready = q_549_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_2_io_right_out_ready = q_35_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_2_io_bottom_out_ready = q_333_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_2_clock = clock;
  assign cols_6_2_reset = reset;
  assign cols_6_2_io_left_in_valid = q_35_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_6_2_io_left_in_bits = q_35_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_6_2_io_top_in_valid = q_347_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_6_2_io_top_in_bits = q_347_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_6_2_io_sum_ready = q_550_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_2_io_right_out_ready = q_36_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_2_io_bottom_out_ready = q_348_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_2_clock = clock;
  assign cols_7_2_reset = reset;
  assign cols_7_2_io_left_in_valid = q_36_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_7_2_io_left_in_bits = q_36_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_7_2_io_top_in_valid = q_362_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_7_2_io_top_in_bits = q_362_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_7_2_io_sum_ready = q_551_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_2_io_right_out_ready = q_37_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_2_io_bottom_out_ready = q_363_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_2_clock = clock;
  assign cols_8_2_reset = reset;
  assign cols_8_2_io_left_in_valid = q_37_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_8_2_io_left_in_bits = q_37_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_8_2_io_top_in_valid = q_377_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_8_2_io_top_in_bits = q_377_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_8_2_io_sum_ready = q_552_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_2_io_right_out_ready = q_38_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_2_io_bottom_out_ready = q_378_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_2_clock = clock;
  assign cols_9_2_reset = reset;
  assign cols_9_2_io_left_in_valid = q_38_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_9_2_io_left_in_bits = q_38_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_9_2_io_top_in_valid = q_392_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_9_2_io_top_in_bits = q_392_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_9_2_io_sum_ready = q_553_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_2_io_right_out_ready = q_39_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_2_io_bottom_out_ready = q_393_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_2_clock = clock;
  assign cols_10_2_reset = reset;
  assign cols_10_2_io_left_in_valid = q_39_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_10_2_io_left_in_bits = q_39_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_10_2_io_top_in_valid = q_407_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_10_2_io_top_in_bits = q_407_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_10_2_io_sum_ready = q_554_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_2_io_right_out_ready = q_40_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_2_io_bottom_out_ready = q_408_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_2_clock = clock;
  assign cols_11_2_reset = reset;
  assign cols_11_2_io_left_in_valid = q_40_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_11_2_io_left_in_bits = q_40_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_11_2_io_top_in_valid = q_422_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_11_2_io_top_in_bits = q_422_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_11_2_io_sum_ready = q_555_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_2_io_right_out_ready = q_41_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_2_io_bottom_out_ready = q_423_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_2_clock = clock;
  assign cols_12_2_reset = reset;
  assign cols_12_2_io_left_in_valid = q_41_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_12_2_io_left_in_bits = q_41_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_12_2_io_top_in_valid = q_437_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_12_2_io_top_in_bits = q_437_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_12_2_io_sum_ready = q_556_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_2_io_right_out_ready = q_42_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_2_io_bottom_out_ready = q_438_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_2_clock = clock;
  assign cols_13_2_reset = reset;
  assign cols_13_2_io_left_in_valid = q_42_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_13_2_io_left_in_bits = q_42_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_13_2_io_top_in_valid = q_452_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_13_2_io_top_in_bits = q_452_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_13_2_io_sum_ready = q_557_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_2_io_right_out_ready = q_43_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_2_io_bottom_out_ready = q_453_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_2_clock = clock;
  assign cols_14_2_reset = reset;
  assign cols_14_2_io_left_in_valid = q_43_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_14_2_io_left_in_bits = q_43_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_14_2_io_top_in_valid = q_467_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_14_2_io_top_in_bits = q_467_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_14_2_io_sum_ready = q_558_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_2_io_right_out_ready = q_44_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_2_io_bottom_out_ready = q_468_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_2_clock = clock;
  assign cols_15_2_reset = reset;
  assign cols_15_2_io_left_in_valid = q_44_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_15_2_io_left_in_bits = q_44_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_15_2_io_top_in_valid = q_482_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_15_2_io_top_in_bits = q_482_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_15_2_io_sum_ready = q_559_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_2_io_right_out_ready = 1'h1; // @[Stab.scala 102:51]
  assign cols_15_2_io_bottom_out_ready = q_483_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_3_clock = clock;
  assign cols_0_3_reset = reset;
  assign cols_0_3_io_left_in_valid = q_499_io_deq_valid; // @[Stab.scala 100:101]
  assign cols_0_3_io_left_in_bits = q_499_io_deq_bits; // @[Stab.scala 100:101]
  assign cols_0_3_io_top_in_valid = q_258_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_0_3_io_top_in_bits = q_258_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_0_3_io_sum_ready = q_560_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_3_io_right_out_ready = q_45_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_3_io_bottom_out_ready = q_259_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_3_clock = clock;
  assign cols_1_3_reset = reset;
  assign cols_1_3_io_left_in_valid = q_45_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_1_3_io_left_in_bits = q_45_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_1_3_io_top_in_valid = q_273_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_1_3_io_top_in_bits = q_273_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_1_3_io_sum_ready = q_561_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_3_io_right_out_ready = q_46_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_3_io_bottom_out_ready = q_274_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_3_clock = clock;
  assign cols_2_3_reset = reset;
  assign cols_2_3_io_left_in_valid = q_46_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_2_3_io_left_in_bits = q_46_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_2_3_io_top_in_valid = q_288_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_2_3_io_top_in_bits = q_288_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_2_3_io_sum_ready = q_562_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_3_io_right_out_ready = q_47_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_3_io_bottom_out_ready = q_289_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_3_clock = clock;
  assign cols_3_3_reset = reset;
  assign cols_3_3_io_left_in_valid = q_47_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_3_3_io_left_in_bits = q_47_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_3_3_io_top_in_valid = q_303_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_3_3_io_top_in_bits = q_303_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_3_3_io_sum_ready = q_563_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_3_io_right_out_ready = q_48_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_3_io_bottom_out_ready = q_304_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_3_clock = clock;
  assign cols_4_3_reset = reset;
  assign cols_4_3_io_left_in_valid = q_48_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_4_3_io_left_in_bits = q_48_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_4_3_io_top_in_valid = q_318_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_4_3_io_top_in_bits = q_318_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_4_3_io_sum_ready = q_564_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_3_io_right_out_ready = q_49_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_3_io_bottom_out_ready = q_319_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_3_clock = clock;
  assign cols_5_3_reset = reset;
  assign cols_5_3_io_left_in_valid = q_49_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_5_3_io_left_in_bits = q_49_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_5_3_io_top_in_valid = q_333_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_5_3_io_top_in_bits = q_333_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_5_3_io_sum_ready = q_565_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_3_io_right_out_ready = q_50_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_3_io_bottom_out_ready = q_334_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_3_clock = clock;
  assign cols_6_3_reset = reset;
  assign cols_6_3_io_left_in_valid = q_50_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_6_3_io_left_in_bits = q_50_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_6_3_io_top_in_valid = q_348_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_6_3_io_top_in_bits = q_348_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_6_3_io_sum_ready = q_566_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_3_io_right_out_ready = q_51_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_3_io_bottom_out_ready = q_349_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_3_clock = clock;
  assign cols_7_3_reset = reset;
  assign cols_7_3_io_left_in_valid = q_51_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_7_3_io_left_in_bits = q_51_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_7_3_io_top_in_valid = q_363_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_7_3_io_top_in_bits = q_363_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_7_3_io_sum_ready = q_567_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_3_io_right_out_ready = q_52_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_3_io_bottom_out_ready = q_364_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_3_clock = clock;
  assign cols_8_3_reset = reset;
  assign cols_8_3_io_left_in_valid = q_52_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_8_3_io_left_in_bits = q_52_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_8_3_io_top_in_valid = q_378_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_8_3_io_top_in_bits = q_378_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_8_3_io_sum_ready = q_568_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_3_io_right_out_ready = q_53_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_3_io_bottom_out_ready = q_379_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_3_clock = clock;
  assign cols_9_3_reset = reset;
  assign cols_9_3_io_left_in_valid = q_53_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_9_3_io_left_in_bits = q_53_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_9_3_io_top_in_valid = q_393_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_9_3_io_top_in_bits = q_393_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_9_3_io_sum_ready = q_569_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_3_io_right_out_ready = q_54_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_3_io_bottom_out_ready = q_394_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_3_clock = clock;
  assign cols_10_3_reset = reset;
  assign cols_10_3_io_left_in_valid = q_54_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_10_3_io_left_in_bits = q_54_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_10_3_io_top_in_valid = q_408_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_10_3_io_top_in_bits = q_408_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_10_3_io_sum_ready = q_570_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_3_io_right_out_ready = q_55_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_3_io_bottom_out_ready = q_409_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_3_clock = clock;
  assign cols_11_3_reset = reset;
  assign cols_11_3_io_left_in_valid = q_55_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_11_3_io_left_in_bits = q_55_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_11_3_io_top_in_valid = q_423_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_11_3_io_top_in_bits = q_423_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_11_3_io_sum_ready = q_571_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_3_io_right_out_ready = q_56_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_3_io_bottom_out_ready = q_424_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_3_clock = clock;
  assign cols_12_3_reset = reset;
  assign cols_12_3_io_left_in_valid = q_56_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_12_3_io_left_in_bits = q_56_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_12_3_io_top_in_valid = q_438_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_12_3_io_top_in_bits = q_438_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_12_3_io_sum_ready = q_572_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_3_io_right_out_ready = q_57_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_3_io_bottom_out_ready = q_439_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_3_clock = clock;
  assign cols_13_3_reset = reset;
  assign cols_13_3_io_left_in_valid = q_57_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_13_3_io_left_in_bits = q_57_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_13_3_io_top_in_valid = q_453_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_13_3_io_top_in_bits = q_453_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_13_3_io_sum_ready = q_573_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_3_io_right_out_ready = q_58_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_3_io_bottom_out_ready = q_454_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_3_clock = clock;
  assign cols_14_3_reset = reset;
  assign cols_14_3_io_left_in_valid = q_58_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_14_3_io_left_in_bits = q_58_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_14_3_io_top_in_valid = q_468_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_14_3_io_top_in_bits = q_468_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_14_3_io_sum_ready = q_574_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_3_io_right_out_ready = q_59_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_3_io_bottom_out_ready = q_469_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_3_clock = clock;
  assign cols_15_3_reset = reset;
  assign cols_15_3_io_left_in_valid = q_59_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_15_3_io_left_in_bits = q_59_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_15_3_io_top_in_valid = q_483_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_15_3_io_top_in_bits = q_483_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_15_3_io_sum_ready = q_575_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_3_io_right_out_ready = 1'h1; // @[Stab.scala 102:51]
  assign cols_15_3_io_bottom_out_ready = q_484_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_4_clock = clock;
  assign cols_0_4_reset = reset;
  assign cols_0_4_io_left_in_valid = q_500_io_deq_valid; // @[Stab.scala 100:101]
  assign cols_0_4_io_left_in_bits = q_500_io_deq_bits; // @[Stab.scala 100:101]
  assign cols_0_4_io_top_in_valid = q_259_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_0_4_io_top_in_bits = q_259_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_0_4_io_sum_ready = q_576_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_4_io_right_out_ready = q_60_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_4_io_bottom_out_ready = q_260_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_4_clock = clock;
  assign cols_1_4_reset = reset;
  assign cols_1_4_io_left_in_valid = q_60_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_1_4_io_left_in_bits = q_60_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_1_4_io_top_in_valid = q_274_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_1_4_io_top_in_bits = q_274_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_1_4_io_sum_ready = q_577_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_4_io_right_out_ready = q_61_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_4_io_bottom_out_ready = q_275_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_4_clock = clock;
  assign cols_2_4_reset = reset;
  assign cols_2_4_io_left_in_valid = q_61_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_2_4_io_left_in_bits = q_61_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_2_4_io_top_in_valid = q_289_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_2_4_io_top_in_bits = q_289_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_2_4_io_sum_ready = q_578_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_4_io_right_out_ready = q_62_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_4_io_bottom_out_ready = q_290_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_4_clock = clock;
  assign cols_3_4_reset = reset;
  assign cols_3_4_io_left_in_valid = q_62_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_3_4_io_left_in_bits = q_62_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_3_4_io_top_in_valid = q_304_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_3_4_io_top_in_bits = q_304_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_3_4_io_sum_ready = q_579_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_4_io_right_out_ready = q_63_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_4_io_bottom_out_ready = q_305_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_4_clock = clock;
  assign cols_4_4_reset = reset;
  assign cols_4_4_io_left_in_valid = q_63_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_4_4_io_left_in_bits = q_63_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_4_4_io_top_in_valid = q_319_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_4_4_io_top_in_bits = q_319_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_4_4_io_sum_ready = q_580_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_4_io_right_out_ready = q_64_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_4_io_bottom_out_ready = q_320_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_4_clock = clock;
  assign cols_5_4_reset = reset;
  assign cols_5_4_io_left_in_valid = q_64_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_5_4_io_left_in_bits = q_64_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_5_4_io_top_in_valid = q_334_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_5_4_io_top_in_bits = q_334_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_5_4_io_sum_ready = q_581_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_4_io_right_out_ready = q_65_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_4_io_bottom_out_ready = q_335_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_4_clock = clock;
  assign cols_6_4_reset = reset;
  assign cols_6_4_io_left_in_valid = q_65_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_6_4_io_left_in_bits = q_65_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_6_4_io_top_in_valid = q_349_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_6_4_io_top_in_bits = q_349_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_6_4_io_sum_ready = q_582_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_4_io_right_out_ready = q_66_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_4_io_bottom_out_ready = q_350_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_4_clock = clock;
  assign cols_7_4_reset = reset;
  assign cols_7_4_io_left_in_valid = q_66_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_7_4_io_left_in_bits = q_66_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_7_4_io_top_in_valid = q_364_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_7_4_io_top_in_bits = q_364_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_7_4_io_sum_ready = q_583_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_4_io_right_out_ready = q_67_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_4_io_bottom_out_ready = q_365_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_4_clock = clock;
  assign cols_8_4_reset = reset;
  assign cols_8_4_io_left_in_valid = q_67_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_8_4_io_left_in_bits = q_67_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_8_4_io_top_in_valid = q_379_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_8_4_io_top_in_bits = q_379_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_8_4_io_sum_ready = q_584_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_4_io_right_out_ready = q_68_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_4_io_bottom_out_ready = q_380_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_4_clock = clock;
  assign cols_9_4_reset = reset;
  assign cols_9_4_io_left_in_valid = q_68_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_9_4_io_left_in_bits = q_68_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_9_4_io_top_in_valid = q_394_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_9_4_io_top_in_bits = q_394_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_9_4_io_sum_ready = q_585_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_4_io_right_out_ready = q_69_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_4_io_bottom_out_ready = q_395_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_4_clock = clock;
  assign cols_10_4_reset = reset;
  assign cols_10_4_io_left_in_valid = q_69_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_10_4_io_left_in_bits = q_69_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_10_4_io_top_in_valid = q_409_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_10_4_io_top_in_bits = q_409_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_10_4_io_sum_ready = q_586_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_4_io_right_out_ready = q_70_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_4_io_bottom_out_ready = q_410_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_4_clock = clock;
  assign cols_11_4_reset = reset;
  assign cols_11_4_io_left_in_valid = q_70_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_11_4_io_left_in_bits = q_70_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_11_4_io_top_in_valid = q_424_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_11_4_io_top_in_bits = q_424_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_11_4_io_sum_ready = q_587_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_4_io_right_out_ready = q_71_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_4_io_bottom_out_ready = q_425_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_4_clock = clock;
  assign cols_12_4_reset = reset;
  assign cols_12_4_io_left_in_valid = q_71_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_12_4_io_left_in_bits = q_71_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_12_4_io_top_in_valid = q_439_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_12_4_io_top_in_bits = q_439_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_12_4_io_sum_ready = q_588_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_4_io_right_out_ready = q_72_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_4_io_bottom_out_ready = q_440_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_4_clock = clock;
  assign cols_13_4_reset = reset;
  assign cols_13_4_io_left_in_valid = q_72_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_13_4_io_left_in_bits = q_72_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_13_4_io_top_in_valid = q_454_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_13_4_io_top_in_bits = q_454_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_13_4_io_sum_ready = q_589_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_4_io_right_out_ready = q_73_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_4_io_bottom_out_ready = q_455_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_4_clock = clock;
  assign cols_14_4_reset = reset;
  assign cols_14_4_io_left_in_valid = q_73_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_14_4_io_left_in_bits = q_73_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_14_4_io_top_in_valid = q_469_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_14_4_io_top_in_bits = q_469_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_14_4_io_sum_ready = q_590_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_4_io_right_out_ready = q_74_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_4_io_bottom_out_ready = q_470_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_4_clock = clock;
  assign cols_15_4_reset = reset;
  assign cols_15_4_io_left_in_valid = q_74_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_15_4_io_left_in_bits = q_74_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_15_4_io_top_in_valid = q_484_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_15_4_io_top_in_bits = q_484_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_15_4_io_sum_ready = q_591_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_4_io_right_out_ready = 1'h1; // @[Stab.scala 102:51]
  assign cols_15_4_io_bottom_out_ready = q_485_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_5_clock = clock;
  assign cols_0_5_reset = reset;
  assign cols_0_5_io_left_in_valid = q_501_io_deq_valid; // @[Stab.scala 100:101]
  assign cols_0_5_io_left_in_bits = q_501_io_deq_bits; // @[Stab.scala 100:101]
  assign cols_0_5_io_top_in_valid = q_260_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_0_5_io_top_in_bits = q_260_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_0_5_io_sum_ready = q_592_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_5_io_right_out_ready = q_75_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_5_io_bottom_out_ready = q_261_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_5_clock = clock;
  assign cols_1_5_reset = reset;
  assign cols_1_5_io_left_in_valid = q_75_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_1_5_io_left_in_bits = q_75_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_1_5_io_top_in_valid = q_275_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_1_5_io_top_in_bits = q_275_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_1_5_io_sum_ready = q_593_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_5_io_right_out_ready = q_76_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_5_io_bottom_out_ready = q_276_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_5_clock = clock;
  assign cols_2_5_reset = reset;
  assign cols_2_5_io_left_in_valid = q_76_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_2_5_io_left_in_bits = q_76_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_2_5_io_top_in_valid = q_290_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_2_5_io_top_in_bits = q_290_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_2_5_io_sum_ready = q_594_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_5_io_right_out_ready = q_77_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_5_io_bottom_out_ready = q_291_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_5_clock = clock;
  assign cols_3_5_reset = reset;
  assign cols_3_5_io_left_in_valid = q_77_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_3_5_io_left_in_bits = q_77_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_3_5_io_top_in_valid = q_305_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_3_5_io_top_in_bits = q_305_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_3_5_io_sum_ready = q_595_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_5_io_right_out_ready = q_78_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_5_io_bottom_out_ready = q_306_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_5_clock = clock;
  assign cols_4_5_reset = reset;
  assign cols_4_5_io_left_in_valid = q_78_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_4_5_io_left_in_bits = q_78_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_4_5_io_top_in_valid = q_320_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_4_5_io_top_in_bits = q_320_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_4_5_io_sum_ready = q_596_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_5_io_right_out_ready = q_79_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_5_io_bottom_out_ready = q_321_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_5_clock = clock;
  assign cols_5_5_reset = reset;
  assign cols_5_5_io_left_in_valid = q_79_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_5_5_io_left_in_bits = q_79_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_5_5_io_top_in_valid = q_335_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_5_5_io_top_in_bits = q_335_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_5_5_io_sum_ready = q_597_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_5_io_right_out_ready = q_80_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_5_io_bottom_out_ready = q_336_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_5_clock = clock;
  assign cols_6_5_reset = reset;
  assign cols_6_5_io_left_in_valid = q_80_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_6_5_io_left_in_bits = q_80_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_6_5_io_top_in_valid = q_350_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_6_5_io_top_in_bits = q_350_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_6_5_io_sum_ready = q_598_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_5_io_right_out_ready = q_81_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_5_io_bottom_out_ready = q_351_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_5_clock = clock;
  assign cols_7_5_reset = reset;
  assign cols_7_5_io_left_in_valid = q_81_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_7_5_io_left_in_bits = q_81_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_7_5_io_top_in_valid = q_365_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_7_5_io_top_in_bits = q_365_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_7_5_io_sum_ready = q_599_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_5_io_right_out_ready = q_82_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_5_io_bottom_out_ready = q_366_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_5_clock = clock;
  assign cols_8_5_reset = reset;
  assign cols_8_5_io_left_in_valid = q_82_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_8_5_io_left_in_bits = q_82_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_8_5_io_top_in_valid = q_380_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_8_5_io_top_in_bits = q_380_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_8_5_io_sum_ready = q_600_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_5_io_right_out_ready = q_83_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_5_io_bottom_out_ready = q_381_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_5_clock = clock;
  assign cols_9_5_reset = reset;
  assign cols_9_5_io_left_in_valid = q_83_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_9_5_io_left_in_bits = q_83_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_9_5_io_top_in_valid = q_395_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_9_5_io_top_in_bits = q_395_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_9_5_io_sum_ready = q_601_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_5_io_right_out_ready = q_84_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_5_io_bottom_out_ready = q_396_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_5_clock = clock;
  assign cols_10_5_reset = reset;
  assign cols_10_5_io_left_in_valid = q_84_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_10_5_io_left_in_bits = q_84_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_10_5_io_top_in_valid = q_410_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_10_5_io_top_in_bits = q_410_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_10_5_io_sum_ready = q_602_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_5_io_right_out_ready = q_85_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_5_io_bottom_out_ready = q_411_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_5_clock = clock;
  assign cols_11_5_reset = reset;
  assign cols_11_5_io_left_in_valid = q_85_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_11_5_io_left_in_bits = q_85_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_11_5_io_top_in_valid = q_425_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_11_5_io_top_in_bits = q_425_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_11_5_io_sum_ready = q_603_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_5_io_right_out_ready = q_86_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_5_io_bottom_out_ready = q_426_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_5_clock = clock;
  assign cols_12_5_reset = reset;
  assign cols_12_5_io_left_in_valid = q_86_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_12_5_io_left_in_bits = q_86_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_12_5_io_top_in_valid = q_440_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_12_5_io_top_in_bits = q_440_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_12_5_io_sum_ready = q_604_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_5_io_right_out_ready = q_87_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_5_io_bottom_out_ready = q_441_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_5_clock = clock;
  assign cols_13_5_reset = reset;
  assign cols_13_5_io_left_in_valid = q_87_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_13_5_io_left_in_bits = q_87_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_13_5_io_top_in_valid = q_455_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_13_5_io_top_in_bits = q_455_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_13_5_io_sum_ready = q_605_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_5_io_right_out_ready = q_88_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_5_io_bottom_out_ready = q_456_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_5_clock = clock;
  assign cols_14_5_reset = reset;
  assign cols_14_5_io_left_in_valid = q_88_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_14_5_io_left_in_bits = q_88_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_14_5_io_top_in_valid = q_470_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_14_5_io_top_in_bits = q_470_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_14_5_io_sum_ready = q_606_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_5_io_right_out_ready = q_89_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_5_io_bottom_out_ready = q_471_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_5_clock = clock;
  assign cols_15_5_reset = reset;
  assign cols_15_5_io_left_in_valid = q_89_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_15_5_io_left_in_bits = q_89_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_15_5_io_top_in_valid = q_485_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_15_5_io_top_in_bits = q_485_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_15_5_io_sum_ready = q_607_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_5_io_right_out_ready = 1'h1; // @[Stab.scala 102:51]
  assign cols_15_5_io_bottom_out_ready = q_486_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_6_clock = clock;
  assign cols_0_6_reset = reset;
  assign cols_0_6_io_left_in_valid = q_502_io_deq_valid; // @[Stab.scala 100:101]
  assign cols_0_6_io_left_in_bits = q_502_io_deq_bits; // @[Stab.scala 100:101]
  assign cols_0_6_io_top_in_valid = q_261_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_0_6_io_top_in_bits = q_261_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_0_6_io_sum_ready = q_608_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_6_io_right_out_ready = q_90_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_6_io_bottom_out_ready = q_262_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_6_clock = clock;
  assign cols_1_6_reset = reset;
  assign cols_1_6_io_left_in_valid = q_90_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_1_6_io_left_in_bits = q_90_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_1_6_io_top_in_valid = q_276_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_1_6_io_top_in_bits = q_276_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_1_6_io_sum_ready = q_609_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_6_io_right_out_ready = q_91_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_6_io_bottom_out_ready = q_277_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_6_clock = clock;
  assign cols_2_6_reset = reset;
  assign cols_2_6_io_left_in_valid = q_91_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_2_6_io_left_in_bits = q_91_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_2_6_io_top_in_valid = q_291_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_2_6_io_top_in_bits = q_291_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_2_6_io_sum_ready = q_610_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_6_io_right_out_ready = q_92_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_6_io_bottom_out_ready = q_292_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_6_clock = clock;
  assign cols_3_6_reset = reset;
  assign cols_3_6_io_left_in_valid = q_92_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_3_6_io_left_in_bits = q_92_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_3_6_io_top_in_valid = q_306_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_3_6_io_top_in_bits = q_306_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_3_6_io_sum_ready = q_611_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_6_io_right_out_ready = q_93_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_6_io_bottom_out_ready = q_307_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_6_clock = clock;
  assign cols_4_6_reset = reset;
  assign cols_4_6_io_left_in_valid = q_93_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_4_6_io_left_in_bits = q_93_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_4_6_io_top_in_valid = q_321_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_4_6_io_top_in_bits = q_321_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_4_6_io_sum_ready = q_612_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_6_io_right_out_ready = q_94_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_6_io_bottom_out_ready = q_322_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_6_clock = clock;
  assign cols_5_6_reset = reset;
  assign cols_5_6_io_left_in_valid = q_94_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_5_6_io_left_in_bits = q_94_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_5_6_io_top_in_valid = q_336_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_5_6_io_top_in_bits = q_336_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_5_6_io_sum_ready = q_613_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_6_io_right_out_ready = q_95_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_6_io_bottom_out_ready = q_337_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_6_clock = clock;
  assign cols_6_6_reset = reset;
  assign cols_6_6_io_left_in_valid = q_95_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_6_6_io_left_in_bits = q_95_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_6_6_io_top_in_valid = q_351_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_6_6_io_top_in_bits = q_351_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_6_6_io_sum_ready = q_614_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_6_io_right_out_ready = q_96_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_6_io_bottom_out_ready = q_352_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_6_clock = clock;
  assign cols_7_6_reset = reset;
  assign cols_7_6_io_left_in_valid = q_96_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_7_6_io_left_in_bits = q_96_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_7_6_io_top_in_valid = q_366_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_7_6_io_top_in_bits = q_366_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_7_6_io_sum_ready = q_615_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_6_io_right_out_ready = q_97_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_6_io_bottom_out_ready = q_367_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_6_clock = clock;
  assign cols_8_6_reset = reset;
  assign cols_8_6_io_left_in_valid = q_97_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_8_6_io_left_in_bits = q_97_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_8_6_io_top_in_valid = q_381_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_8_6_io_top_in_bits = q_381_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_8_6_io_sum_ready = q_616_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_6_io_right_out_ready = q_98_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_6_io_bottom_out_ready = q_382_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_6_clock = clock;
  assign cols_9_6_reset = reset;
  assign cols_9_6_io_left_in_valid = q_98_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_9_6_io_left_in_bits = q_98_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_9_6_io_top_in_valid = q_396_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_9_6_io_top_in_bits = q_396_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_9_6_io_sum_ready = q_617_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_6_io_right_out_ready = q_99_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_6_io_bottom_out_ready = q_397_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_6_clock = clock;
  assign cols_10_6_reset = reset;
  assign cols_10_6_io_left_in_valid = q_99_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_10_6_io_left_in_bits = q_99_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_10_6_io_top_in_valid = q_411_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_10_6_io_top_in_bits = q_411_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_10_6_io_sum_ready = q_618_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_6_io_right_out_ready = q_100_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_6_io_bottom_out_ready = q_412_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_6_clock = clock;
  assign cols_11_6_reset = reset;
  assign cols_11_6_io_left_in_valid = q_100_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_11_6_io_left_in_bits = q_100_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_11_6_io_top_in_valid = q_426_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_11_6_io_top_in_bits = q_426_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_11_6_io_sum_ready = q_619_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_6_io_right_out_ready = q_101_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_6_io_bottom_out_ready = q_427_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_6_clock = clock;
  assign cols_12_6_reset = reset;
  assign cols_12_6_io_left_in_valid = q_101_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_12_6_io_left_in_bits = q_101_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_12_6_io_top_in_valid = q_441_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_12_6_io_top_in_bits = q_441_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_12_6_io_sum_ready = q_620_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_6_io_right_out_ready = q_102_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_6_io_bottom_out_ready = q_442_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_6_clock = clock;
  assign cols_13_6_reset = reset;
  assign cols_13_6_io_left_in_valid = q_102_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_13_6_io_left_in_bits = q_102_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_13_6_io_top_in_valid = q_456_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_13_6_io_top_in_bits = q_456_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_13_6_io_sum_ready = q_621_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_6_io_right_out_ready = q_103_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_6_io_bottom_out_ready = q_457_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_6_clock = clock;
  assign cols_14_6_reset = reset;
  assign cols_14_6_io_left_in_valid = q_103_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_14_6_io_left_in_bits = q_103_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_14_6_io_top_in_valid = q_471_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_14_6_io_top_in_bits = q_471_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_14_6_io_sum_ready = q_622_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_6_io_right_out_ready = q_104_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_6_io_bottom_out_ready = q_472_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_6_clock = clock;
  assign cols_15_6_reset = reset;
  assign cols_15_6_io_left_in_valid = q_104_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_15_6_io_left_in_bits = q_104_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_15_6_io_top_in_valid = q_486_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_15_6_io_top_in_bits = q_486_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_15_6_io_sum_ready = q_623_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_6_io_right_out_ready = 1'h1; // @[Stab.scala 102:51]
  assign cols_15_6_io_bottom_out_ready = q_487_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_7_clock = clock;
  assign cols_0_7_reset = reset;
  assign cols_0_7_io_left_in_valid = q_503_io_deq_valid; // @[Stab.scala 100:101]
  assign cols_0_7_io_left_in_bits = q_503_io_deq_bits; // @[Stab.scala 100:101]
  assign cols_0_7_io_top_in_valid = q_262_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_0_7_io_top_in_bits = q_262_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_0_7_io_sum_ready = q_624_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_7_io_right_out_ready = q_105_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_7_io_bottom_out_ready = q_263_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_7_clock = clock;
  assign cols_1_7_reset = reset;
  assign cols_1_7_io_left_in_valid = q_105_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_1_7_io_left_in_bits = q_105_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_1_7_io_top_in_valid = q_277_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_1_7_io_top_in_bits = q_277_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_1_7_io_sum_ready = q_625_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_7_io_right_out_ready = q_106_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_7_io_bottom_out_ready = q_278_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_7_clock = clock;
  assign cols_2_7_reset = reset;
  assign cols_2_7_io_left_in_valid = q_106_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_2_7_io_left_in_bits = q_106_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_2_7_io_top_in_valid = q_292_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_2_7_io_top_in_bits = q_292_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_2_7_io_sum_ready = q_626_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_7_io_right_out_ready = q_107_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_7_io_bottom_out_ready = q_293_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_7_clock = clock;
  assign cols_3_7_reset = reset;
  assign cols_3_7_io_left_in_valid = q_107_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_3_7_io_left_in_bits = q_107_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_3_7_io_top_in_valid = q_307_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_3_7_io_top_in_bits = q_307_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_3_7_io_sum_ready = q_627_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_7_io_right_out_ready = q_108_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_7_io_bottom_out_ready = q_308_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_7_clock = clock;
  assign cols_4_7_reset = reset;
  assign cols_4_7_io_left_in_valid = q_108_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_4_7_io_left_in_bits = q_108_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_4_7_io_top_in_valid = q_322_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_4_7_io_top_in_bits = q_322_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_4_7_io_sum_ready = q_628_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_7_io_right_out_ready = q_109_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_7_io_bottom_out_ready = q_323_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_7_clock = clock;
  assign cols_5_7_reset = reset;
  assign cols_5_7_io_left_in_valid = q_109_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_5_7_io_left_in_bits = q_109_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_5_7_io_top_in_valid = q_337_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_5_7_io_top_in_bits = q_337_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_5_7_io_sum_ready = q_629_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_7_io_right_out_ready = q_110_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_7_io_bottom_out_ready = q_338_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_7_clock = clock;
  assign cols_6_7_reset = reset;
  assign cols_6_7_io_left_in_valid = q_110_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_6_7_io_left_in_bits = q_110_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_6_7_io_top_in_valid = q_352_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_6_7_io_top_in_bits = q_352_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_6_7_io_sum_ready = q_630_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_7_io_right_out_ready = q_111_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_7_io_bottom_out_ready = q_353_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_7_clock = clock;
  assign cols_7_7_reset = reset;
  assign cols_7_7_io_left_in_valid = q_111_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_7_7_io_left_in_bits = q_111_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_7_7_io_top_in_valid = q_367_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_7_7_io_top_in_bits = q_367_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_7_7_io_sum_ready = q_631_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_7_io_right_out_ready = q_112_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_7_io_bottom_out_ready = q_368_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_7_clock = clock;
  assign cols_8_7_reset = reset;
  assign cols_8_7_io_left_in_valid = q_112_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_8_7_io_left_in_bits = q_112_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_8_7_io_top_in_valid = q_382_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_8_7_io_top_in_bits = q_382_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_8_7_io_sum_ready = q_632_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_7_io_right_out_ready = q_113_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_7_io_bottom_out_ready = q_383_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_7_clock = clock;
  assign cols_9_7_reset = reset;
  assign cols_9_7_io_left_in_valid = q_113_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_9_7_io_left_in_bits = q_113_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_9_7_io_top_in_valid = q_397_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_9_7_io_top_in_bits = q_397_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_9_7_io_sum_ready = q_633_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_7_io_right_out_ready = q_114_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_7_io_bottom_out_ready = q_398_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_7_clock = clock;
  assign cols_10_7_reset = reset;
  assign cols_10_7_io_left_in_valid = q_114_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_10_7_io_left_in_bits = q_114_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_10_7_io_top_in_valid = q_412_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_10_7_io_top_in_bits = q_412_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_10_7_io_sum_ready = q_634_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_7_io_right_out_ready = q_115_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_7_io_bottom_out_ready = q_413_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_7_clock = clock;
  assign cols_11_7_reset = reset;
  assign cols_11_7_io_left_in_valid = q_115_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_11_7_io_left_in_bits = q_115_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_11_7_io_top_in_valid = q_427_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_11_7_io_top_in_bits = q_427_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_11_7_io_sum_ready = q_635_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_7_io_right_out_ready = q_116_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_7_io_bottom_out_ready = q_428_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_7_clock = clock;
  assign cols_12_7_reset = reset;
  assign cols_12_7_io_left_in_valid = q_116_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_12_7_io_left_in_bits = q_116_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_12_7_io_top_in_valid = q_442_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_12_7_io_top_in_bits = q_442_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_12_7_io_sum_ready = q_636_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_7_io_right_out_ready = q_117_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_7_io_bottom_out_ready = q_443_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_7_clock = clock;
  assign cols_13_7_reset = reset;
  assign cols_13_7_io_left_in_valid = q_117_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_13_7_io_left_in_bits = q_117_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_13_7_io_top_in_valid = q_457_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_13_7_io_top_in_bits = q_457_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_13_7_io_sum_ready = q_637_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_7_io_right_out_ready = q_118_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_7_io_bottom_out_ready = q_458_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_7_clock = clock;
  assign cols_14_7_reset = reset;
  assign cols_14_7_io_left_in_valid = q_118_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_14_7_io_left_in_bits = q_118_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_14_7_io_top_in_valid = q_472_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_14_7_io_top_in_bits = q_472_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_14_7_io_sum_ready = q_638_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_7_io_right_out_ready = q_119_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_7_io_bottom_out_ready = q_473_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_7_clock = clock;
  assign cols_15_7_reset = reset;
  assign cols_15_7_io_left_in_valid = q_119_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_15_7_io_left_in_bits = q_119_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_15_7_io_top_in_valid = q_487_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_15_7_io_top_in_bits = q_487_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_15_7_io_sum_ready = q_639_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_7_io_right_out_ready = 1'h1; // @[Stab.scala 102:51]
  assign cols_15_7_io_bottom_out_ready = q_488_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_8_clock = clock;
  assign cols_0_8_reset = reset;
  assign cols_0_8_io_left_in_valid = q_504_io_deq_valid; // @[Stab.scala 100:101]
  assign cols_0_8_io_left_in_bits = q_504_io_deq_bits; // @[Stab.scala 100:101]
  assign cols_0_8_io_top_in_valid = q_263_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_0_8_io_top_in_bits = q_263_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_0_8_io_sum_ready = q_640_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_8_io_right_out_ready = q_120_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_8_io_bottom_out_ready = q_264_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_8_clock = clock;
  assign cols_1_8_reset = reset;
  assign cols_1_8_io_left_in_valid = q_120_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_1_8_io_left_in_bits = q_120_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_1_8_io_top_in_valid = q_278_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_1_8_io_top_in_bits = q_278_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_1_8_io_sum_ready = q_641_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_8_io_right_out_ready = q_121_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_8_io_bottom_out_ready = q_279_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_8_clock = clock;
  assign cols_2_8_reset = reset;
  assign cols_2_8_io_left_in_valid = q_121_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_2_8_io_left_in_bits = q_121_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_2_8_io_top_in_valid = q_293_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_2_8_io_top_in_bits = q_293_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_2_8_io_sum_ready = q_642_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_8_io_right_out_ready = q_122_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_8_io_bottom_out_ready = q_294_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_8_clock = clock;
  assign cols_3_8_reset = reset;
  assign cols_3_8_io_left_in_valid = q_122_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_3_8_io_left_in_bits = q_122_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_3_8_io_top_in_valid = q_308_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_3_8_io_top_in_bits = q_308_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_3_8_io_sum_ready = q_643_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_8_io_right_out_ready = q_123_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_8_io_bottom_out_ready = q_309_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_8_clock = clock;
  assign cols_4_8_reset = reset;
  assign cols_4_8_io_left_in_valid = q_123_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_4_8_io_left_in_bits = q_123_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_4_8_io_top_in_valid = q_323_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_4_8_io_top_in_bits = q_323_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_4_8_io_sum_ready = q_644_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_8_io_right_out_ready = q_124_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_8_io_bottom_out_ready = q_324_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_8_clock = clock;
  assign cols_5_8_reset = reset;
  assign cols_5_8_io_left_in_valid = q_124_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_5_8_io_left_in_bits = q_124_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_5_8_io_top_in_valid = q_338_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_5_8_io_top_in_bits = q_338_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_5_8_io_sum_ready = q_645_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_8_io_right_out_ready = q_125_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_8_io_bottom_out_ready = q_339_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_8_clock = clock;
  assign cols_6_8_reset = reset;
  assign cols_6_8_io_left_in_valid = q_125_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_6_8_io_left_in_bits = q_125_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_6_8_io_top_in_valid = q_353_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_6_8_io_top_in_bits = q_353_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_6_8_io_sum_ready = q_646_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_8_io_right_out_ready = q_126_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_8_io_bottom_out_ready = q_354_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_8_clock = clock;
  assign cols_7_8_reset = reset;
  assign cols_7_8_io_left_in_valid = q_126_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_7_8_io_left_in_bits = q_126_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_7_8_io_top_in_valid = q_368_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_7_8_io_top_in_bits = q_368_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_7_8_io_sum_ready = q_647_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_8_io_right_out_ready = q_127_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_8_io_bottom_out_ready = q_369_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_8_clock = clock;
  assign cols_8_8_reset = reset;
  assign cols_8_8_io_left_in_valid = q_127_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_8_8_io_left_in_bits = q_127_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_8_8_io_top_in_valid = q_383_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_8_8_io_top_in_bits = q_383_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_8_8_io_sum_ready = q_648_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_8_io_right_out_ready = q_128_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_8_io_bottom_out_ready = q_384_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_8_clock = clock;
  assign cols_9_8_reset = reset;
  assign cols_9_8_io_left_in_valid = q_128_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_9_8_io_left_in_bits = q_128_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_9_8_io_top_in_valid = q_398_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_9_8_io_top_in_bits = q_398_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_9_8_io_sum_ready = q_649_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_8_io_right_out_ready = q_129_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_8_io_bottom_out_ready = q_399_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_8_clock = clock;
  assign cols_10_8_reset = reset;
  assign cols_10_8_io_left_in_valid = q_129_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_10_8_io_left_in_bits = q_129_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_10_8_io_top_in_valid = q_413_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_10_8_io_top_in_bits = q_413_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_10_8_io_sum_ready = q_650_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_8_io_right_out_ready = q_130_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_8_io_bottom_out_ready = q_414_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_8_clock = clock;
  assign cols_11_8_reset = reset;
  assign cols_11_8_io_left_in_valid = q_130_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_11_8_io_left_in_bits = q_130_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_11_8_io_top_in_valid = q_428_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_11_8_io_top_in_bits = q_428_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_11_8_io_sum_ready = q_651_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_8_io_right_out_ready = q_131_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_8_io_bottom_out_ready = q_429_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_8_clock = clock;
  assign cols_12_8_reset = reset;
  assign cols_12_8_io_left_in_valid = q_131_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_12_8_io_left_in_bits = q_131_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_12_8_io_top_in_valid = q_443_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_12_8_io_top_in_bits = q_443_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_12_8_io_sum_ready = q_652_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_8_io_right_out_ready = q_132_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_8_io_bottom_out_ready = q_444_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_8_clock = clock;
  assign cols_13_8_reset = reset;
  assign cols_13_8_io_left_in_valid = q_132_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_13_8_io_left_in_bits = q_132_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_13_8_io_top_in_valid = q_458_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_13_8_io_top_in_bits = q_458_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_13_8_io_sum_ready = q_653_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_8_io_right_out_ready = q_133_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_8_io_bottom_out_ready = q_459_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_8_clock = clock;
  assign cols_14_8_reset = reset;
  assign cols_14_8_io_left_in_valid = q_133_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_14_8_io_left_in_bits = q_133_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_14_8_io_top_in_valid = q_473_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_14_8_io_top_in_bits = q_473_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_14_8_io_sum_ready = q_654_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_8_io_right_out_ready = q_134_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_8_io_bottom_out_ready = q_474_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_8_clock = clock;
  assign cols_15_8_reset = reset;
  assign cols_15_8_io_left_in_valid = q_134_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_15_8_io_left_in_bits = q_134_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_15_8_io_top_in_valid = q_488_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_15_8_io_top_in_bits = q_488_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_15_8_io_sum_ready = q_655_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_8_io_right_out_ready = 1'h1; // @[Stab.scala 102:51]
  assign cols_15_8_io_bottom_out_ready = q_489_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_9_clock = clock;
  assign cols_0_9_reset = reset;
  assign cols_0_9_io_left_in_valid = q_505_io_deq_valid; // @[Stab.scala 100:101]
  assign cols_0_9_io_left_in_bits = q_505_io_deq_bits; // @[Stab.scala 100:101]
  assign cols_0_9_io_top_in_valid = q_264_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_0_9_io_top_in_bits = q_264_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_0_9_io_sum_ready = q_656_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_9_io_right_out_ready = q_135_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_9_io_bottom_out_ready = q_265_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_9_clock = clock;
  assign cols_1_9_reset = reset;
  assign cols_1_9_io_left_in_valid = q_135_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_1_9_io_left_in_bits = q_135_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_1_9_io_top_in_valid = q_279_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_1_9_io_top_in_bits = q_279_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_1_9_io_sum_ready = q_657_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_9_io_right_out_ready = q_136_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_9_io_bottom_out_ready = q_280_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_9_clock = clock;
  assign cols_2_9_reset = reset;
  assign cols_2_9_io_left_in_valid = q_136_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_2_9_io_left_in_bits = q_136_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_2_9_io_top_in_valid = q_294_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_2_9_io_top_in_bits = q_294_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_2_9_io_sum_ready = q_658_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_9_io_right_out_ready = q_137_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_9_io_bottom_out_ready = q_295_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_9_clock = clock;
  assign cols_3_9_reset = reset;
  assign cols_3_9_io_left_in_valid = q_137_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_3_9_io_left_in_bits = q_137_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_3_9_io_top_in_valid = q_309_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_3_9_io_top_in_bits = q_309_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_3_9_io_sum_ready = q_659_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_9_io_right_out_ready = q_138_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_9_io_bottom_out_ready = q_310_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_9_clock = clock;
  assign cols_4_9_reset = reset;
  assign cols_4_9_io_left_in_valid = q_138_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_4_9_io_left_in_bits = q_138_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_4_9_io_top_in_valid = q_324_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_4_9_io_top_in_bits = q_324_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_4_9_io_sum_ready = q_660_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_9_io_right_out_ready = q_139_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_9_io_bottom_out_ready = q_325_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_9_clock = clock;
  assign cols_5_9_reset = reset;
  assign cols_5_9_io_left_in_valid = q_139_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_5_9_io_left_in_bits = q_139_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_5_9_io_top_in_valid = q_339_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_5_9_io_top_in_bits = q_339_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_5_9_io_sum_ready = q_661_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_9_io_right_out_ready = q_140_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_9_io_bottom_out_ready = q_340_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_9_clock = clock;
  assign cols_6_9_reset = reset;
  assign cols_6_9_io_left_in_valid = q_140_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_6_9_io_left_in_bits = q_140_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_6_9_io_top_in_valid = q_354_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_6_9_io_top_in_bits = q_354_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_6_9_io_sum_ready = q_662_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_9_io_right_out_ready = q_141_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_9_io_bottom_out_ready = q_355_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_9_clock = clock;
  assign cols_7_9_reset = reset;
  assign cols_7_9_io_left_in_valid = q_141_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_7_9_io_left_in_bits = q_141_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_7_9_io_top_in_valid = q_369_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_7_9_io_top_in_bits = q_369_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_7_9_io_sum_ready = q_663_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_9_io_right_out_ready = q_142_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_9_io_bottom_out_ready = q_370_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_9_clock = clock;
  assign cols_8_9_reset = reset;
  assign cols_8_9_io_left_in_valid = q_142_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_8_9_io_left_in_bits = q_142_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_8_9_io_top_in_valid = q_384_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_8_9_io_top_in_bits = q_384_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_8_9_io_sum_ready = q_664_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_9_io_right_out_ready = q_143_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_9_io_bottom_out_ready = q_385_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_9_clock = clock;
  assign cols_9_9_reset = reset;
  assign cols_9_9_io_left_in_valid = q_143_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_9_9_io_left_in_bits = q_143_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_9_9_io_top_in_valid = q_399_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_9_9_io_top_in_bits = q_399_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_9_9_io_sum_ready = q_665_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_9_io_right_out_ready = q_144_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_9_io_bottom_out_ready = q_400_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_9_clock = clock;
  assign cols_10_9_reset = reset;
  assign cols_10_9_io_left_in_valid = q_144_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_10_9_io_left_in_bits = q_144_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_10_9_io_top_in_valid = q_414_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_10_9_io_top_in_bits = q_414_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_10_9_io_sum_ready = q_666_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_9_io_right_out_ready = q_145_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_9_io_bottom_out_ready = q_415_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_9_clock = clock;
  assign cols_11_9_reset = reset;
  assign cols_11_9_io_left_in_valid = q_145_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_11_9_io_left_in_bits = q_145_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_11_9_io_top_in_valid = q_429_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_11_9_io_top_in_bits = q_429_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_11_9_io_sum_ready = q_667_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_9_io_right_out_ready = q_146_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_9_io_bottom_out_ready = q_430_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_9_clock = clock;
  assign cols_12_9_reset = reset;
  assign cols_12_9_io_left_in_valid = q_146_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_12_9_io_left_in_bits = q_146_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_12_9_io_top_in_valid = q_444_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_12_9_io_top_in_bits = q_444_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_12_9_io_sum_ready = q_668_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_9_io_right_out_ready = q_147_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_9_io_bottom_out_ready = q_445_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_9_clock = clock;
  assign cols_13_9_reset = reset;
  assign cols_13_9_io_left_in_valid = q_147_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_13_9_io_left_in_bits = q_147_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_13_9_io_top_in_valid = q_459_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_13_9_io_top_in_bits = q_459_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_13_9_io_sum_ready = q_669_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_9_io_right_out_ready = q_148_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_9_io_bottom_out_ready = q_460_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_9_clock = clock;
  assign cols_14_9_reset = reset;
  assign cols_14_9_io_left_in_valid = q_148_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_14_9_io_left_in_bits = q_148_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_14_9_io_top_in_valid = q_474_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_14_9_io_top_in_bits = q_474_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_14_9_io_sum_ready = q_670_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_9_io_right_out_ready = q_149_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_9_io_bottom_out_ready = q_475_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_9_clock = clock;
  assign cols_15_9_reset = reset;
  assign cols_15_9_io_left_in_valid = q_149_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_15_9_io_left_in_bits = q_149_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_15_9_io_top_in_valid = q_489_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_15_9_io_top_in_bits = q_489_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_15_9_io_sum_ready = q_671_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_9_io_right_out_ready = 1'h1; // @[Stab.scala 102:51]
  assign cols_15_9_io_bottom_out_ready = q_490_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_10_clock = clock;
  assign cols_0_10_reset = reset;
  assign cols_0_10_io_left_in_valid = q_506_io_deq_valid; // @[Stab.scala 100:101]
  assign cols_0_10_io_left_in_bits = q_506_io_deq_bits; // @[Stab.scala 100:101]
  assign cols_0_10_io_top_in_valid = q_265_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_0_10_io_top_in_bits = q_265_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_0_10_io_sum_ready = q_672_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_10_io_right_out_ready = q_150_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_10_io_bottom_out_ready = q_266_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_10_clock = clock;
  assign cols_1_10_reset = reset;
  assign cols_1_10_io_left_in_valid = q_150_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_1_10_io_left_in_bits = q_150_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_1_10_io_top_in_valid = q_280_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_1_10_io_top_in_bits = q_280_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_1_10_io_sum_ready = q_673_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_10_io_right_out_ready = q_151_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_10_io_bottom_out_ready = q_281_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_10_clock = clock;
  assign cols_2_10_reset = reset;
  assign cols_2_10_io_left_in_valid = q_151_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_2_10_io_left_in_bits = q_151_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_2_10_io_top_in_valid = q_295_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_2_10_io_top_in_bits = q_295_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_2_10_io_sum_ready = q_674_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_10_io_right_out_ready = q_152_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_10_io_bottom_out_ready = q_296_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_10_clock = clock;
  assign cols_3_10_reset = reset;
  assign cols_3_10_io_left_in_valid = q_152_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_3_10_io_left_in_bits = q_152_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_3_10_io_top_in_valid = q_310_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_3_10_io_top_in_bits = q_310_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_3_10_io_sum_ready = q_675_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_10_io_right_out_ready = q_153_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_10_io_bottom_out_ready = q_311_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_10_clock = clock;
  assign cols_4_10_reset = reset;
  assign cols_4_10_io_left_in_valid = q_153_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_4_10_io_left_in_bits = q_153_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_4_10_io_top_in_valid = q_325_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_4_10_io_top_in_bits = q_325_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_4_10_io_sum_ready = q_676_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_10_io_right_out_ready = q_154_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_10_io_bottom_out_ready = q_326_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_10_clock = clock;
  assign cols_5_10_reset = reset;
  assign cols_5_10_io_left_in_valid = q_154_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_5_10_io_left_in_bits = q_154_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_5_10_io_top_in_valid = q_340_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_5_10_io_top_in_bits = q_340_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_5_10_io_sum_ready = q_677_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_10_io_right_out_ready = q_155_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_10_io_bottom_out_ready = q_341_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_10_clock = clock;
  assign cols_6_10_reset = reset;
  assign cols_6_10_io_left_in_valid = q_155_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_6_10_io_left_in_bits = q_155_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_6_10_io_top_in_valid = q_355_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_6_10_io_top_in_bits = q_355_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_6_10_io_sum_ready = q_678_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_10_io_right_out_ready = q_156_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_10_io_bottom_out_ready = q_356_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_10_clock = clock;
  assign cols_7_10_reset = reset;
  assign cols_7_10_io_left_in_valid = q_156_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_7_10_io_left_in_bits = q_156_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_7_10_io_top_in_valid = q_370_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_7_10_io_top_in_bits = q_370_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_7_10_io_sum_ready = q_679_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_10_io_right_out_ready = q_157_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_10_io_bottom_out_ready = q_371_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_10_clock = clock;
  assign cols_8_10_reset = reset;
  assign cols_8_10_io_left_in_valid = q_157_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_8_10_io_left_in_bits = q_157_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_8_10_io_top_in_valid = q_385_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_8_10_io_top_in_bits = q_385_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_8_10_io_sum_ready = q_680_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_10_io_right_out_ready = q_158_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_10_io_bottom_out_ready = q_386_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_10_clock = clock;
  assign cols_9_10_reset = reset;
  assign cols_9_10_io_left_in_valid = q_158_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_9_10_io_left_in_bits = q_158_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_9_10_io_top_in_valid = q_400_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_9_10_io_top_in_bits = q_400_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_9_10_io_sum_ready = q_681_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_10_io_right_out_ready = q_159_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_10_io_bottom_out_ready = q_401_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_10_clock = clock;
  assign cols_10_10_reset = reset;
  assign cols_10_10_io_left_in_valid = q_159_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_10_10_io_left_in_bits = q_159_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_10_10_io_top_in_valid = q_415_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_10_10_io_top_in_bits = q_415_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_10_10_io_sum_ready = q_682_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_10_io_right_out_ready = q_160_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_10_io_bottom_out_ready = q_416_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_10_clock = clock;
  assign cols_11_10_reset = reset;
  assign cols_11_10_io_left_in_valid = q_160_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_11_10_io_left_in_bits = q_160_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_11_10_io_top_in_valid = q_430_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_11_10_io_top_in_bits = q_430_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_11_10_io_sum_ready = q_683_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_10_io_right_out_ready = q_161_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_10_io_bottom_out_ready = q_431_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_10_clock = clock;
  assign cols_12_10_reset = reset;
  assign cols_12_10_io_left_in_valid = q_161_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_12_10_io_left_in_bits = q_161_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_12_10_io_top_in_valid = q_445_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_12_10_io_top_in_bits = q_445_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_12_10_io_sum_ready = q_684_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_10_io_right_out_ready = q_162_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_10_io_bottom_out_ready = q_446_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_10_clock = clock;
  assign cols_13_10_reset = reset;
  assign cols_13_10_io_left_in_valid = q_162_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_13_10_io_left_in_bits = q_162_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_13_10_io_top_in_valid = q_460_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_13_10_io_top_in_bits = q_460_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_13_10_io_sum_ready = q_685_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_10_io_right_out_ready = q_163_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_10_io_bottom_out_ready = q_461_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_10_clock = clock;
  assign cols_14_10_reset = reset;
  assign cols_14_10_io_left_in_valid = q_163_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_14_10_io_left_in_bits = q_163_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_14_10_io_top_in_valid = q_475_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_14_10_io_top_in_bits = q_475_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_14_10_io_sum_ready = q_686_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_10_io_right_out_ready = q_164_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_10_io_bottom_out_ready = q_476_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_10_clock = clock;
  assign cols_15_10_reset = reset;
  assign cols_15_10_io_left_in_valid = q_164_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_15_10_io_left_in_bits = q_164_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_15_10_io_top_in_valid = q_490_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_15_10_io_top_in_bits = q_490_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_15_10_io_sum_ready = q_687_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_10_io_right_out_ready = 1'h1; // @[Stab.scala 102:51]
  assign cols_15_10_io_bottom_out_ready = q_491_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_11_clock = clock;
  assign cols_0_11_reset = reset;
  assign cols_0_11_io_left_in_valid = q_507_io_deq_valid; // @[Stab.scala 100:101]
  assign cols_0_11_io_left_in_bits = q_507_io_deq_bits; // @[Stab.scala 100:101]
  assign cols_0_11_io_top_in_valid = q_266_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_0_11_io_top_in_bits = q_266_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_0_11_io_sum_ready = q_688_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_11_io_right_out_ready = q_165_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_11_io_bottom_out_ready = q_267_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_11_clock = clock;
  assign cols_1_11_reset = reset;
  assign cols_1_11_io_left_in_valid = q_165_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_1_11_io_left_in_bits = q_165_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_1_11_io_top_in_valid = q_281_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_1_11_io_top_in_bits = q_281_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_1_11_io_sum_ready = q_689_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_11_io_right_out_ready = q_166_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_11_io_bottom_out_ready = q_282_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_11_clock = clock;
  assign cols_2_11_reset = reset;
  assign cols_2_11_io_left_in_valid = q_166_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_2_11_io_left_in_bits = q_166_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_2_11_io_top_in_valid = q_296_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_2_11_io_top_in_bits = q_296_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_2_11_io_sum_ready = q_690_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_11_io_right_out_ready = q_167_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_11_io_bottom_out_ready = q_297_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_11_clock = clock;
  assign cols_3_11_reset = reset;
  assign cols_3_11_io_left_in_valid = q_167_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_3_11_io_left_in_bits = q_167_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_3_11_io_top_in_valid = q_311_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_3_11_io_top_in_bits = q_311_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_3_11_io_sum_ready = q_691_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_11_io_right_out_ready = q_168_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_11_io_bottom_out_ready = q_312_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_11_clock = clock;
  assign cols_4_11_reset = reset;
  assign cols_4_11_io_left_in_valid = q_168_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_4_11_io_left_in_bits = q_168_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_4_11_io_top_in_valid = q_326_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_4_11_io_top_in_bits = q_326_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_4_11_io_sum_ready = q_692_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_11_io_right_out_ready = q_169_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_11_io_bottom_out_ready = q_327_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_11_clock = clock;
  assign cols_5_11_reset = reset;
  assign cols_5_11_io_left_in_valid = q_169_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_5_11_io_left_in_bits = q_169_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_5_11_io_top_in_valid = q_341_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_5_11_io_top_in_bits = q_341_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_5_11_io_sum_ready = q_693_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_11_io_right_out_ready = q_170_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_11_io_bottom_out_ready = q_342_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_11_clock = clock;
  assign cols_6_11_reset = reset;
  assign cols_6_11_io_left_in_valid = q_170_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_6_11_io_left_in_bits = q_170_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_6_11_io_top_in_valid = q_356_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_6_11_io_top_in_bits = q_356_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_6_11_io_sum_ready = q_694_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_11_io_right_out_ready = q_171_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_11_io_bottom_out_ready = q_357_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_11_clock = clock;
  assign cols_7_11_reset = reset;
  assign cols_7_11_io_left_in_valid = q_171_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_7_11_io_left_in_bits = q_171_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_7_11_io_top_in_valid = q_371_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_7_11_io_top_in_bits = q_371_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_7_11_io_sum_ready = q_695_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_11_io_right_out_ready = q_172_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_11_io_bottom_out_ready = q_372_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_11_clock = clock;
  assign cols_8_11_reset = reset;
  assign cols_8_11_io_left_in_valid = q_172_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_8_11_io_left_in_bits = q_172_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_8_11_io_top_in_valid = q_386_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_8_11_io_top_in_bits = q_386_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_8_11_io_sum_ready = q_696_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_11_io_right_out_ready = q_173_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_11_io_bottom_out_ready = q_387_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_11_clock = clock;
  assign cols_9_11_reset = reset;
  assign cols_9_11_io_left_in_valid = q_173_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_9_11_io_left_in_bits = q_173_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_9_11_io_top_in_valid = q_401_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_9_11_io_top_in_bits = q_401_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_9_11_io_sum_ready = q_697_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_11_io_right_out_ready = q_174_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_11_io_bottom_out_ready = q_402_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_11_clock = clock;
  assign cols_10_11_reset = reset;
  assign cols_10_11_io_left_in_valid = q_174_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_10_11_io_left_in_bits = q_174_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_10_11_io_top_in_valid = q_416_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_10_11_io_top_in_bits = q_416_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_10_11_io_sum_ready = q_698_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_11_io_right_out_ready = q_175_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_11_io_bottom_out_ready = q_417_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_11_clock = clock;
  assign cols_11_11_reset = reset;
  assign cols_11_11_io_left_in_valid = q_175_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_11_11_io_left_in_bits = q_175_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_11_11_io_top_in_valid = q_431_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_11_11_io_top_in_bits = q_431_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_11_11_io_sum_ready = q_699_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_11_io_right_out_ready = q_176_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_11_io_bottom_out_ready = q_432_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_11_clock = clock;
  assign cols_12_11_reset = reset;
  assign cols_12_11_io_left_in_valid = q_176_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_12_11_io_left_in_bits = q_176_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_12_11_io_top_in_valid = q_446_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_12_11_io_top_in_bits = q_446_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_12_11_io_sum_ready = q_700_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_11_io_right_out_ready = q_177_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_11_io_bottom_out_ready = q_447_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_11_clock = clock;
  assign cols_13_11_reset = reset;
  assign cols_13_11_io_left_in_valid = q_177_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_13_11_io_left_in_bits = q_177_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_13_11_io_top_in_valid = q_461_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_13_11_io_top_in_bits = q_461_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_13_11_io_sum_ready = q_701_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_11_io_right_out_ready = q_178_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_11_io_bottom_out_ready = q_462_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_11_clock = clock;
  assign cols_14_11_reset = reset;
  assign cols_14_11_io_left_in_valid = q_178_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_14_11_io_left_in_bits = q_178_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_14_11_io_top_in_valid = q_476_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_14_11_io_top_in_bits = q_476_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_14_11_io_sum_ready = q_702_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_11_io_right_out_ready = q_179_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_11_io_bottom_out_ready = q_477_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_11_clock = clock;
  assign cols_15_11_reset = reset;
  assign cols_15_11_io_left_in_valid = q_179_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_15_11_io_left_in_bits = q_179_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_15_11_io_top_in_valid = q_491_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_15_11_io_top_in_bits = q_491_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_15_11_io_sum_ready = q_703_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_11_io_right_out_ready = 1'h1; // @[Stab.scala 102:51]
  assign cols_15_11_io_bottom_out_ready = q_492_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_12_clock = clock;
  assign cols_0_12_reset = reset;
  assign cols_0_12_io_left_in_valid = q_508_io_deq_valid; // @[Stab.scala 100:101]
  assign cols_0_12_io_left_in_bits = q_508_io_deq_bits; // @[Stab.scala 100:101]
  assign cols_0_12_io_top_in_valid = q_267_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_0_12_io_top_in_bits = q_267_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_0_12_io_sum_ready = q_704_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_12_io_right_out_ready = q_180_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_12_io_bottom_out_ready = q_268_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_12_clock = clock;
  assign cols_1_12_reset = reset;
  assign cols_1_12_io_left_in_valid = q_180_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_1_12_io_left_in_bits = q_180_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_1_12_io_top_in_valid = q_282_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_1_12_io_top_in_bits = q_282_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_1_12_io_sum_ready = q_705_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_12_io_right_out_ready = q_181_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_12_io_bottom_out_ready = q_283_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_12_clock = clock;
  assign cols_2_12_reset = reset;
  assign cols_2_12_io_left_in_valid = q_181_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_2_12_io_left_in_bits = q_181_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_2_12_io_top_in_valid = q_297_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_2_12_io_top_in_bits = q_297_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_2_12_io_sum_ready = q_706_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_12_io_right_out_ready = q_182_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_12_io_bottom_out_ready = q_298_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_12_clock = clock;
  assign cols_3_12_reset = reset;
  assign cols_3_12_io_left_in_valid = q_182_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_3_12_io_left_in_bits = q_182_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_3_12_io_top_in_valid = q_312_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_3_12_io_top_in_bits = q_312_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_3_12_io_sum_ready = q_707_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_12_io_right_out_ready = q_183_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_12_io_bottom_out_ready = q_313_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_12_clock = clock;
  assign cols_4_12_reset = reset;
  assign cols_4_12_io_left_in_valid = q_183_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_4_12_io_left_in_bits = q_183_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_4_12_io_top_in_valid = q_327_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_4_12_io_top_in_bits = q_327_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_4_12_io_sum_ready = q_708_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_12_io_right_out_ready = q_184_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_12_io_bottom_out_ready = q_328_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_12_clock = clock;
  assign cols_5_12_reset = reset;
  assign cols_5_12_io_left_in_valid = q_184_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_5_12_io_left_in_bits = q_184_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_5_12_io_top_in_valid = q_342_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_5_12_io_top_in_bits = q_342_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_5_12_io_sum_ready = q_709_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_12_io_right_out_ready = q_185_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_12_io_bottom_out_ready = q_343_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_12_clock = clock;
  assign cols_6_12_reset = reset;
  assign cols_6_12_io_left_in_valid = q_185_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_6_12_io_left_in_bits = q_185_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_6_12_io_top_in_valid = q_357_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_6_12_io_top_in_bits = q_357_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_6_12_io_sum_ready = q_710_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_12_io_right_out_ready = q_186_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_12_io_bottom_out_ready = q_358_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_12_clock = clock;
  assign cols_7_12_reset = reset;
  assign cols_7_12_io_left_in_valid = q_186_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_7_12_io_left_in_bits = q_186_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_7_12_io_top_in_valid = q_372_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_7_12_io_top_in_bits = q_372_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_7_12_io_sum_ready = q_711_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_12_io_right_out_ready = q_187_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_12_io_bottom_out_ready = q_373_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_12_clock = clock;
  assign cols_8_12_reset = reset;
  assign cols_8_12_io_left_in_valid = q_187_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_8_12_io_left_in_bits = q_187_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_8_12_io_top_in_valid = q_387_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_8_12_io_top_in_bits = q_387_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_8_12_io_sum_ready = q_712_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_12_io_right_out_ready = q_188_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_12_io_bottom_out_ready = q_388_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_12_clock = clock;
  assign cols_9_12_reset = reset;
  assign cols_9_12_io_left_in_valid = q_188_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_9_12_io_left_in_bits = q_188_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_9_12_io_top_in_valid = q_402_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_9_12_io_top_in_bits = q_402_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_9_12_io_sum_ready = q_713_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_12_io_right_out_ready = q_189_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_12_io_bottom_out_ready = q_403_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_12_clock = clock;
  assign cols_10_12_reset = reset;
  assign cols_10_12_io_left_in_valid = q_189_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_10_12_io_left_in_bits = q_189_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_10_12_io_top_in_valid = q_417_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_10_12_io_top_in_bits = q_417_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_10_12_io_sum_ready = q_714_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_12_io_right_out_ready = q_190_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_12_io_bottom_out_ready = q_418_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_12_clock = clock;
  assign cols_11_12_reset = reset;
  assign cols_11_12_io_left_in_valid = q_190_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_11_12_io_left_in_bits = q_190_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_11_12_io_top_in_valid = q_432_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_11_12_io_top_in_bits = q_432_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_11_12_io_sum_ready = q_715_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_12_io_right_out_ready = q_191_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_12_io_bottom_out_ready = q_433_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_12_clock = clock;
  assign cols_12_12_reset = reset;
  assign cols_12_12_io_left_in_valid = q_191_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_12_12_io_left_in_bits = q_191_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_12_12_io_top_in_valid = q_447_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_12_12_io_top_in_bits = q_447_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_12_12_io_sum_ready = q_716_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_12_io_right_out_ready = q_192_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_12_io_bottom_out_ready = q_448_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_12_clock = clock;
  assign cols_13_12_reset = reset;
  assign cols_13_12_io_left_in_valid = q_192_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_13_12_io_left_in_bits = q_192_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_13_12_io_top_in_valid = q_462_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_13_12_io_top_in_bits = q_462_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_13_12_io_sum_ready = q_717_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_12_io_right_out_ready = q_193_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_12_io_bottom_out_ready = q_463_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_12_clock = clock;
  assign cols_14_12_reset = reset;
  assign cols_14_12_io_left_in_valid = q_193_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_14_12_io_left_in_bits = q_193_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_14_12_io_top_in_valid = q_477_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_14_12_io_top_in_bits = q_477_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_14_12_io_sum_ready = q_718_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_12_io_right_out_ready = q_194_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_12_io_bottom_out_ready = q_478_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_12_clock = clock;
  assign cols_15_12_reset = reset;
  assign cols_15_12_io_left_in_valid = q_194_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_15_12_io_left_in_bits = q_194_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_15_12_io_top_in_valid = q_492_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_15_12_io_top_in_bits = q_492_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_15_12_io_sum_ready = q_719_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_12_io_right_out_ready = 1'h1; // @[Stab.scala 102:51]
  assign cols_15_12_io_bottom_out_ready = q_493_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_13_clock = clock;
  assign cols_0_13_reset = reset;
  assign cols_0_13_io_left_in_valid = q_509_io_deq_valid; // @[Stab.scala 100:101]
  assign cols_0_13_io_left_in_bits = q_509_io_deq_bits; // @[Stab.scala 100:101]
  assign cols_0_13_io_top_in_valid = q_268_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_0_13_io_top_in_bits = q_268_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_0_13_io_sum_ready = q_720_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_13_io_right_out_ready = q_195_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_13_io_bottom_out_ready = q_269_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_13_clock = clock;
  assign cols_1_13_reset = reset;
  assign cols_1_13_io_left_in_valid = q_195_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_1_13_io_left_in_bits = q_195_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_1_13_io_top_in_valid = q_283_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_1_13_io_top_in_bits = q_283_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_1_13_io_sum_ready = q_721_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_13_io_right_out_ready = q_196_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_13_io_bottom_out_ready = q_284_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_13_clock = clock;
  assign cols_2_13_reset = reset;
  assign cols_2_13_io_left_in_valid = q_196_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_2_13_io_left_in_bits = q_196_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_2_13_io_top_in_valid = q_298_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_2_13_io_top_in_bits = q_298_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_2_13_io_sum_ready = q_722_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_13_io_right_out_ready = q_197_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_13_io_bottom_out_ready = q_299_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_13_clock = clock;
  assign cols_3_13_reset = reset;
  assign cols_3_13_io_left_in_valid = q_197_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_3_13_io_left_in_bits = q_197_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_3_13_io_top_in_valid = q_313_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_3_13_io_top_in_bits = q_313_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_3_13_io_sum_ready = q_723_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_13_io_right_out_ready = q_198_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_13_io_bottom_out_ready = q_314_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_13_clock = clock;
  assign cols_4_13_reset = reset;
  assign cols_4_13_io_left_in_valid = q_198_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_4_13_io_left_in_bits = q_198_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_4_13_io_top_in_valid = q_328_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_4_13_io_top_in_bits = q_328_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_4_13_io_sum_ready = q_724_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_13_io_right_out_ready = q_199_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_13_io_bottom_out_ready = q_329_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_13_clock = clock;
  assign cols_5_13_reset = reset;
  assign cols_5_13_io_left_in_valid = q_199_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_5_13_io_left_in_bits = q_199_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_5_13_io_top_in_valid = q_343_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_5_13_io_top_in_bits = q_343_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_5_13_io_sum_ready = q_725_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_13_io_right_out_ready = q_200_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_13_io_bottom_out_ready = q_344_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_13_clock = clock;
  assign cols_6_13_reset = reset;
  assign cols_6_13_io_left_in_valid = q_200_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_6_13_io_left_in_bits = q_200_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_6_13_io_top_in_valid = q_358_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_6_13_io_top_in_bits = q_358_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_6_13_io_sum_ready = q_726_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_13_io_right_out_ready = q_201_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_13_io_bottom_out_ready = q_359_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_13_clock = clock;
  assign cols_7_13_reset = reset;
  assign cols_7_13_io_left_in_valid = q_201_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_7_13_io_left_in_bits = q_201_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_7_13_io_top_in_valid = q_373_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_7_13_io_top_in_bits = q_373_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_7_13_io_sum_ready = q_727_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_13_io_right_out_ready = q_202_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_13_io_bottom_out_ready = q_374_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_13_clock = clock;
  assign cols_8_13_reset = reset;
  assign cols_8_13_io_left_in_valid = q_202_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_8_13_io_left_in_bits = q_202_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_8_13_io_top_in_valid = q_388_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_8_13_io_top_in_bits = q_388_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_8_13_io_sum_ready = q_728_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_13_io_right_out_ready = q_203_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_13_io_bottom_out_ready = q_389_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_13_clock = clock;
  assign cols_9_13_reset = reset;
  assign cols_9_13_io_left_in_valid = q_203_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_9_13_io_left_in_bits = q_203_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_9_13_io_top_in_valid = q_403_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_9_13_io_top_in_bits = q_403_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_9_13_io_sum_ready = q_729_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_13_io_right_out_ready = q_204_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_13_io_bottom_out_ready = q_404_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_13_clock = clock;
  assign cols_10_13_reset = reset;
  assign cols_10_13_io_left_in_valid = q_204_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_10_13_io_left_in_bits = q_204_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_10_13_io_top_in_valid = q_418_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_10_13_io_top_in_bits = q_418_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_10_13_io_sum_ready = q_730_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_13_io_right_out_ready = q_205_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_13_io_bottom_out_ready = q_419_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_13_clock = clock;
  assign cols_11_13_reset = reset;
  assign cols_11_13_io_left_in_valid = q_205_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_11_13_io_left_in_bits = q_205_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_11_13_io_top_in_valid = q_433_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_11_13_io_top_in_bits = q_433_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_11_13_io_sum_ready = q_731_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_13_io_right_out_ready = q_206_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_13_io_bottom_out_ready = q_434_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_13_clock = clock;
  assign cols_12_13_reset = reset;
  assign cols_12_13_io_left_in_valid = q_206_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_12_13_io_left_in_bits = q_206_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_12_13_io_top_in_valid = q_448_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_12_13_io_top_in_bits = q_448_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_12_13_io_sum_ready = q_732_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_13_io_right_out_ready = q_207_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_13_io_bottom_out_ready = q_449_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_13_clock = clock;
  assign cols_13_13_reset = reset;
  assign cols_13_13_io_left_in_valid = q_207_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_13_13_io_left_in_bits = q_207_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_13_13_io_top_in_valid = q_463_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_13_13_io_top_in_bits = q_463_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_13_13_io_sum_ready = q_733_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_13_io_right_out_ready = q_208_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_13_io_bottom_out_ready = q_464_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_13_clock = clock;
  assign cols_14_13_reset = reset;
  assign cols_14_13_io_left_in_valid = q_208_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_14_13_io_left_in_bits = q_208_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_14_13_io_top_in_valid = q_478_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_14_13_io_top_in_bits = q_478_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_14_13_io_sum_ready = q_734_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_13_io_right_out_ready = q_209_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_13_io_bottom_out_ready = q_479_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_13_clock = clock;
  assign cols_15_13_reset = reset;
  assign cols_15_13_io_left_in_valid = q_209_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_15_13_io_left_in_bits = q_209_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_15_13_io_top_in_valid = q_493_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_15_13_io_top_in_bits = q_493_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_15_13_io_sum_ready = q_735_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_13_io_right_out_ready = 1'h1; // @[Stab.scala 102:51]
  assign cols_15_13_io_bottom_out_ready = q_494_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_14_clock = clock;
  assign cols_0_14_reset = reset;
  assign cols_0_14_io_left_in_valid = q_510_io_deq_valid; // @[Stab.scala 100:101]
  assign cols_0_14_io_left_in_bits = q_510_io_deq_bits; // @[Stab.scala 100:101]
  assign cols_0_14_io_top_in_valid = q_269_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_0_14_io_top_in_bits = q_269_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_0_14_io_sum_ready = q_736_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_14_io_right_out_ready = q_210_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_14_io_bottom_out_ready = q_270_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_14_clock = clock;
  assign cols_1_14_reset = reset;
  assign cols_1_14_io_left_in_valid = q_210_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_1_14_io_left_in_bits = q_210_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_1_14_io_top_in_valid = q_284_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_1_14_io_top_in_bits = q_284_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_1_14_io_sum_ready = q_737_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_14_io_right_out_ready = q_211_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_14_io_bottom_out_ready = q_285_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_14_clock = clock;
  assign cols_2_14_reset = reset;
  assign cols_2_14_io_left_in_valid = q_211_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_2_14_io_left_in_bits = q_211_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_2_14_io_top_in_valid = q_299_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_2_14_io_top_in_bits = q_299_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_2_14_io_sum_ready = q_738_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_14_io_right_out_ready = q_212_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_14_io_bottom_out_ready = q_300_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_14_clock = clock;
  assign cols_3_14_reset = reset;
  assign cols_3_14_io_left_in_valid = q_212_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_3_14_io_left_in_bits = q_212_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_3_14_io_top_in_valid = q_314_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_3_14_io_top_in_bits = q_314_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_3_14_io_sum_ready = q_739_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_14_io_right_out_ready = q_213_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_14_io_bottom_out_ready = q_315_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_14_clock = clock;
  assign cols_4_14_reset = reset;
  assign cols_4_14_io_left_in_valid = q_213_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_4_14_io_left_in_bits = q_213_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_4_14_io_top_in_valid = q_329_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_4_14_io_top_in_bits = q_329_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_4_14_io_sum_ready = q_740_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_14_io_right_out_ready = q_214_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_14_io_bottom_out_ready = q_330_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_14_clock = clock;
  assign cols_5_14_reset = reset;
  assign cols_5_14_io_left_in_valid = q_214_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_5_14_io_left_in_bits = q_214_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_5_14_io_top_in_valid = q_344_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_5_14_io_top_in_bits = q_344_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_5_14_io_sum_ready = q_741_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_14_io_right_out_ready = q_215_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_14_io_bottom_out_ready = q_345_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_14_clock = clock;
  assign cols_6_14_reset = reset;
  assign cols_6_14_io_left_in_valid = q_215_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_6_14_io_left_in_bits = q_215_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_6_14_io_top_in_valid = q_359_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_6_14_io_top_in_bits = q_359_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_6_14_io_sum_ready = q_742_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_14_io_right_out_ready = q_216_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_14_io_bottom_out_ready = q_360_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_14_clock = clock;
  assign cols_7_14_reset = reset;
  assign cols_7_14_io_left_in_valid = q_216_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_7_14_io_left_in_bits = q_216_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_7_14_io_top_in_valid = q_374_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_7_14_io_top_in_bits = q_374_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_7_14_io_sum_ready = q_743_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_14_io_right_out_ready = q_217_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_14_io_bottom_out_ready = q_375_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_14_clock = clock;
  assign cols_8_14_reset = reset;
  assign cols_8_14_io_left_in_valid = q_217_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_8_14_io_left_in_bits = q_217_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_8_14_io_top_in_valid = q_389_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_8_14_io_top_in_bits = q_389_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_8_14_io_sum_ready = q_744_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_14_io_right_out_ready = q_218_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_14_io_bottom_out_ready = q_390_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_14_clock = clock;
  assign cols_9_14_reset = reset;
  assign cols_9_14_io_left_in_valid = q_218_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_9_14_io_left_in_bits = q_218_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_9_14_io_top_in_valid = q_404_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_9_14_io_top_in_bits = q_404_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_9_14_io_sum_ready = q_745_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_14_io_right_out_ready = q_219_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_14_io_bottom_out_ready = q_405_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_14_clock = clock;
  assign cols_10_14_reset = reset;
  assign cols_10_14_io_left_in_valid = q_219_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_10_14_io_left_in_bits = q_219_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_10_14_io_top_in_valid = q_419_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_10_14_io_top_in_bits = q_419_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_10_14_io_sum_ready = q_746_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_14_io_right_out_ready = q_220_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_14_io_bottom_out_ready = q_420_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_14_clock = clock;
  assign cols_11_14_reset = reset;
  assign cols_11_14_io_left_in_valid = q_220_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_11_14_io_left_in_bits = q_220_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_11_14_io_top_in_valid = q_434_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_11_14_io_top_in_bits = q_434_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_11_14_io_sum_ready = q_747_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_14_io_right_out_ready = q_221_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_14_io_bottom_out_ready = q_435_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_14_clock = clock;
  assign cols_12_14_reset = reset;
  assign cols_12_14_io_left_in_valid = q_221_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_12_14_io_left_in_bits = q_221_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_12_14_io_top_in_valid = q_449_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_12_14_io_top_in_bits = q_449_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_12_14_io_sum_ready = q_748_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_14_io_right_out_ready = q_222_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_14_io_bottom_out_ready = q_450_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_14_clock = clock;
  assign cols_13_14_reset = reset;
  assign cols_13_14_io_left_in_valid = q_222_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_13_14_io_left_in_bits = q_222_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_13_14_io_top_in_valid = q_464_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_13_14_io_top_in_bits = q_464_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_13_14_io_sum_ready = q_749_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_14_io_right_out_ready = q_223_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_14_io_bottom_out_ready = q_465_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_14_clock = clock;
  assign cols_14_14_reset = reset;
  assign cols_14_14_io_left_in_valid = q_223_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_14_14_io_left_in_bits = q_223_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_14_14_io_top_in_valid = q_479_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_14_14_io_top_in_bits = q_479_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_14_14_io_sum_ready = q_750_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_14_io_right_out_ready = q_224_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_14_io_bottom_out_ready = q_480_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_14_clock = clock;
  assign cols_15_14_reset = reset;
  assign cols_15_14_io_left_in_valid = q_224_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_15_14_io_left_in_bits = q_224_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_15_14_io_top_in_valid = q_494_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_15_14_io_top_in_bits = q_494_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_15_14_io_sum_ready = q_751_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_14_io_right_out_ready = 1'h1; // @[Stab.scala 102:51]
  assign cols_15_14_io_bottom_out_ready = q_495_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_15_clock = clock;
  assign cols_0_15_reset = reset;
  assign cols_0_15_io_left_in_valid = q_511_io_deq_valid; // @[Stab.scala 100:101]
  assign cols_0_15_io_left_in_bits = q_511_io_deq_bits; // @[Stab.scala 100:101]
  assign cols_0_15_io_top_in_valid = q_270_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_0_15_io_top_in_bits = q_270_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_0_15_io_sum_ready = q_752_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_15_io_right_out_ready = q_225_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_0_15_io_bottom_out_ready = 1'h1; // @[Stab.scala 94:52]
  assign cols_1_15_clock = clock;
  assign cols_1_15_reset = reset;
  assign cols_1_15_io_left_in_valid = q_225_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_1_15_io_left_in_bits = q_225_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_1_15_io_top_in_valid = q_285_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_1_15_io_top_in_bits = q_285_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_1_15_io_sum_ready = q_753_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_15_io_right_out_ready = q_226_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_1_15_io_bottom_out_ready = 1'h1; // @[Stab.scala 94:52]
  assign cols_2_15_clock = clock;
  assign cols_2_15_reset = reset;
  assign cols_2_15_io_left_in_valid = q_226_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_2_15_io_left_in_bits = q_226_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_2_15_io_top_in_valid = q_300_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_2_15_io_top_in_bits = q_300_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_2_15_io_sum_ready = q_754_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_15_io_right_out_ready = q_227_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_2_15_io_bottom_out_ready = 1'h1; // @[Stab.scala 94:52]
  assign cols_3_15_clock = clock;
  assign cols_3_15_reset = reset;
  assign cols_3_15_io_left_in_valid = q_227_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_3_15_io_left_in_bits = q_227_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_3_15_io_top_in_valid = q_315_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_3_15_io_top_in_bits = q_315_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_3_15_io_sum_ready = q_755_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_15_io_right_out_ready = q_228_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_3_15_io_bottom_out_ready = 1'h1; // @[Stab.scala 94:52]
  assign cols_4_15_clock = clock;
  assign cols_4_15_reset = reset;
  assign cols_4_15_io_left_in_valid = q_228_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_4_15_io_left_in_bits = q_228_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_4_15_io_top_in_valid = q_330_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_4_15_io_top_in_bits = q_330_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_4_15_io_sum_ready = q_756_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_15_io_right_out_ready = q_229_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_4_15_io_bottom_out_ready = 1'h1; // @[Stab.scala 94:52]
  assign cols_5_15_clock = clock;
  assign cols_5_15_reset = reset;
  assign cols_5_15_io_left_in_valid = q_229_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_5_15_io_left_in_bits = q_229_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_5_15_io_top_in_valid = q_345_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_5_15_io_top_in_bits = q_345_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_5_15_io_sum_ready = q_757_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_15_io_right_out_ready = q_230_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_5_15_io_bottom_out_ready = 1'h1; // @[Stab.scala 94:52]
  assign cols_6_15_clock = clock;
  assign cols_6_15_reset = reset;
  assign cols_6_15_io_left_in_valid = q_230_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_6_15_io_left_in_bits = q_230_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_6_15_io_top_in_valid = q_360_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_6_15_io_top_in_bits = q_360_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_6_15_io_sum_ready = q_758_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_15_io_right_out_ready = q_231_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_6_15_io_bottom_out_ready = 1'h1; // @[Stab.scala 94:52]
  assign cols_7_15_clock = clock;
  assign cols_7_15_reset = reset;
  assign cols_7_15_io_left_in_valid = q_231_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_7_15_io_left_in_bits = q_231_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_7_15_io_top_in_valid = q_375_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_7_15_io_top_in_bits = q_375_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_7_15_io_sum_ready = q_759_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_15_io_right_out_ready = q_232_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_7_15_io_bottom_out_ready = 1'h1; // @[Stab.scala 94:52]
  assign cols_8_15_clock = clock;
  assign cols_8_15_reset = reset;
  assign cols_8_15_io_left_in_valid = q_232_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_8_15_io_left_in_bits = q_232_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_8_15_io_top_in_valid = q_390_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_8_15_io_top_in_bits = q_390_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_8_15_io_sum_ready = q_760_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_15_io_right_out_ready = q_233_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_8_15_io_bottom_out_ready = 1'h1; // @[Stab.scala 94:52]
  assign cols_9_15_clock = clock;
  assign cols_9_15_reset = reset;
  assign cols_9_15_io_left_in_valid = q_233_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_9_15_io_left_in_bits = q_233_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_9_15_io_top_in_valid = q_405_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_9_15_io_top_in_bits = q_405_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_9_15_io_sum_ready = q_761_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_15_io_right_out_ready = q_234_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_9_15_io_bottom_out_ready = 1'h1; // @[Stab.scala 94:52]
  assign cols_10_15_clock = clock;
  assign cols_10_15_reset = reset;
  assign cols_10_15_io_left_in_valid = q_234_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_10_15_io_left_in_bits = q_234_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_10_15_io_top_in_valid = q_420_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_10_15_io_top_in_bits = q_420_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_10_15_io_sum_ready = q_762_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_15_io_right_out_ready = q_235_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_10_15_io_bottom_out_ready = 1'h1; // @[Stab.scala 94:52]
  assign cols_11_15_clock = clock;
  assign cols_11_15_reset = reset;
  assign cols_11_15_io_left_in_valid = q_235_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_11_15_io_left_in_bits = q_235_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_11_15_io_top_in_valid = q_435_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_11_15_io_top_in_bits = q_435_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_11_15_io_sum_ready = q_763_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_15_io_right_out_ready = q_236_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_11_15_io_bottom_out_ready = 1'h1; // @[Stab.scala 94:52]
  assign cols_12_15_clock = clock;
  assign cols_12_15_reset = reset;
  assign cols_12_15_io_left_in_valid = q_236_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_12_15_io_left_in_bits = q_236_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_12_15_io_top_in_valid = q_450_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_12_15_io_top_in_bits = q_450_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_12_15_io_sum_ready = q_764_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_15_io_right_out_ready = q_237_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_12_15_io_bottom_out_ready = 1'h1; // @[Stab.scala 94:52]
  assign cols_13_15_clock = clock;
  assign cols_13_15_reset = reset;
  assign cols_13_15_io_left_in_valid = q_237_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_13_15_io_left_in_bits = q_237_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_13_15_io_top_in_valid = q_465_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_13_15_io_top_in_bits = q_465_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_13_15_io_sum_ready = q_765_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_15_io_right_out_ready = q_238_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_13_15_io_bottom_out_ready = 1'h1; // @[Stab.scala 94:52]
  assign cols_14_15_clock = clock;
  assign cols_14_15_reset = reset;
  assign cols_14_15_io_left_in_valid = q_238_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_14_15_io_left_in_bits = q_238_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_14_15_io_top_in_valid = q_480_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_14_15_io_top_in_bits = q_480_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_14_15_io_sum_ready = q_766_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_15_io_right_out_ready = q_239_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_14_15_io_bottom_out_ready = 1'h1; // @[Stab.scala 94:52]
  assign cols_15_15_clock = clock;
  assign cols_15_15_reset = reset;
  assign cols_15_15_io_left_in_valid = q_239_io_deq_valid; // @[Stab.scala 89:69]
  assign cols_15_15_io_left_in_bits = q_239_io_deq_bits; // @[Stab.scala 89:69]
  assign cols_15_15_io_top_in_valid = q_495_io_deq_valid; // @[Stab.scala 97:70]
  assign cols_15_15_io_top_in_bits = q_495_io_deq_bits; // @[Stab.scala 97:70]
  assign cols_15_15_io_sum_ready = q_767_io_enq_ready; // @[Decoupled.scala 365:17]
  assign cols_15_15_io_right_out_ready = 1'h1; // @[Stab.scala 102:51]
  assign cols_15_15_io_bottom_out_ready = 1'h1; // @[Stab.scala 94:52]
  assign q_clock = clock;
  assign q_reset = reset;
  assign q_io_enq_valid = cols_0_0_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_io_enq_bits = cols_0_0_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_io_deq_ready = cols_1_0_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_1_clock = clock;
  assign q_1_reset = reset;
  assign q_1_io_enq_valid = cols_1_0_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_1_io_enq_bits = cols_1_0_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_1_io_deq_ready = cols_2_0_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_2_clock = clock;
  assign q_2_reset = reset;
  assign q_2_io_enq_valid = cols_2_0_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_2_io_enq_bits = cols_2_0_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_2_io_deq_ready = cols_3_0_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_3_clock = clock;
  assign q_3_reset = reset;
  assign q_3_io_enq_valid = cols_3_0_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_3_io_enq_bits = cols_3_0_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_3_io_deq_ready = cols_4_0_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_4_clock = clock;
  assign q_4_reset = reset;
  assign q_4_io_enq_valid = cols_4_0_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_4_io_enq_bits = cols_4_0_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_4_io_deq_ready = cols_5_0_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_5_clock = clock;
  assign q_5_reset = reset;
  assign q_5_io_enq_valid = cols_5_0_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_5_io_enq_bits = cols_5_0_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_5_io_deq_ready = cols_6_0_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_6_clock = clock;
  assign q_6_reset = reset;
  assign q_6_io_enq_valid = cols_6_0_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_6_io_enq_bits = cols_6_0_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_6_io_deq_ready = cols_7_0_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_7_clock = clock;
  assign q_7_reset = reset;
  assign q_7_io_enq_valid = cols_7_0_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_7_io_enq_bits = cols_7_0_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_7_io_deq_ready = cols_8_0_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_8_clock = clock;
  assign q_8_reset = reset;
  assign q_8_io_enq_valid = cols_8_0_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_8_io_enq_bits = cols_8_0_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_8_io_deq_ready = cols_9_0_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_9_clock = clock;
  assign q_9_reset = reset;
  assign q_9_io_enq_valid = cols_9_0_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_9_io_enq_bits = cols_9_0_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_9_io_deq_ready = cols_10_0_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_10_clock = clock;
  assign q_10_reset = reset;
  assign q_10_io_enq_valid = cols_10_0_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_10_io_enq_bits = cols_10_0_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_10_io_deq_ready = cols_11_0_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_11_clock = clock;
  assign q_11_reset = reset;
  assign q_11_io_enq_valid = cols_11_0_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_11_io_enq_bits = cols_11_0_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_11_io_deq_ready = cols_12_0_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_12_clock = clock;
  assign q_12_reset = reset;
  assign q_12_io_enq_valid = cols_12_0_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_12_io_enq_bits = cols_12_0_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_12_io_deq_ready = cols_13_0_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_13_clock = clock;
  assign q_13_reset = reset;
  assign q_13_io_enq_valid = cols_13_0_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_13_io_enq_bits = cols_13_0_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_13_io_deq_ready = cols_14_0_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_14_clock = clock;
  assign q_14_reset = reset;
  assign q_14_io_enq_valid = cols_14_0_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_14_io_enq_bits = cols_14_0_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_14_io_deq_ready = cols_15_0_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_15_clock = clock;
  assign q_15_reset = reset;
  assign q_15_io_enq_valid = cols_0_1_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_15_io_enq_bits = cols_0_1_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_15_io_deq_ready = cols_1_1_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_16_clock = clock;
  assign q_16_reset = reset;
  assign q_16_io_enq_valid = cols_1_1_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_16_io_enq_bits = cols_1_1_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_16_io_deq_ready = cols_2_1_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_17_clock = clock;
  assign q_17_reset = reset;
  assign q_17_io_enq_valid = cols_2_1_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_17_io_enq_bits = cols_2_1_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_17_io_deq_ready = cols_3_1_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_18_clock = clock;
  assign q_18_reset = reset;
  assign q_18_io_enq_valid = cols_3_1_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_18_io_enq_bits = cols_3_1_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_18_io_deq_ready = cols_4_1_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_19_clock = clock;
  assign q_19_reset = reset;
  assign q_19_io_enq_valid = cols_4_1_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_19_io_enq_bits = cols_4_1_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_19_io_deq_ready = cols_5_1_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_20_clock = clock;
  assign q_20_reset = reset;
  assign q_20_io_enq_valid = cols_5_1_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_20_io_enq_bits = cols_5_1_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_20_io_deq_ready = cols_6_1_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_21_clock = clock;
  assign q_21_reset = reset;
  assign q_21_io_enq_valid = cols_6_1_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_21_io_enq_bits = cols_6_1_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_21_io_deq_ready = cols_7_1_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_22_clock = clock;
  assign q_22_reset = reset;
  assign q_22_io_enq_valid = cols_7_1_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_22_io_enq_bits = cols_7_1_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_22_io_deq_ready = cols_8_1_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_23_clock = clock;
  assign q_23_reset = reset;
  assign q_23_io_enq_valid = cols_8_1_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_23_io_enq_bits = cols_8_1_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_23_io_deq_ready = cols_9_1_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_24_clock = clock;
  assign q_24_reset = reset;
  assign q_24_io_enq_valid = cols_9_1_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_24_io_enq_bits = cols_9_1_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_24_io_deq_ready = cols_10_1_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_25_clock = clock;
  assign q_25_reset = reset;
  assign q_25_io_enq_valid = cols_10_1_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_25_io_enq_bits = cols_10_1_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_25_io_deq_ready = cols_11_1_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_26_clock = clock;
  assign q_26_reset = reset;
  assign q_26_io_enq_valid = cols_11_1_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_26_io_enq_bits = cols_11_1_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_26_io_deq_ready = cols_12_1_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_27_clock = clock;
  assign q_27_reset = reset;
  assign q_27_io_enq_valid = cols_12_1_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_27_io_enq_bits = cols_12_1_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_27_io_deq_ready = cols_13_1_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_28_clock = clock;
  assign q_28_reset = reset;
  assign q_28_io_enq_valid = cols_13_1_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_28_io_enq_bits = cols_13_1_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_28_io_deq_ready = cols_14_1_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_29_clock = clock;
  assign q_29_reset = reset;
  assign q_29_io_enq_valid = cols_14_1_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_29_io_enq_bits = cols_14_1_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_29_io_deq_ready = cols_15_1_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_30_clock = clock;
  assign q_30_reset = reset;
  assign q_30_io_enq_valid = cols_0_2_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_30_io_enq_bits = cols_0_2_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_30_io_deq_ready = cols_1_2_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_31_clock = clock;
  assign q_31_reset = reset;
  assign q_31_io_enq_valid = cols_1_2_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_31_io_enq_bits = cols_1_2_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_31_io_deq_ready = cols_2_2_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_32_clock = clock;
  assign q_32_reset = reset;
  assign q_32_io_enq_valid = cols_2_2_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_32_io_enq_bits = cols_2_2_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_32_io_deq_ready = cols_3_2_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_33_clock = clock;
  assign q_33_reset = reset;
  assign q_33_io_enq_valid = cols_3_2_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_33_io_enq_bits = cols_3_2_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_33_io_deq_ready = cols_4_2_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_34_clock = clock;
  assign q_34_reset = reset;
  assign q_34_io_enq_valid = cols_4_2_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_34_io_enq_bits = cols_4_2_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_34_io_deq_ready = cols_5_2_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_35_clock = clock;
  assign q_35_reset = reset;
  assign q_35_io_enq_valid = cols_5_2_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_35_io_enq_bits = cols_5_2_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_35_io_deq_ready = cols_6_2_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_36_clock = clock;
  assign q_36_reset = reset;
  assign q_36_io_enq_valid = cols_6_2_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_36_io_enq_bits = cols_6_2_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_36_io_deq_ready = cols_7_2_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_37_clock = clock;
  assign q_37_reset = reset;
  assign q_37_io_enq_valid = cols_7_2_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_37_io_enq_bits = cols_7_2_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_37_io_deq_ready = cols_8_2_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_38_clock = clock;
  assign q_38_reset = reset;
  assign q_38_io_enq_valid = cols_8_2_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_38_io_enq_bits = cols_8_2_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_38_io_deq_ready = cols_9_2_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_39_clock = clock;
  assign q_39_reset = reset;
  assign q_39_io_enq_valid = cols_9_2_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_39_io_enq_bits = cols_9_2_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_39_io_deq_ready = cols_10_2_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_40_clock = clock;
  assign q_40_reset = reset;
  assign q_40_io_enq_valid = cols_10_2_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_40_io_enq_bits = cols_10_2_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_40_io_deq_ready = cols_11_2_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_41_clock = clock;
  assign q_41_reset = reset;
  assign q_41_io_enq_valid = cols_11_2_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_41_io_enq_bits = cols_11_2_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_41_io_deq_ready = cols_12_2_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_42_clock = clock;
  assign q_42_reset = reset;
  assign q_42_io_enq_valid = cols_12_2_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_42_io_enq_bits = cols_12_2_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_42_io_deq_ready = cols_13_2_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_43_clock = clock;
  assign q_43_reset = reset;
  assign q_43_io_enq_valid = cols_13_2_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_43_io_enq_bits = cols_13_2_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_43_io_deq_ready = cols_14_2_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_44_clock = clock;
  assign q_44_reset = reset;
  assign q_44_io_enq_valid = cols_14_2_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_44_io_enq_bits = cols_14_2_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_44_io_deq_ready = cols_15_2_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_45_clock = clock;
  assign q_45_reset = reset;
  assign q_45_io_enq_valid = cols_0_3_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_45_io_enq_bits = cols_0_3_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_45_io_deq_ready = cols_1_3_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_46_clock = clock;
  assign q_46_reset = reset;
  assign q_46_io_enq_valid = cols_1_3_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_46_io_enq_bits = cols_1_3_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_46_io_deq_ready = cols_2_3_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_47_clock = clock;
  assign q_47_reset = reset;
  assign q_47_io_enq_valid = cols_2_3_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_47_io_enq_bits = cols_2_3_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_47_io_deq_ready = cols_3_3_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_48_clock = clock;
  assign q_48_reset = reset;
  assign q_48_io_enq_valid = cols_3_3_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_48_io_enq_bits = cols_3_3_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_48_io_deq_ready = cols_4_3_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_49_clock = clock;
  assign q_49_reset = reset;
  assign q_49_io_enq_valid = cols_4_3_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_49_io_enq_bits = cols_4_3_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_49_io_deq_ready = cols_5_3_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_50_clock = clock;
  assign q_50_reset = reset;
  assign q_50_io_enq_valid = cols_5_3_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_50_io_enq_bits = cols_5_3_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_50_io_deq_ready = cols_6_3_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_51_clock = clock;
  assign q_51_reset = reset;
  assign q_51_io_enq_valid = cols_6_3_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_51_io_enq_bits = cols_6_3_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_51_io_deq_ready = cols_7_3_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_52_clock = clock;
  assign q_52_reset = reset;
  assign q_52_io_enq_valid = cols_7_3_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_52_io_enq_bits = cols_7_3_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_52_io_deq_ready = cols_8_3_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_53_clock = clock;
  assign q_53_reset = reset;
  assign q_53_io_enq_valid = cols_8_3_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_53_io_enq_bits = cols_8_3_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_53_io_deq_ready = cols_9_3_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_54_clock = clock;
  assign q_54_reset = reset;
  assign q_54_io_enq_valid = cols_9_3_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_54_io_enq_bits = cols_9_3_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_54_io_deq_ready = cols_10_3_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_55_clock = clock;
  assign q_55_reset = reset;
  assign q_55_io_enq_valid = cols_10_3_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_55_io_enq_bits = cols_10_3_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_55_io_deq_ready = cols_11_3_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_56_clock = clock;
  assign q_56_reset = reset;
  assign q_56_io_enq_valid = cols_11_3_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_56_io_enq_bits = cols_11_3_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_56_io_deq_ready = cols_12_3_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_57_clock = clock;
  assign q_57_reset = reset;
  assign q_57_io_enq_valid = cols_12_3_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_57_io_enq_bits = cols_12_3_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_57_io_deq_ready = cols_13_3_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_58_clock = clock;
  assign q_58_reset = reset;
  assign q_58_io_enq_valid = cols_13_3_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_58_io_enq_bits = cols_13_3_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_58_io_deq_ready = cols_14_3_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_59_clock = clock;
  assign q_59_reset = reset;
  assign q_59_io_enq_valid = cols_14_3_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_59_io_enq_bits = cols_14_3_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_59_io_deq_ready = cols_15_3_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_60_clock = clock;
  assign q_60_reset = reset;
  assign q_60_io_enq_valid = cols_0_4_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_60_io_enq_bits = cols_0_4_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_60_io_deq_ready = cols_1_4_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_61_clock = clock;
  assign q_61_reset = reset;
  assign q_61_io_enq_valid = cols_1_4_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_61_io_enq_bits = cols_1_4_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_61_io_deq_ready = cols_2_4_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_62_clock = clock;
  assign q_62_reset = reset;
  assign q_62_io_enq_valid = cols_2_4_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_62_io_enq_bits = cols_2_4_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_62_io_deq_ready = cols_3_4_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_63_clock = clock;
  assign q_63_reset = reset;
  assign q_63_io_enq_valid = cols_3_4_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_63_io_enq_bits = cols_3_4_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_63_io_deq_ready = cols_4_4_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_64_clock = clock;
  assign q_64_reset = reset;
  assign q_64_io_enq_valid = cols_4_4_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_64_io_enq_bits = cols_4_4_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_64_io_deq_ready = cols_5_4_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_65_clock = clock;
  assign q_65_reset = reset;
  assign q_65_io_enq_valid = cols_5_4_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_65_io_enq_bits = cols_5_4_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_65_io_deq_ready = cols_6_4_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_66_clock = clock;
  assign q_66_reset = reset;
  assign q_66_io_enq_valid = cols_6_4_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_66_io_enq_bits = cols_6_4_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_66_io_deq_ready = cols_7_4_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_67_clock = clock;
  assign q_67_reset = reset;
  assign q_67_io_enq_valid = cols_7_4_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_67_io_enq_bits = cols_7_4_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_67_io_deq_ready = cols_8_4_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_68_clock = clock;
  assign q_68_reset = reset;
  assign q_68_io_enq_valid = cols_8_4_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_68_io_enq_bits = cols_8_4_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_68_io_deq_ready = cols_9_4_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_69_clock = clock;
  assign q_69_reset = reset;
  assign q_69_io_enq_valid = cols_9_4_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_69_io_enq_bits = cols_9_4_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_69_io_deq_ready = cols_10_4_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_70_clock = clock;
  assign q_70_reset = reset;
  assign q_70_io_enq_valid = cols_10_4_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_70_io_enq_bits = cols_10_4_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_70_io_deq_ready = cols_11_4_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_71_clock = clock;
  assign q_71_reset = reset;
  assign q_71_io_enq_valid = cols_11_4_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_71_io_enq_bits = cols_11_4_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_71_io_deq_ready = cols_12_4_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_72_clock = clock;
  assign q_72_reset = reset;
  assign q_72_io_enq_valid = cols_12_4_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_72_io_enq_bits = cols_12_4_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_72_io_deq_ready = cols_13_4_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_73_clock = clock;
  assign q_73_reset = reset;
  assign q_73_io_enq_valid = cols_13_4_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_73_io_enq_bits = cols_13_4_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_73_io_deq_ready = cols_14_4_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_74_clock = clock;
  assign q_74_reset = reset;
  assign q_74_io_enq_valid = cols_14_4_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_74_io_enq_bits = cols_14_4_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_74_io_deq_ready = cols_15_4_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_75_clock = clock;
  assign q_75_reset = reset;
  assign q_75_io_enq_valid = cols_0_5_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_75_io_enq_bits = cols_0_5_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_75_io_deq_ready = cols_1_5_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_76_clock = clock;
  assign q_76_reset = reset;
  assign q_76_io_enq_valid = cols_1_5_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_76_io_enq_bits = cols_1_5_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_76_io_deq_ready = cols_2_5_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_77_clock = clock;
  assign q_77_reset = reset;
  assign q_77_io_enq_valid = cols_2_5_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_77_io_enq_bits = cols_2_5_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_77_io_deq_ready = cols_3_5_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_78_clock = clock;
  assign q_78_reset = reset;
  assign q_78_io_enq_valid = cols_3_5_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_78_io_enq_bits = cols_3_5_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_78_io_deq_ready = cols_4_5_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_79_clock = clock;
  assign q_79_reset = reset;
  assign q_79_io_enq_valid = cols_4_5_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_79_io_enq_bits = cols_4_5_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_79_io_deq_ready = cols_5_5_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_80_clock = clock;
  assign q_80_reset = reset;
  assign q_80_io_enq_valid = cols_5_5_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_80_io_enq_bits = cols_5_5_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_80_io_deq_ready = cols_6_5_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_81_clock = clock;
  assign q_81_reset = reset;
  assign q_81_io_enq_valid = cols_6_5_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_81_io_enq_bits = cols_6_5_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_81_io_deq_ready = cols_7_5_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_82_clock = clock;
  assign q_82_reset = reset;
  assign q_82_io_enq_valid = cols_7_5_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_82_io_enq_bits = cols_7_5_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_82_io_deq_ready = cols_8_5_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_83_clock = clock;
  assign q_83_reset = reset;
  assign q_83_io_enq_valid = cols_8_5_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_83_io_enq_bits = cols_8_5_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_83_io_deq_ready = cols_9_5_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_84_clock = clock;
  assign q_84_reset = reset;
  assign q_84_io_enq_valid = cols_9_5_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_84_io_enq_bits = cols_9_5_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_84_io_deq_ready = cols_10_5_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_85_clock = clock;
  assign q_85_reset = reset;
  assign q_85_io_enq_valid = cols_10_5_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_85_io_enq_bits = cols_10_5_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_85_io_deq_ready = cols_11_5_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_86_clock = clock;
  assign q_86_reset = reset;
  assign q_86_io_enq_valid = cols_11_5_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_86_io_enq_bits = cols_11_5_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_86_io_deq_ready = cols_12_5_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_87_clock = clock;
  assign q_87_reset = reset;
  assign q_87_io_enq_valid = cols_12_5_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_87_io_enq_bits = cols_12_5_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_87_io_deq_ready = cols_13_5_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_88_clock = clock;
  assign q_88_reset = reset;
  assign q_88_io_enq_valid = cols_13_5_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_88_io_enq_bits = cols_13_5_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_88_io_deq_ready = cols_14_5_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_89_clock = clock;
  assign q_89_reset = reset;
  assign q_89_io_enq_valid = cols_14_5_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_89_io_enq_bits = cols_14_5_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_89_io_deq_ready = cols_15_5_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_90_clock = clock;
  assign q_90_reset = reset;
  assign q_90_io_enq_valid = cols_0_6_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_90_io_enq_bits = cols_0_6_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_90_io_deq_ready = cols_1_6_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_91_clock = clock;
  assign q_91_reset = reset;
  assign q_91_io_enq_valid = cols_1_6_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_91_io_enq_bits = cols_1_6_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_91_io_deq_ready = cols_2_6_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_92_clock = clock;
  assign q_92_reset = reset;
  assign q_92_io_enq_valid = cols_2_6_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_92_io_enq_bits = cols_2_6_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_92_io_deq_ready = cols_3_6_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_93_clock = clock;
  assign q_93_reset = reset;
  assign q_93_io_enq_valid = cols_3_6_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_93_io_enq_bits = cols_3_6_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_93_io_deq_ready = cols_4_6_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_94_clock = clock;
  assign q_94_reset = reset;
  assign q_94_io_enq_valid = cols_4_6_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_94_io_enq_bits = cols_4_6_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_94_io_deq_ready = cols_5_6_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_95_clock = clock;
  assign q_95_reset = reset;
  assign q_95_io_enq_valid = cols_5_6_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_95_io_enq_bits = cols_5_6_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_95_io_deq_ready = cols_6_6_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_96_clock = clock;
  assign q_96_reset = reset;
  assign q_96_io_enq_valid = cols_6_6_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_96_io_enq_bits = cols_6_6_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_96_io_deq_ready = cols_7_6_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_97_clock = clock;
  assign q_97_reset = reset;
  assign q_97_io_enq_valid = cols_7_6_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_97_io_enq_bits = cols_7_6_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_97_io_deq_ready = cols_8_6_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_98_clock = clock;
  assign q_98_reset = reset;
  assign q_98_io_enq_valid = cols_8_6_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_98_io_enq_bits = cols_8_6_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_98_io_deq_ready = cols_9_6_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_99_clock = clock;
  assign q_99_reset = reset;
  assign q_99_io_enq_valid = cols_9_6_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_99_io_enq_bits = cols_9_6_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_99_io_deq_ready = cols_10_6_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_100_clock = clock;
  assign q_100_reset = reset;
  assign q_100_io_enq_valid = cols_10_6_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_100_io_enq_bits = cols_10_6_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_100_io_deq_ready = cols_11_6_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_101_clock = clock;
  assign q_101_reset = reset;
  assign q_101_io_enq_valid = cols_11_6_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_101_io_enq_bits = cols_11_6_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_101_io_deq_ready = cols_12_6_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_102_clock = clock;
  assign q_102_reset = reset;
  assign q_102_io_enq_valid = cols_12_6_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_102_io_enq_bits = cols_12_6_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_102_io_deq_ready = cols_13_6_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_103_clock = clock;
  assign q_103_reset = reset;
  assign q_103_io_enq_valid = cols_13_6_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_103_io_enq_bits = cols_13_6_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_103_io_deq_ready = cols_14_6_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_104_clock = clock;
  assign q_104_reset = reset;
  assign q_104_io_enq_valid = cols_14_6_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_104_io_enq_bits = cols_14_6_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_104_io_deq_ready = cols_15_6_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_105_clock = clock;
  assign q_105_reset = reset;
  assign q_105_io_enq_valid = cols_0_7_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_105_io_enq_bits = cols_0_7_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_105_io_deq_ready = cols_1_7_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_106_clock = clock;
  assign q_106_reset = reset;
  assign q_106_io_enq_valid = cols_1_7_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_106_io_enq_bits = cols_1_7_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_106_io_deq_ready = cols_2_7_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_107_clock = clock;
  assign q_107_reset = reset;
  assign q_107_io_enq_valid = cols_2_7_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_107_io_enq_bits = cols_2_7_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_107_io_deq_ready = cols_3_7_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_108_clock = clock;
  assign q_108_reset = reset;
  assign q_108_io_enq_valid = cols_3_7_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_108_io_enq_bits = cols_3_7_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_108_io_deq_ready = cols_4_7_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_109_clock = clock;
  assign q_109_reset = reset;
  assign q_109_io_enq_valid = cols_4_7_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_109_io_enq_bits = cols_4_7_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_109_io_deq_ready = cols_5_7_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_110_clock = clock;
  assign q_110_reset = reset;
  assign q_110_io_enq_valid = cols_5_7_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_110_io_enq_bits = cols_5_7_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_110_io_deq_ready = cols_6_7_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_111_clock = clock;
  assign q_111_reset = reset;
  assign q_111_io_enq_valid = cols_6_7_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_111_io_enq_bits = cols_6_7_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_111_io_deq_ready = cols_7_7_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_112_clock = clock;
  assign q_112_reset = reset;
  assign q_112_io_enq_valid = cols_7_7_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_112_io_enq_bits = cols_7_7_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_112_io_deq_ready = cols_8_7_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_113_clock = clock;
  assign q_113_reset = reset;
  assign q_113_io_enq_valid = cols_8_7_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_113_io_enq_bits = cols_8_7_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_113_io_deq_ready = cols_9_7_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_114_clock = clock;
  assign q_114_reset = reset;
  assign q_114_io_enq_valid = cols_9_7_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_114_io_enq_bits = cols_9_7_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_114_io_deq_ready = cols_10_7_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_115_clock = clock;
  assign q_115_reset = reset;
  assign q_115_io_enq_valid = cols_10_7_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_115_io_enq_bits = cols_10_7_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_115_io_deq_ready = cols_11_7_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_116_clock = clock;
  assign q_116_reset = reset;
  assign q_116_io_enq_valid = cols_11_7_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_116_io_enq_bits = cols_11_7_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_116_io_deq_ready = cols_12_7_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_117_clock = clock;
  assign q_117_reset = reset;
  assign q_117_io_enq_valid = cols_12_7_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_117_io_enq_bits = cols_12_7_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_117_io_deq_ready = cols_13_7_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_118_clock = clock;
  assign q_118_reset = reset;
  assign q_118_io_enq_valid = cols_13_7_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_118_io_enq_bits = cols_13_7_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_118_io_deq_ready = cols_14_7_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_119_clock = clock;
  assign q_119_reset = reset;
  assign q_119_io_enq_valid = cols_14_7_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_119_io_enq_bits = cols_14_7_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_119_io_deq_ready = cols_15_7_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_120_clock = clock;
  assign q_120_reset = reset;
  assign q_120_io_enq_valid = cols_0_8_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_120_io_enq_bits = cols_0_8_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_120_io_deq_ready = cols_1_8_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_121_clock = clock;
  assign q_121_reset = reset;
  assign q_121_io_enq_valid = cols_1_8_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_121_io_enq_bits = cols_1_8_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_121_io_deq_ready = cols_2_8_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_122_clock = clock;
  assign q_122_reset = reset;
  assign q_122_io_enq_valid = cols_2_8_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_122_io_enq_bits = cols_2_8_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_122_io_deq_ready = cols_3_8_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_123_clock = clock;
  assign q_123_reset = reset;
  assign q_123_io_enq_valid = cols_3_8_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_123_io_enq_bits = cols_3_8_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_123_io_deq_ready = cols_4_8_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_124_clock = clock;
  assign q_124_reset = reset;
  assign q_124_io_enq_valid = cols_4_8_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_124_io_enq_bits = cols_4_8_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_124_io_deq_ready = cols_5_8_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_125_clock = clock;
  assign q_125_reset = reset;
  assign q_125_io_enq_valid = cols_5_8_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_125_io_enq_bits = cols_5_8_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_125_io_deq_ready = cols_6_8_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_126_clock = clock;
  assign q_126_reset = reset;
  assign q_126_io_enq_valid = cols_6_8_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_126_io_enq_bits = cols_6_8_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_126_io_deq_ready = cols_7_8_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_127_clock = clock;
  assign q_127_reset = reset;
  assign q_127_io_enq_valid = cols_7_8_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_127_io_enq_bits = cols_7_8_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_127_io_deq_ready = cols_8_8_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_128_clock = clock;
  assign q_128_reset = reset;
  assign q_128_io_enq_valid = cols_8_8_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_128_io_enq_bits = cols_8_8_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_128_io_deq_ready = cols_9_8_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_129_clock = clock;
  assign q_129_reset = reset;
  assign q_129_io_enq_valid = cols_9_8_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_129_io_enq_bits = cols_9_8_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_129_io_deq_ready = cols_10_8_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_130_clock = clock;
  assign q_130_reset = reset;
  assign q_130_io_enq_valid = cols_10_8_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_130_io_enq_bits = cols_10_8_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_130_io_deq_ready = cols_11_8_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_131_clock = clock;
  assign q_131_reset = reset;
  assign q_131_io_enq_valid = cols_11_8_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_131_io_enq_bits = cols_11_8_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_131_io_deq_ready = cols_12_8_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_132_clock = clock;
  assign q_132_reset = reset;
  assign q_132_io_enq_valid = cols_12_8_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_132_io_enq_bits = cols_12_8_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_132_io_deq_ready = cols_13_8_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_133_clock = clock;
  assign q_133_reset = reset;
  assign q_133_io_enq_valid = cols_13_8_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_133_io_enq_bits = cols_13_8_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_133_io_deq_ready = cols_14_8_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_134_clock = clock;
  assign q_134_reset = reset;
  assign q_134_io_enq_valid = cols_14_8_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_134_io_enq_bits = cols_14_8_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_134_io_deq_ready = cols_15_8_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_135_clock = clock;
  assign q_135_reset = reset;
  assign q_135_io_enq_valid = cols_0_9_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_135_io_enq_bits = cols_0_9_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_135_io_deq_ready = cols_1_9_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_136_clock = clock;
  assign q_136_reset = reset;
  assign q_136_io_enq_valid = cols_1_9_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_136_io_enq_bits = cols_1_9_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_136_io_deq_ready = cols_2_9_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_137_clock = clock;
  assign q_137_reset = reset;
  assign q_137_io_enq_valid = cols_2_9_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_137_io_enq_bits = cols_2_9_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_137_io_deq_ready = cols_3_9_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_138_clock = clock;
  assign q_138_reset = reset;
  assign q_138_io_enq_valid = cols_3_9_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_138_io_enq_bits = cols_3_9_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_138_io_deq_ready = cols_4_9_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_139_clock = clock;
  assign q_139_reset = reset;
  assign q_139_io_enq_valid = cols_4_9_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_139_io_enq_bits = cols_4_9_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_139_io_deq_ready = cols_5_9_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_140_clock = clock;
  assign q_140_reset = reset;
  assign q_140_io_enq_valid = cols_5_9_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_140_io_enq_bits = cols_5_9_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_140_io_deq_ready = cols_6_9_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_141_clock = clock;
  assign q_141_reset = reset;
  assign q_141_io_enq_valid = cols_6_9_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_141_io_enq_bits = cols_6_9_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_141_io_deq_ready = cols_7_9_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_142_clock = clock;
  assign q_142_reset = reset;
  assign q_142_io_enq_valid = cols_7_9_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_142_io_enq_bits = cols_7_9_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_142_io_deq_ready = cols_8_9_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_143_clock = clock;
  assign q_143_reset = reset;
  assign q_143_io_enq_valid = cols_8_9_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_143_io_enq_bits = cols_8_9_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_143_io_deq_ready = cols_9_9_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_144_clock = clock;
  assign q_144_reset = reset;
  assign q_144_io_enq_valid = cols_9_9_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_144_io_enq_bits = cols_9_9_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_144_io_deq_ready = cols_10_9_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_145_clock = clock;
  assign q_145_reset = reset;
  assign q_145_io_enq_valid = cols_10_9_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_145_io_enq_bits = cols_10_9_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_145_io_deq_ready = cols_11_9_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_146_clock = clock;
  assign q_146_reset = reset;
  assign q_146_io_enq_valid = cols_11_9_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_146_io_enq_bits = cols_11_9_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_146_io_deq_ready = cols_12_9_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_147_clock = clock;
  assign q_147_reset = reset;
  assign q_147_io_enq_valid = cols_12_9_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_147_io_enq_bits = cols_12_9_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_147_io_deq_ready = cols_13_9_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_148_clock = clock;
  assign q_148_reset = reset;
  assign q_148_io_enq_valid = cols_13_9_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_148_io_enq_bits = cols_13_9_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_148_io_deq_ready = cols_14_9_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_149_clock = clock;
  assign q_149_reset = reset;
  assign q_149_io_enq_valid = cols_14_9_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_149_io_enq_bits = cols_14_9_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_149_io_deq_ready = cols_15_9_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_150_clock = clock;
  assign q_150_reset = reset;
  assign q_150_io_enq_valid = cols_0_10_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_150_io_enq_bits = cols_0_10_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_150_io_deq_ready = cols_1_10_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_151_clock = clock;
  assign q_151_reset = reset;
  assign q_151_io_enq_valid = cols_1_10_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_151_io_enq_bits = cols_1_10_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_151_io_deq_ready = cols_2_10_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_152_clock = clock;
  assign q_152_reset = reset;
  assign q_152_io_enq_valid = cols_2_10_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_152_io_enq_bits = cols_2_10_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_152_io_deq_ready = cols_3_10_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_153_clock = clock;
  assign q_153_reset = reset;
  assign q_153_io_enq_valid = cols_3_10_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_153_io_enq_bits = cols_3_10_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_153_io_deq_ready = cols_4_10_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_154_clock = clock;
  assign q_154_reset = reset;
  assign q_154_io_enq_valid = cols_4_10_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_154_io_enq_bits = cols_4_10_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_154_io_deq_ready = cols_5_10_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_155_clock = clock;
  assign q_155_reset = reset;
  assign q_155_io_enq_valid = cols_5_10_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_155_io_enq_bits = cols_5_10_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_155_io_deq_ready = cols_6_10_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_156_clock = clock;
  assign q_156_reset = reset;
  assign q_156_io_enq_valid = cols_6_10_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_156_io_enq_bits = cols_6_10_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_156_io_deq_ready = cols_7_10_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_157_clock = clock;
  assign q_157_reset = reset;
  assign q_157_io_enq_valid = cols_7_10_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_157_io_enq_bits = cols_7_10_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_157_io_deq_ready = cols_8_10_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_158_clock = clock;
  assign q_158_reset = reset;
  assign q_158_io_enq_valid = cols_8_10_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_158_io_enq_bits = cols_8_10_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_158_io_deq_ready = cols_9_10_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_159_clock = clock;
  assign q_159_reset = reset;
  assign q_159_io_enq_valid = cols_9_10_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_159_io_enq_bits = cols_9_10_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_159_io_deq_ready = cols_10_10_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_160_clock = clock;
  assign q_160_reset = reset;
  assign q_160_io_enq_valid = cols_10_10_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_160_io_enq_bits = cols_10_10_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_160_io_deq_ready = cols_11_10_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_161_clock = clock;
  assign q_161_reset = reset;
  assign q_161_io_enq_valid = cols_11_10_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_161_io_enq_bits = cols_11_10_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_161_io_deq_ready = cols_12_10_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_162_clock = clock;
  assign q_162_reset = reset;
  assign q_162_io_enq_valid = cols_12_10_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_162_io_enq_bits = cols_12_10_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_162_io_deq_ready = cols_13_10_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_163_clock = clock;
  assign q_163_reset = reset;
  assign q_163_io_enq_valid = cols_13_10_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_163_io_enq_bits = cols_13_10_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_163_io_deq_ready = cols_14_10_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_164_clock = clock;
  assign q_164_reset = reset;
  assign q_164_io_enq_valid = cols_14_10_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_164_io_enq_bits = cols_14_10_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_164_io_deq_ready = cols_15_10_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_165_clock = clock;
  assign q_165_reset = reset;
  assign q_165_io_enq_valid = cols_0_11_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_165_io_enq_bits = cols_0_11_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_165_io_deq_ready = cols_1_11_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_166_clock = clock;
  assign q_166_reset = reset;
  assign q_166_io_enq_valid = cols_1_11_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_166_io_enq_bits = cols_1_11_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_166_io_deq_ready = cols_2_11_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_167_clock = clock;
  assign q_167_reset = reset;
  assign q_167_io_enq_valid = cols_2_11_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_167_io_enq_bits = cols_2_11_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_167_io_deq_ready = cols_3_11_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_168_clock = clock;
  assign q_168_reset = reset;
  assign q_168_io_enq_valid = cols_3_11_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_168_io_enq_bits = cols_3_11_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_168_io_deq_ready = cols_4_11_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_169_clock = clock;
  assign q_169_reset = reset;
  assign q_169_io_enq_valid = cols_4_11_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_169_io_enq_bits = cols_4_11_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_169_io_deq_ready = cols_5_11_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_170_clock = clock;
  assign q_170_reset = reset;
  assign q_170_io_enq_valid = cols_5_11_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_170_io_enq_bits = cols_5_11_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_170_io_deq_ready = cols_6_11_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_171_clock = clock;
  assign q_171_reset = reset;
  assign q_171_io_enq_valid = cols_6_11_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_171_io_enq_bits = cols_6_11_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_171_io_deq_ready = cols_7_11_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_172_clock = clock;
  assign q_172_reset = reset;
  assign q_172_io_enq_valid = cols_7_11_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_172_io_enq_bits = cols_7_11_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_172_io_deq_ready = cols_8_11_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_173_clock = clock;
  assign q_173_reset = reset;
  assign q_173_io_enq_valid = cols_8_11_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_173_io_enq_bits = cols_8_11_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_173_io_deq_ready = cols_9_11_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_174_clock = clock;
  assign q_174_reset = reset;
  assign q_174_io_enq_valid = cols_9_11_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_174_io_enq_bits = cols_9_11_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_174_io_deq_ready = cols_10_11_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_175_clock = clock;
  assign q_175_reset = reset;
  assign q_175_io_enq_valid = cols_10_11_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_175_io_enq_bits = cols_10_11_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_175_io_deq_ready = cols_11_11_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_176_clock = clock;
  assign q_176_reset = reset;
  assign q_176_io_enq_valid = cols_11_11_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_176_io_enq_bits = cols_11_11_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_176_io_deq_ready = cols_12_11_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_177_clock = clock;
  assign q_177_reset = reset;
  assign q_177_io_enq_valid = cols_12_11_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_177_io_enq_bits = cols_12_11_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_177_io_deq_ready = cols_13_11_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_178_clock = clock;
  assign q_178_reset = reset;
  assign q_178_io_enq_valid = cols_13_11_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_178_io_enq_bits = cols_13_11_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_178_io_deq_ready = cols_14_11_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_179_clock = clock;
  assign q_179_reset = reset;
  assign q_179_io_enq_valid = cols_14_11_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_179_io_enq_bits = cols_14_11_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_179_io_deq_ready = cols_15_11_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_180_clock = clock;
  assign q_180_reset = reset;
  assign q_180_io_enq_valid = cols_0_12_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_180_io_enq_bits = cols_0_12_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_180_io_deq_ready = cols_1_12_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_181_clock = clock;
  assign q_181_reset = reset;
  assign q_181_io_enq_valid = cols_1_12_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_181_io_enq_bits = cols_1_12_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_181_io_deq_ready = cols_2_12_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_182_clock = clock;
  assign q_182_reset = reset;
  assign q_182_io_enq_valid = cols_2_12_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_182_io_enq_bits = cols_2_12_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_182_io_deq_ready = cols_3_12_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_183_clock = clock;
  assign q_183_reset = reset;
  assign q_183_io_enq_valid = cols_3_12_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_183_io_enq_bits = cols_3_12_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_183_io_deq_ready = cols_4_12_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_184_clock = clock;
  assign q_184_reset = reset;
  assign q_184_io_enq_valid = cols_4_12_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_184_io_enq_bits = cols_4_12_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_184_io_deq_ready = cols_5_12_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_185_clock = clock;
  assign q_185_reset = reset;
  assign q_185_io_enq_valid = cols_5_12_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_185_io_enq_bits = cols_5_12_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_185_io_deq_ready = cols_6_12_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_186_clock = clock;
  assign q_186_reset = reset;
  assign q_186_io_enq_valid = cols_6_12_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_186_io_enq_bits = cols_6_12_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_186_io_deq_ready = cols_7_12_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_187_clock = clock;
  assign q_187_reset = reset;
  assign q_187_io_enq_valid = cols_7_12_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_187_io_enq_bits = cols_7_12_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_187_io_deq_ready = cols_8_12_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_188_clock = clock;
  assign q_188_reset = reset;
  assign q_188_io_enq_valid = cols_8_12_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_188_io_enq_bits = cols_8_12_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_188_io_deq_ready = cols_9_12_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_189_clock = clock;
  assign q_189_reset = reset;
  assign q_189_io_enq_valid = cols_9_12_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_189_io_enq_bits = cols_9_12_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_189_io_deq_ready = cols_10_12_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_190_clock = clock;
  assign q_190_reset = reset;
  assign q_190_io_enq_valid = cols_10_12_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_190_io_enq_bits = cols_10_12_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_190_io_deq_ready = cols_11_12_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_191_clock = clock;
  assign q_191_reset = reset;
  assign q_191_io_enq_valid = cols_11_12_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_191_io_enq_bits = cols_11_12_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_191_io_deq_ready = cols_12_12_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_192_clock = clock;
  assign q_192_reset = reset;
  assign q_192_io_enq_valid = cols_12_12_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_192_io_enq_bits = cols_12_12_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_192_io_deq_ready = cols_13_12_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_193_clock = clock;
  assign q_193_reset = reset;
  assign q_193_io_enq_valid = cols_13_12_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_193_io_enq_bits = cols_13_12_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_193_io_deq_ready = cols_14_12_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_194_clock = clock;
  assign q_194_reset = reset;
  assign q_194_io_enq_valid = cols_14_12_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_194_io_enq_bits = cols_14_12_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_194_io_deq_ready = cols_15_12_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_195_clock = clock;
  assign q_195_reset = reset;
  assign q_195_io_enq_valid = cols_0_13_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_195_io_enq_bits = cols_0_13_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_195_io_deq_ready = cols_1_13_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_196_clock = clock;
  assign q_196_reset = reset;
  assign q_196_io_enq_valid = cols_1_13_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_196_io_enq_bits = cols_1_13_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_196_io_deq_ready = cols_2_13_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_197_clock = clock;
  assign q_197_reset = reset;
  assign q_197_io_enq_valid = cols_2_13_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_197_io_enq_bits = cols_2_13_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_197_io_deq_ready = cols_3_13_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_198_clock = clock;
  assign q_198_reset = reset;
  assign q_198_io_enq_valid = cols_3_13_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_198_io_enq_bits = cols_3_13_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_198_io_deq_ready = cols_4_13_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_199_clock = clock;
  assign q_199_reset = reset;
  assign q_199_io_enq_valid = cols_4_13_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_199_io_enq_bits = cols_4_13_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_199_io_deq_ready = cols_5_13_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_200_clock = clock;
  assign q_200_reset = reset;
  assign q_200_io_enq_valid = cols_5_13_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_200_io_enq_bits = cols_5_13_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_200_io_deq_ready = cols_6_13_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_201_clock = clock;
  assign q_201_reset = reset;
  assign q_201_io_enq_valid = cols_6_13_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_201_io_enq_bits = cols_6_13_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_201_io_deq_ready = cols_7_13_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_202_clock = clock;
  assign q_202_reset = reset;
  assign q_202_io_enq_valid = cols_7_13_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_202_io_enq_bits = cols_7_13_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_202_io_deq_ready = cols_8_13_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_203_clock = clock;
  assign q_203_reset = reset;
  assign q_203_io_enq_valid = cols_8_13_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_203_io_enq_bits = cols_8_13_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_203_io_deq_ready = cols_9_13_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_204_clock = clock;
  assign q_204_reset = reset;
  assign q_204_io_enq_valid = cols_9_13_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_204_io_enq_bits = cols_9_13_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_204_io_deq_ready = cols_10_13_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_205_clock = clock;
  assign q_205_reset = reset;
  assign q_205_io_enq_valid = cols_10_13_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_205_io_enq_bits = cols_10_13_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_205_io_deq_ready = cols_11_13_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_206_clock = clock;
  assign q_206_reset = reset;
  assign q_206_io_enq_valid = cols_11_13_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_206_io_enq_bits = cols_11_13_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_206_io_deq_ready = cols_12_13_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_207_clock = clock;
  assign q_207_reset = reset;
  assign q_207_io_enq_valid = cols_12_13_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_207_io_enq_bits = cols_12_13_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_207_io_deq_ready = cols_13_13_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_208_clock = clock;
  assign q_208_reset = reset;
  assign q_208_io_enq_valid = cols_13_13_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_208_io_enq_bits = cols_13_13_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_208_io_deq_ready = cols_14_13_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_209_clock = clock;
  assign q_209_reset = reset;
  assign q_209_io_enq_valid = cols_14_13_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_209_io_enq_bits = cols_14_13_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_209_io_deq_ready = cols_15_13_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_210_clock = clock;
  assign q_210_reset = reset;
  assign q_210_io_enq_valid = cols_0_14_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_210_io_enq_bits = cols_0_14_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_210_io_deq_ready = cols_1_14_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_211_clock = clock;
  assign q_211_reset = reset;
  assign q_211_io_enq_valid = cols_1_14_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_211_io_enq_bits = cols_1_14_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_211_io_deq_ready = cols_2_14_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_212_clock = clock;
  assign q_212_reset = reset;
  assign q_212_io_enq_valid = cols_2_14_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_212_io_enq_bits = cols_2_14_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_212_io_deq_ready = cols_3_14_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_213_clock = clock;
  assign q_213_reset = reset;
  assign q_213_io_enq_valid = cols_3_14_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_213_io_enq_bits = cols_3_14_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_213_io_deq_ready = cols_4_14_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_214_clock = clock;
  assign q_214_reset = reset;
  assign q_214_io_enq_valid = cols_4_14_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_214_io_enq_bits = cols_4_14_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_214_io_deq_ready = cols_5_14_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_215_clock = clock;
  assign q_215_reset = reset;
  assign q_215_io_enq_valid = cols_5_14_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_215_io_enq_bits = cols_5_14_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_215_io_deq_ready = cols_6_14_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_216_clock = clock;
  assign q_216_reset = reset;
  assign q_216_io_enq_valid = cols_6_14_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_216_io_enq_bits = cols_6_14_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_216_io_deq_ready = cols_7_14_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_217_clock = clock;
  assign q_217_reset = reset;
  assign q_217_io_enq_valid = cols_7_14_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_217_io_enq_bits = cols_7_14_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_217_io_deq_ready = cols_8_14_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_218_clock = clock;
  assign q_218_reset = reset;
  assign q_218_io_enq_valid = cols_8_14_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_218_io_enq_bits = cols_8_14_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_218_io_deq_ready = cols_9_14_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_219_clock = clock;
  assign q_219_reset = reset;
  assign q_219_io_enq_valid = cols_9_14_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_219_io_enq_bits = cols_9_14_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_219_io_deq_ready = cols_10_14_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_220_clock = clock;
  assign q_220_reset = reset;
  assign q_220_io_enq_valid = cols_10_14_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_220_io_enq_bits = cols_10_14_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_220_io_deq_ready = cols_11_14_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_221_clock = clock;
  assign q_221_reset = reset;
  assign q_221_io_enq_valid = cols_11_14_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_221_io_enq_bits = cols_11_14_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_221_io_deq_ready = cols_12_14_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_222_clock = clock;
  assign q_222_reset = reset;
  assign q_222_io_enq_valid = cols_12_14_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_222_io_enq_bits = cols_12_14_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_222_io_deq_ready = cols_13_14_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_223_clock = clock;
  assign q_223_reset = reset;
  assign q_223_io_enq_valid = cols_13_14_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_223_io_enq_bits = cols_13_14_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_223_io_deq_ready = cols_14_14_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_224_clock = clock;
  assign q_224_reset = reset;
  assign q_224_io_enq_valid = cols_14_14_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_224_io_enq_bits = cols_14_14_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_224_io_deq_ready = cols_15_14_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_225_clock = clock;
  assign q_225_reset = reset;
  assign q_225_io_enq_valid = cols_0_15_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_225_io_enq_bits = cols_0_15_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_225_io_deq_ready = cols_1_15_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_226_clock = clock;
  assign q_226_reset = reset;
  assign q_226_io_enq_valid = cols_1_15_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_226_io_enq_bits = cols_1_15_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_226_io_deq_ready = cols_2_15_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_227_clock = clock;
  assign q_227_reset = reset;
  assign q_227_io_enq_valid = cols_2_15_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_227_io_enq_bits = cols_2_15_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_227_io_deq_ready = cols_3_15_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_228_clock = clock;
  assign q_228_reset = reset;
  assign q_228_io_enq_valid = cols_3_15_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_228_io_enq_bits = cols_3_15_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_228_io_deq_ready = cols_4_15_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_229_clock = clock;
  assign q_229_reset = reset;
  assign q_229_io_enq_valid = cols_4_15_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_229_io_enq_bits = cols_4_15_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_229_io_deq_ready = cols_5_15_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_230_clock = clock;
  assign q_230_reset = reset;
  assign q_230_io_enq_valid = cols_5_15_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_230_io_enq_bits = cols_5_15_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_230_io_deq_ready = cols_6_15_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_231_clock = clock;
  assign q_231_reset = reset;
  assign q_231_io_enq_valid = cols_6_15_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_231_io_enq_bits = cols_6_15_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_231_io_deq_ready = cols_7_15_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_232_clock = clock;
  assign q_232_reset = reset;
  assign q_232_io_enq_valid = cols_7_15_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_232_io_enq_bits = cols_7_15_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_232_io_deq_ready = cols_8_15_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_233_clock = clock;
  assign q_233_reset = reset;
  assign q_233_io_enq_valid = cols_8_15_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_233_io_enq_bits = cols_8_15_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_233_io_deq_ready = cols_9_15_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_234_clock = clock;
  assign q_234_reset = reset;
  assign q_234_io_enq_valid = cols_9_15_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_234_io_enq_bits = cols_9_15_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_234_io_deq_ready = cols_10_15_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_235_clock = clock;
  assign q_235_reset = reset;
  assign q_235_io_enq_valid = cols_10_15_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_235_io_enq_bits = cols_10_15_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_235_io_deq_ready = cols_11_15_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_236_clock = clock;
  assign q_236_reset = reset;
  assign q_236_io_enq_valid = cols_11_15_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_236_io_enq_bits = cols_11_15_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_236_io_deq_ready = cols_12_15_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_237_clock = clock;
  assign q_237_reset = reset;
  assign q_237_io_enq_valid = cols_12_15_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_237_io_enq_bits = cols_12_15_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_237_io_deq_ready = cols_13_15_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_238_clock = clock;
  assign q_238_reset = reset;
  assign q_238_io_enq_valid = cols_13_15_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_238_io_enq_bits = cols_13_15_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_238_io_deq_ready = cols_14_15_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_239_clock = clock;
  assign q_239_reset = reset;
  assign q_239_io_enq_valid = cols_14_15_io_right_out_valid; // @[Decoupled.scala 363:22]
  assign q_239_io_enq_bits = cols_14_15_io_right_out_bits; // @[Decoupled.scala 364:21]
  assign q_239_io_deq_ready = cols_15_15_io_left_in_ready; // @[Stab.scala 89:69]
  assign q_240_clock = clock;
  assign q_240_reset = reset;
  assign q_240_io_enq_valid = io_weight_in_0_valid; // @[Decoupled.scala 363:22]
  assign q_240_io_enq_bits = io_weight_in_0_bits; // @[Decoupled.scala 364:21]
  assign q_240_io_deq_ready = cols_0_0_io_top_in_ready; // @[Stab.scala 93:102]
  assign q_241_clock = clock;
  assign q_241_reset = reset;
  assign q_241_io_enq_valid = io_weight_in_1_valid; // @[Decoupled.scala 363:22]
  assign q_241_io_enq_bits = io_weight_in_1_bits; // @[Decoupled.scala 364:21]
  assign q_241_io_deq_ready = cols_1_0_io_top_in_ready; // @[Stab.scala 93:102]
  assign q_242_clock = clock;
  assign q_242_reset = reset;
  assign q_242_io_enq_valid = io_weight_in_2_valid; // @[Decoupled.scala 363:22]
  assign q_242_io_enq_bits = io_weight_in_2_bits; // @[Decoupled.scala 364:21]
  assign q_242_io_deq_ready = cols_2_0_io_top_in_ready; // @[Stab.scala 93:102]
  assign q_243_clock = clock;
  assign q_243_reset = reset;
  assign q_243_io_enq_valid = io_weight_in_3_valid; // @[Decoupled.scala 363:22]
  assign q_243_io_enq_bits = io_weight_in_3_bits; // @[Decoupled.scala 364:21]
  assign q_243_io_deq_ready = cols_3_0_io_top_in_ready; // @[Stab.scala 93:102]
  assign q_244_clock = clock;
  assign q_244_reset = reset;
  assign q_244_io_enq_valid = io_weight_in_4_valid; // @[Decoupled.scala 363:22]
  assign q_244_io_enq_bits = io_weight_in_4_bits; // @[Decoupled.scala 364:21]
  assign q_244_io_deq_ready = cols_4_0_io_top_in_ready; // @[Stab.scala 93:102]
  assign q_245_clock = clock;
  assign q_245_reset = reset;
  assign q_245_io_enq_valid = io_weight_in_5_valid; // @[Decoupled.scala 363:22]
  assign q_245_io_enq_bits = io_weight_in_5_bits; // @[Decoupled.scala 364:21]
  assign q_245_io_deq_ready = cols_5_0_io_top_in_ready; // @[Stab.scala 93:102]
  assign q_246_clock = clock;
  assign q_246_reset = reset;
  assign q_246_io_enq_valid = io_weight_in_6_valid; // @[Decoupled.scala 363:22]
  assign q_246_io_enq_bits = io_weight_in_6_bits; // @[Decoupled.scala 364:21]
  assign q_246_io_deq_ready = cols_6_0_io_top_in_ready; // @[Stab.scala 93:102]
  assign q_247_clock = clock;
  assign q_247_reset = reset;
  assign q_247_io_enq_valid = io_weight_in_7_valid; // @[Decoupled.scala 363:22]
  assign q_247_io_enq_bits = io_weight_in_7_bits; // @[Decoupled.scala 364:21]
  assign q_247_io_deq_ready = cols_7_0_io_top_in_ready; // @[Stab.scala 93:102]
  assign q_248_clock = clock;
  assign q_248_reset = reset;
  assign q_248_io_enq_valid = io_weight_in_8_valid; // @[Decoupled.scala 363:22]
  assign q_248_io_enq_bits = io_weight_in_8_bits; // @[Decoupled.scala 364:21]
  assign q_248_io_deq_ready = cols_8_0_io_top_in_ready; // @[Stab.scala 93:102]
  assign q_249_clock = clock;
  assign q_249_reset = reset;
  assign q_249_io_enq_valid = io_weight_in_9_valid; // @[Decoupled.scala 363:22]
  assign q_249_io_enq_bits = io_weight_in_9_bits; // @[Decoupled.scala 364:21]
  assign q_249_io_deq_ready = cols_9_0_io_top_in_ready; // @[Stab.scala 93:102]
  assign q_250_clock = clock;
  assign q_250_reset = reset;
  assign q_250_io_enq_valid = io_weight_in_10_valid; // @[Decoupled.scala 363:22]
  assign q_250_io_enq_bits = io_weight_in_10_bits; // @[Decoupled.scala 364:21]
  assign q_250_io_deq_ready = cols_10_0_io_top_in_ready; // @[Stab.scala 93:102]
  assign q_251_clock = clock;
  assign q_251_reset = reset;
  assign q_251_io_enq_valid = io_weight_in_11_valid; // @[Decoupled.scala 363:22]
  assign q_251_io_enq_bits = io_weight_in_11_bits; // @[Decoupled.scala 364:21]
  assign q_251_io_deq_ready = cols_11_0_io_top_in_ready; // @[Stab.scala 93:102]
  assign q_252_clock = clock;
  assign q_252_reset = reset;
  assign q_252_io_enq_valid = io_weight_in_12_valid; // @[Decoupled.scala 363:22]
  assign q_252_io_enq_bits = io_weight_in_12_bits; // @[Decoupled.scala 364:21]
  assign q_252_io_deq_ready = cols_12_0_io_top_in_ready; // @[Stab.scala 93:102]
  assign q_253_clock = clock;
  assign q_253_reset = reset;
  assign q_253_io_enq_valid = io_weight_in_13_valid; // @[Decoupled.scala 363:22]
  assign q_253_io_enq_bits = io_weight_in_13_bits; // @[Decoupled.scala 364:21]
  assign q_253_io_deq_ready = cols_13_0_io_top_in_ready; // @[Stab.scala 93:102]
  assign q_254_clock = clock;
  assign q_254_reset = reset;
  assign q_254_io_enq_valid = io_weight_in_14_valid; // @[Decoupled.scala 363:22]
  assign q_254_io_enq_bits = io_weight_in_14_bits; // @[Decoupled.scala 364:21]
  assign q_254_io_deq_ready = cols_14_0_io_top_in_ready; // @[Stab.scala 93:102]
  assign q_255_clock = clock;
  assign q_255_reset = reset;
  assign q_255_io_enq_valid = io_weight_in_15_valid; // @[Decoupled.scala 363:22]
  assign q_255_io_enq_bits = io_weight_in_15_bits; // @[Decoupled.scala 364:21]
  assign q_255_io_deq_ready = cols_15_0_io_top_in_ready; // @[Stab.scala 93:102]
  assign q_256_clock = clock;
  assign q_256_reset = reset;
  assign q_256_io_enq_valid = cols_0_0_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_256_io_enq_bits = cols_0_0_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_256_io_deq_ready = cols_0_1_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_257_clock = clock;
  assign q_257_reset = reset;
  assign q_257_io_enq_valid = cols_0_1_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_257_io_enq_bits = cols_0_1_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_257_io_deq_ready = cols_0_2_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_258_clock = clock;
  assign q_258_reset = reset;
  assign q_258_io_enq_valid = cols_0_2_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_258_io_enq_bits = cols_0_2_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_258_io_deq_ready = cols_0_3_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_259_clock = clock;
  assign q_259_reset = reset;
  assign q_259_io_enq_valid = cols_0_3_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_259_io_enq_bits = cols_0_3_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_259_io_deq_ready = cols_0_4_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_260_clock = clock;
  assign q_260_reset = reset;
  assign q_260_io_enq_valid = cols_0_4_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_260_io_enq_bits = cols_0_4_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_260_io_deq_ready = cols_0_5_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_261_clock = clock;
  assign q_261_reset = reset;
  assign q_261_io_enq_valid = cols_0_5_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_261_io_enq_bits = cols_0_5_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_261_io_deq_ready = cols_0_6_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_262_clock = clock;
  assign q_262_reset = reset;
  assign q_262_io_enq_valid = cols_0_6_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_262_io_enq_bits = cols_0_6_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_262_io_deq_ready = cols_0_7_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_263_clock = clock;
  assign q_263_reset = reset;
  assign q_263_io_enq_valid = cols_0_7_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_263_io_enq_bits = cols_0_7_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_263_io_deq_ready = cols_0_8_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_264_clock = clock;
  assign q_264_reset = reset;
  assign q_264_io_enq_valid = cols_0_8_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_264_io_enq_bits = cols_0_8_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_264_io_deq_ready = cols_0_9_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_265_clock = clock;
  assign q_265_reset = reset;
  assign q_265_io_enq_valid = cols_0_9_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_265_io_enq_bits = cols_0_9_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_265_io_deq_ready = cols_0_10_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_266_clock = clock;
  assign q_266_reset = reset;
  assign q_266_io_enq_valid = cols_0_10_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_266_io_enq_bits = cols_0_10_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_266_io_deq_ready = cols_0_11_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_267_clock = clock;
  assign q_267_reset = reset;
  assign q_267_io_enq_valid = cols_0_11_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_267_io_enq_bits = cols_0_11_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_267_io_deq_ready = cols_0_12_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_268_clock = clock;
  assign q_268_reset = reset;
  assign q_268_io_enq_valid = cols_0_12_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_268_io_enq_bits = cols_0_12_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_268_io_deq_ready = cols_0_13_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_269_clock = clock;
  assign q_269_reset = reset;
  assign q_269_io_enq_valid = cols_0_13_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_269_io_enq_bits = cols_0_13_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_269_io_deq_ready = cols_0_14_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_270_clock = clock;
  assign q_270_reset = reset;
  assign q_270_io_enq_valid = cols_0_14_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_270_io_enq_bits = cols_0_14_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_270_io_deq_ready = cols_0_15_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_271_clock = clock;
  assign q_271_reset = reset;
  assign q_271_io_enq_valid = cols_1_0_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_271_io_enq_bits = cols_1_0_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_271_io_deq_ready = cols_1_1_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_272_clock = clock;
  assign q_272_reset = reset;
  assign q_272_io_enq_valid = cols_1_1_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_272_io_enq_bits = cols_1_1_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_272_io_deq_ready = cols_1_2_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_273_clock = clock;
  assign q_273_reset = reset;
  assign q_273_io_enq_valid = cols_1_2_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_273_io_enq_bits = cols_1_2_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_273_io_deq_ready = cols_1_3_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_274_clock = clock;
  assign q_274_reset = reset;
  assign q_274_io_enq_valid = cols_1_3_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_274_io_enq_bits = cols_1_3_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_274_io_deq_ready = cols_1_4_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_275_clock = clock;
  assign q_275_reset = reset;
  assign q_275_io_enq_valid = cols_1_4_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_275_io_enq_bits = cols_1_4_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_275_io_deq_ready = cols_1_5_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_276_clock = clock;
  assign q_276_reset = reset;
  assign q_276_io_enq_valid = cols_1_5_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_276_io_enq_bits = cols_1_5_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_276_io_deq_ready = cols_1_6_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_277_clock = clock;
  assign q_277_reset = reset;
  assign q_277_io_enq_valid = cols_1_6_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_277_io_enq_bits = cols_1_6_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_277_io_deq_ready = cols_1_7_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_278_clock = clock;
  assign q_278_reset = reset;
  assign q_278_io_enq_valid = cols_1_7_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_278_io_enq_bits = cols_1_7_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_278_io_deq_ready = cols_1_8_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_279_clock = clock;
  assign q_279_reset = reset;
  assign q_279_io_enq_valid = cols_1_8_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_279_io_enq_bits = cols_1_8_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_279_io_deq_ready = cols_1_9_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_280_clock = clock;
  assign q_280_reset = reset;
  assign q_280_io_enq_valid = cols_1_9_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_280_io_enq_bits = cols_1_9_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_280_io_deq_ready = cols_1_10_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_281_clock = clock;
  assign q_281_reset = reset;
  assign q_281_io_enq_valid = cols_1_10_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_281_io_enq_bits = cols_1_10_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_281_io_deq_ready = cols_1_11_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_282_clock = clock;
  assign q_282_reset = reset;
  assign q_282_io_enq_valid = cols_1_11_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_282_io_enq_bits = cols_1_11_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_282_io_deq_ready = cols_1_12_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_283_clock = clock;
  assign q_283_reset = reset;
  assign q_283_io_enq_valid = cols_1_12_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_283_io_enq_bits = cols_1_12_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_283_io_deq_ready = cols_1_13_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_284_clock = clock;
  assign q_284_reset = reset;
  assign q_284_io_enq_valid = cols_1_13_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_284_io_enq_bits = cols_1_13_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_284_io_deq_ready = cols_1_14_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_285_clock = clock;
  assign q_285_reset = reset;
  assign q_285_io_enq_valid = cols_1_14_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_285_io_enq_bits = cols_1_14_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_285_io_deq_ready = cols_1_15_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_286_clock = clock;
  assign q_286_reset = reset;
  assign q_286_io_enq_valid = cols_2_0_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_286_io_enq_bits = cols_2_0_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_286_io_deq_ready = cols_2_1_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_287_clock = clock;
  assign q_287_reset = reset;
  assign q_287_io_enq_valid = cols_2_1_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_287_io_enq_bits = cols_2_1_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_287_io_deq_ready = cols_2_2_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_288_clock = clock;
  assign q_288_reset = reset;
  assign q_288_io_enq_valid = cols_2_2_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_288_io_enq_bits = cols_2_2_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_288_io_deq_ready = cols_2_3_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_289_clock = clock;
  assign q_289_reset = reset;
  assign q_289_io_enq_valid = cols_2_3_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_289_io_enq_bits = cols_2_3_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_289_io_deq_ready = cols_2_4_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_290_clock = clock;
  assign q_290_reset = reset;
  assign q_290_io_enq_valid = cols_2_4_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_290_io_enq_bits = cols_2_4_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_290_io_deq_ready = cols_2_5_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_291_clock = clock;
  assign q_291_reset = reset;
  assign q_291_io_enq_valid = cols_2_5_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_291_io_enq_bits = cols_2_5_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_291_io_deq_ready = cols_2_6_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_292_clock = clock;
  assign q_292_reset = reset;
  assign q_292_io_enq_valid = cols_2_6_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_292_io_enq_bits = cols_2_6_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_292_io_deq_ready = cols_2_7_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_293_clock = clock;
  assign q_293_reset = reset;
  assign q_293_io_enq_valid = cols_2_7_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_293_io_enq_bits = cols_2_7_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_293_io_deq_ready = cols_2_8_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_294_clock = clock;
  assign q_294_reset = reset;
  assign q_294_io_enq_valid = cols_2_8_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_294_io_enq_bits = cols_2_8_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_294_io_deq_ready = cols_2_9_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_295_clock = clock;
  assign q_295_reset = reset;
  assign q_295_io_enq_valid = cols_2_9_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_295_io_enq_bits = cols_2_9_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_295_io_deq_ready = cols_2_10_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_296_clock = clock;
  assign q_296_reset = reset;
  assign q_296_io_enq_valid = cols_2_10_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_296_io_enq_bits = cols_2_10_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_296_io_deq_ready = cols_2_11_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_297_clock = clock;
  assign q_297_reset = reset;
  assign q_297_io_enq_valid = cols_2_11_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_297_io_enq_bits = cols_2_11_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_297_io_deq_ready = cols_2_12_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_298_clock = clock;
  assign q_298_reset = reset;
  assign q_298_io_enq_valid = cols_2_12_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_298_io_enq_bits = cols_2_12_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_298_io_deq_ready = cols_2_13_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_299_clock = clock;
  assign q_299_reset = reset;
  assign q_299_io_enq_valid = cols_2_13_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_299_io_enq_bits = cols_2_13_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_299_io_deq_ready = cols_2_14_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_300_clock = clock;
  assign q_300_reset = reset;
  assign q_300_io_enq_valid = cols_2_14_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_300_io_enq_bits = cols_2_14_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_300_io_deq_ready = cols_2_15_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_301_clock = clock;
  assign q_301_reset = reset;
  assign q_301_io_enq_valid = cols_3_0_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_301_io_enq_bits = cols_3_0_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_301_io_deq_ready = cols_3_1_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_302_clock = clock;
  assign q_302_reset = reset;
  assign q_302_io_enq_valid = cols_3_1_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_302_io_enq_bits = cols_3_1_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_302_io_deq_ready = cols_3_2_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_303_clock = clock;
  assign q_303_reset = reset;
  assign q_303_io_enq_valid = cols_3_2_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_303_io_enq_bits = cols_3_2_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_303_io_deq_ready = cols_3_3_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_304_clock = clock;
  assign q_304_reset = reset;
  assign q_304_io_enq_valid = cols_3_3_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_304_io_enq_bits = cols_3_3_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_304_io_deq_ready = cols_3_4_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_305_clock = clock;
  assign q_305_reset = reset;
  assign q_305_io_enq_valid = cols_3_4_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_305_io_enq_bits = cols_3_4_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_305_io_deq_ready = cols_3_5_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_306_clock = clock;
  assign q_306_reset = reset;
  assign q_306_io_enq_valid = cols_3_5_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_306_io_enq_bits = cols_3_5_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_306_io_deq_ready = cols_3_6_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_307_clock = clock;
  assign q_307_reset = reset;
  assign q_307_io_enq_valid = cols_3_6_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_307_io_enq_bits = cols_3_6_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_307_io_deq_ready = cols_3_7_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_308_clock = clock;
  assign q_308_reset = reset;
  assign q_308_io_enq_valid = cols_3_7_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_308_io_enq_bits = cols_3_7_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_308_io_deq_ready = cols_3_8_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_309_clock = clock;
  assign q_309_reset = reset;
  assign q_309_io_enq_valid = cols_3_8_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_309_io_enq_bits = cols_3_8_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_309_io_deq_ready = cols_3_9_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_310_clock = clock;
  assign q_310_reset = reset;
  assign q_310_io_enq_valid = cols_3_9_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_310_io_enq_bits = cols_3_9_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_310_io_deq_ready = cols_3_10_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_311_clock = clock;
  assign q_311_reset = reset;
  assign q_311_io_enq_valid = cols_3_10_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_311_io_enq_bits = cols_3_10_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_311_io_deq_ready = cols_3_11_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_312_clock = clock;
  assign q_312_reset = reset;
  assign q_312_io_enq_valid = cols_3_11_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_312_io_enq_bits = cols_3_11_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_312_io_deq_ready = cols_3_12_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_313_clock = clock;
  assign q_313_reset = reset;
  assign q_313_io_enq_valid = cols_3_12_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_313_io_enq_bits = cols_3_12_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_313_io_deq_ready = cols_3_13_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_314_clock = clock;
  assign q_314_reset = reset;
  assign q_314_io_enq_valid = cols_3_13_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_314_io_enq_bits = cols_3_13_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_314_io_deq_ready = cols_3_14_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_315_clock = clock;
  assign q_315_reset = reset;
  assign q_315_io_enq_valid = cols_3_14_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_315_io_enq_bits = cols_3_14_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_315_io_deq_ready = cols_3_15_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_316_clock = clock;
  assign q_316_reset = reset;
  assign q_316_io_enq_valid = cols_4_0_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_316_io_enq_bits = cols_4_0_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_316_io_deq_ready = cols_4_1_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_317_clock = clock;
  assign q_317_reset = reset;
  assign q_317_io_enq_valid = cols_4_1_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_317_io_enq_bits = cols_4_1_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_317_io_deq_ready = cols_4_2_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_318_clock = clock;
  assign q_318_reset = reset;
  assign q_318_io_enq_valid = cols_4_2_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_318_io_enq_bits = cols_4_2_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_318_io_deq_ready = cols_4_3_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_319_clock = clock;
  assign q_319_reset = reset;
  assign q_319_io_enq_valid = cols_4_3_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_319_io_enq_bits = cols_4_3_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_319_io_deq_ready = cols_4_4_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_320_clock = clock;
  assign q_320_reset = reset;
  assign q_320_io_enq_valid = cols_4_4_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_320_io_enq_bits = cols_4_4_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_320_io_deq_ready = cols_4_5_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_321_clock = clock;
  assign q_321_reset = reset;
  assign q_321_io_enq_valid = cols_4_5_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_321_io_enq_bits = cols_4_5_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_321_io_deq_ready = cols_4_6_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_322_clock = clock;
  assign q_322_reset = reset;
  assign q_322_io_enq_valid = cols_4_6_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_322_io_enq_bits = cols_4_6_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_322_io_deq_ready = cols_4_7_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_323_clock = clock;
  assign q_323_reset = reset;
  assign q_323_io_enq_valid = cols_4_7_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_323_io_enq_bits = cols_4_7_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_323_io_deq_ready = cols_4_8_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_324_clock = clock;
  assign q_324_reset = reset;
  assign q_324_io_enq_valid = cols_4_8_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_324_io_enq_bits = cols_4_8_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_324_io_deq_ready = cols_4_9_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_325_clock = clock;
  assign q_325_reset = reset;
  assign q_325_io_enq_valid = cols_4_9_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_325_io_enq_bits = cols_4_9_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_325_io_deq_ready = cols_4_10_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_326_clock = clock;
  assign q_326_reset = reset;
  assign q_326_io_enq_valid = cols_4_10_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_326_io_enq_bits = cols_4_10_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_326_io_deq_ready = cols_4_11_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_327_clock = clock;
  assign q_327_reset = reset;
  assign q_327_io_enq_valid = cols_4_11_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_327_io_enq_bits = cols_4_11_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_327_io_deq_ready = cols_4_12_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_328_clock = clock;
  assign q_328_reset = reset;
  assign q_328_io_enq_valid = cols_4_12_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_328_io_enq_bits = cols_4_12_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_328_io_deq_ready = cols_4_13_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_329_clock = clock;
  assign q_329_reset = reset;
  assign q_329_io_enq_valid = cols_4_13_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_329_io_enq_bits = cols_4_13_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_329_io_deq_ready = cols_4_14_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_330_clock = clock;
  assign q_330_reset = reset;
  assign q_330_io_enq_valid = cols_4_14_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_330_io_enq_bits = cols_4_14_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_330_io_deq_ready = cols_4_15_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_331_clock = clock;
  assign q_331_reset = reset;
  assign q_331_io_enq_valid = cols_5_0_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_331_io_enq_bits = cols_5_0_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_331_io_deq_ready = cols_5_1_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_332_clock = clock;
  assign q_332_reset = reset;
  assign q_332_io_enq_valid = cols_5_1_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_332_io_enq_bits = cols_5_1_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_332_io_deq_ready = cols_5_2_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_333_clock = clock;
  assign q_333_reset = reset;
  assign q_333_io_enq_valid = cols_5_2_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_333_io_enq_bits = cols_5_2_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_333_io_deq_ready = cols_5_3_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_334_clock = clock;
  assign q_334_reset = reset;
  assign q_334_io_enq_valid = cols_5_3_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_334_io_enq_bits = cols_5_3_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_334_io_deq_ready = cols_5_4_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_335_clock = clock;
  assign q_335_reset = reset;
  assign q_335_io_enq_valid = cols_5_4_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_335_io_enq_bits = cols_5_4_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_335_io_deq_ready = cols_5_5_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_336_clock = clock;
  assign q_336_reset = reset;
  assign q_336_io_enq_valid = cols_5_5_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_336_io_enq_bits = cols_5_5_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_336_io_deq_ready = cols_5_6_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_337_clock = clock;
  assign q_337_reset = reset;
  assign q_337_io_enq_valid = cols_5_6_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_337_io_enq_bits = cols_5_6_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_337_io_deq_ready = cols_5_7_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_338_clock = clock;
  assign q_338_reset = reset;
  assign q_338_io_enq_valid = cols_5_7_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_338_io_enq_bits = cols_5_7_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_338_io_deq_ready = cols_5_8_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_339_clock = clock;
  assign q_339_reset = reset;
  assign q_339_io_enq_valid = cols_5_8_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_339_io_enq_bits = cols_5_8_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_339_io_deq_ready = cols_5_9_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_340_clock = clock;
  assign q_340_reset = reset;
  assign q_340_io_enq_valid = cols_5_9_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_340_io_enq_bits = cols_5_9_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_340_io_deq_ready = cols_5_10_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_341_clock = clock;
  assign q_341_reset = reset;
  assign q_341_io_enq_valid = cols_5_10_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_341_io_enq_bits = cols_5_10_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_341_io_deq_ready = cols_5_11_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_342_clock = clock;
  assign q_342_reset = reset;
  assign q_342_io_enq_valid = cols_5_11_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_342_io_enq_bits = cols_5_11_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_342_io_deq_ready = cols_5_12_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_343_clock = clock;
  assign q_343_reset = reset;
  assign q_343_io_enq_valid = cols_5_12_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_343_io_enq_bits = cols_5_12_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_343_io_deq_ready = cols_5_13_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_344_clock = clock;
  assign q_344_reset = reset;
  assign q_344_io_enq_valid = cols_5_13_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_344_io_enq_bits = cols_5_13_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_344_io_deq_ready = cols_5_14_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_345_clock = clock;
  assign q_345_reset = reset;
  assign q_345_io_enq_valid = cols_5_14_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_345_io_enq_bits = cols_5_14_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_345_io_deq_ready = cols_5_15_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_346_clock = clock;
  assign q_346_reset = reset;
  assign q_346_io_enq_valid = cols_6_0_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_346_io_enq_bits = cols_6_0_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_346_io_deq_ready = cols_6_1_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_347_clock = clock;
  assign q_347_reset = reset;
  assign q_347_io_enq_valid = cols_6_1_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_347_io_enq_bits = cols_6_1_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_347_io_deq_ready = cols_6_2_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_348_clock = clock;
  assign q_348_reset = reset;
  assign q_348_io_enq_valid = cols_6_2_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_348_io_enq_bits = cols_6_2_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_348_io_deq_ready = cols_6_3_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_349_clock = clock;
  assign q_349_reset = reset;
  assign q_349_io_enq_valid = cols_6_3_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_349_io_enq_bits = cols_6_3_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_349_io_deq_ready = cols_6_4_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_350_clock = clock;
  assign q_350_reset = reset;
  assign q_350_io_enq_valid = cols_6_4_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_350_io_enq_bits = cols_6_4_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_350_io_deq_ready = cols_6_5_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_351_clock = clock;
  assign q_351_reset = reset;
  assign q_351_io_enq_valid = cols_6_5_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_351_io_enq_bits = cols_6_5_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_351_io_deq_ready = cols_6_6_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_352_clock = clock;
  assign q_352_reset = reset;
  assign q_352_io_enq_valid = cols_6_6_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_352_io_enq_bits = cols_6_6_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_352_io_deq_ready = cols_6_7_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_353_clock = clock;
  assign q_353_reset = reset;
  assign q_353_io_enq_valid = cols_6_7_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_353_io_enq_bits = cols_6_7_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_353_io_deq_ready = cols_6_8_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_354_clock = clock;
  assign q_354_reset = reset;
  assign q_354_io_enq_valid = cols_6_8_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_354_io_enq_bits = cols_6_8_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_354_io_deq_ready = cols_6_9_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_355_clock = clock;
  assign q_355_reset = reset;
  assign q_355_io_enq_valid = cols_6_9_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_355_io_enq_bits = cols_6_9_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_355_io_deq_ready = cols_6_10_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_356_clock = clock;
  assign q_356_reset = reset;
  assign q_356_io_enq_valid = cols_6_10_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_356_io_enq_bits = cols_6_10_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_356_io_deq_ready = cols_6_11_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_357_clock = clock;
  assign q_357_reset = reset;
  assign q_357_io_enq_valid = cols_6_11_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_357_io_enq_bits = cols_6_11_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_357_io_deq_ready = cols_6_12_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_358_clock = clock;
  assign q_358_reset = reset;
  assign q_358_io_enq_valid = cols_6_12_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_358_io_enq_bits = cols_6_12_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_358_io_deq_ready = cols_6_13_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_359_clock = clock;
  assign q_359_reset = reset;
  assign q_359_io_enq_valid = cols_6_13_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_359_io_enq_bits = cols_6_13_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_359_io_deq_ready = cols_6_14_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_360_clock = clock;
  assign q_360_reset = reset;
  assign q_360_io_enq_valid = cols_6_14_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_360_io_enq_bits = cols_6_14_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_360_io_deq_ready = cols_6_15_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_361_clock = clock;
  assign q_361_reset = reset;
  assign q_361_io_enq_valid = cols_7_0_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_361_io_enq_bits = cols_7_0_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_361_io_deq_ready = cols_7_1_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_362_clock = clock;
  assign q_362_reset = reset;
  assign q_362_io_enq_valid = cols_7_1_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_362_io_enq_bits = cols_7_1_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_362_io_deq_ready = cols_7_2_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_363_clock = clock;
  assign q_363_reset = reset;
  assign q_363_io_enq_valid = cols_7_2_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_363_io_enq_bits = cols_7_2_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_363_io_deq_ready = cols_7_3_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_364_clock = clock;
  assign q_364_reset = reset;
  assign q_364_io_enq_valid = cols_7_3_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_364_io_enq_bits = cols_7_3_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_364_io_deq_ready = cols_7_4_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_365_clock = clock;
  assign q_365_reset = reset;
  assign q_365_io_enq_valid = cols_7_4_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_365_io_enq_bits = cols_7_4_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_365_io_deq_ready = cols_7_5_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_366_clock = clock;
  assign q_366_reset = reset;
  assign q_366_io_enq_valid = cols_7_5_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_366_io_enq_bits = cols_7_5_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_366_io_deq_ready = cols_7_6_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_367_clock = clock;
  assign q_367_reset = reset;
  assign q_367_io_enq_valid = cols_7_6_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_367_io_enq_bits = cols_7_6_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_367_io_deq_ready = cols_7_7_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_368_clock = clock;
  assign q_368_reset = reset;
  assign q_368_io_enq_valid = cols_7_7_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_368_io_enq_bits = cols_7_7_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_368_io_deq_ready = cols_7_8_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_369_clock = clock;
  assign q_369_reset = reset;
  assign q_369_io_enq_valid = cols_7_8_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_369_io_enq_bits = cols_7_8_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_369_io_deq_ready = cols_7_9_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_370_clock = clock;
  assign q_370_reset = reset;
  assign q_370_io_enq_valid = cols_7_9_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_370_io_enq_bits = cols_7_9_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_370_io_deq_ready = cols_7_10_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_371_clock = clock;
  assign q_371_reset = reset;
  assign q_371_io_enq_valid = cols_7_10_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_371_io_enq_bits = cols_7_10_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_371_io_deq_ready = cols_7_11_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_372_clock = clock;
  assign q_372_reset = reset;
  assign q_372_io_enq_valid = cols_7_11_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_372_io_enq_bits = cols_7_11_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_372_io_deq_ready = cols_7_12_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_373_clock = clock;
  assign q_373_reset = reset;
  assign q_373_io_enq_valid = cols_7_12_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_373_io_enq_bits = cols_7_12_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_373_io_deq_ready = cols_7_13_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_374_clock = clock;
  assign q_374_reset = reset;
  assign q_374_io_enq_valid = cols_7_13_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_374_io_enq_bits = cols_7_13_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_374_io_deq_ready = cols_7_14_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_375_clock = clock;
  assign q_375_reset = reset;
  assign q_375_io_enq_valid = cols_7_14_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_375_io_enq_bits = cols_7_14_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_375_io_deq_ready = cols_7_15_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_376_clock = clock;
  assign q_376_reset = reset;
  assign q_376_io_enq_valid = cols_8_0_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_376_io_enq_bits = cols_8_0_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_376_io_deq_ready = cols_8_1_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_377_clock = clock;
  assign q_377_reset = reset;
  assign q_377_io_enq_valid = cols_8_1_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_377_io_enq_bits = cols_8_1_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_377_io_deq_ready = cols_8_2_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_378_clock = clock;
  assign q_378_reset = reset;
  assign q_378_io_enq_valid = cols_8_2_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_378_io_enq_bits = cols_8_2_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_378_io_deq_ready = cols_8_3_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_379_clock = clock;
  assign q_379_reset = reset;
  assign q_379_io_enq_valid = cols_8_3_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_379_io_enq_bits = cols_8_3_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_379_io_deq_ready = cols_8_4_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_380_clock = clock;
  assign q_380_reset = reset;
  assign q_380_io_enq_valid = cols_8_4_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_380_io_enq_bits = cols_8_4_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_380_io_deq_ready = cols_8_5_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_381_clock = clock;
  assign q_381_reset = reset;
  assign q_381_io_enq_valid = cols_8_5_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_381_io_enq_bits = cols_8_5_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_381_io_deq_ready = cols_8_6_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_382_clock = clock;
  assign q_382_reset = reset;
  assign q_382_io_enq_valid = cols_8_6_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_382_io_enq_bits = cols_8_6_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_382_io_deq_ready = cols_8_7_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_383_clock = clock;
  assign q_383_reset = reset;
  assign q_383_io_enq_valid = cols_8_7_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_383_io_enq_bits = cols_8_7_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_383_io_deq_ready = cols_8_8_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_384_clock = clock;
  assign q_384_reset = reset;
  assign q_384_io_enq_valid = cols_8_8_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_384_io_enq_bits = cols_8_8_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_384_io_deq_ready = cols_8_9_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_385_clock = clock;
  assign q_385_reset = reset;
  assign q_385_io_enq_valid = cols_8_9_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_385_io_enq_bits = cols_8_9_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_385_io_deq_ready = cols_8_10_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_386_clock = clock;
  assign q_386_reset = reset;
  assign q_386_io_enq_valid = cols_8_10_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_386_io_enq_bits = cols_8_10_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_386_io_deq_ready = cols_8_11_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_387_clock = clock;
  assign q_387_reset = reset;
  assign q_387_io_enq_valid = cols_8_11_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_387_io_enq_bits = cols_8_11_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_387_io_deq_ready = cols_8_12_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_388_clock = clock;
  assign q_388_reset = reset;
  assign q_388_io_enq_valid = cols_8_12_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_388_io_enq_bits = cols_8_12_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_388_io_deq_ready = cols_8_13_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_389_clock = clock;
  assign q_389_reset = reset;
  assign q_389_io_enq_valid = cols_8_13_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_389_io_enq_bits = cols_8_13_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_389_io_deq_ready = cols_8_14_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_390_clock = clock;
  assign q_390_reset = reset;
  assign q_390_io_enq_valid = cols_8_14_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_390_io_enq_bits = cols_8_14_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_390_io_deq_ready = cols_8_15_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_391_clock = clock;
  assign q_391_reset = reset;
  assign q_391_io_enq_valid = cols_9_0_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_391_io_enq_bits = cols_9_0_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_391_io_deq_ready = cols_9_1_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_392_clock = clock;
  assign q_392_reset = reset;
  assign q_392_io_enq_valid = cols_9_1_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_392_io_enq_bits = cols_9_1_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_392_io_deq_ready = cols_9_2_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_393_clock = clock;
  assign q_393_reset = reset;
  assign q_393_io_enq_valid = cols_9_2_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_393_io_enq_bits = cols_9_2_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_393_io_deq_ready = cols_9_3_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_394_clock = clock;
  assign q_394_reset = reset;
  assign q_394_io_enq_valid = cols_9_3_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_394_io_enq_bits = cols_9_3_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_394_io_deq_ready = cols_9_4_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_395_clock = clock;
  assign q_395_reset = reset;
  assign q_395_io_enq_valid = cols_9_4_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_395_io_enq_bits = cols_9_4_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_395_io_deq_ready = cols_9_5_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_396_clock = clock;
  assign q_396_reset = reset;
  assign q_396_io_enq_valid = cols_9_5_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_396_io_enq_bits = cols_9_5_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_396_io_deq_ready = cols_9_6_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_397_clock = clock;
  assign q_397_reset = reset;
  assign q_397_io_enq_valid = cols_9_6_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_397_io_enq_bits = cols_9_6_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_397_io_deq_ready = cols_9_7_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_398_clock = clock;
  assign q_398_reset = reset;
  assign q_398_io_enq_valid = cols_9_7_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_398_io_enq_bits = cols_9_7_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_398_io_deq_ready = cols_9_8_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_399_clock = clock;
  assign q_399_reset = reset;
  assign q_399_io_enq_valid = cols_9_8_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_399_io_enq_bits = cols_9_8_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_399_io_deq_ready = cols_9_9_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_400_clock = clock;
  assign q_400_reset = reset;
  assign q_400_io_enq_valid = cols_9_9_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_400_io_enq_bits = cols_9_9_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_400_io_deq_ready = cols_9_10_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_401_clock = clock;
  assign q_401_reset = reset;
  assign q_401_io_enq_valid = cols_9_10_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_401_io_enq_bits = cols_9_10_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_401_io_deq_ready = cols_9_11_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_402_clock = clock;
  assign q_402_reset = reset;
  assign q_402_io_enq_valid = cols_9_11_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_402_io_enq_bits = cols_9_11_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_402_io_deq_ready = cols_9_12_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_403_clock = clock;
  assign q_403_reset = reset;
  assign q_403_io_enq_valid = cols_9_12_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_403_io_enq_bits = cols_9_12_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_403_io_deq_ready = cols_9_13_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_404_clock = clock;
  assign q_404_reset = reset;
  assign q_404_io_enq_valid = cols_9_13_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_404_io_enq_bits = cols_9_13_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_404_io_deq_ready = cols_9_14_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_405_clock = clock;
  assign q_405_reset = reset;
  assign q_405_io_enq_valid = cols_9_14_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_405_io_enq_bits = cols_9_14_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_405_io_deq_ready = cols_9_15_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_406_clock = clock;
  assign q_406_reset = reset;
  assign q_406_io_enq_valid = cols_10_0_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_406_io_enq_bits = cols_10_0_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_406_io_deq_ready = cols_10_1_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_407_clock = clock;
  assign q_407_reset = reset;
  assign q_407_io_enq_valid = cols_10_1_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_407_io_enq_bits = cols_10_1_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_407_io_deq_ready = cols_10_2_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_408_clock = clock;
  assign q_408_reset = reset;
  assign q_408_io_enq_valid = cols_10_2_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_408_io_enq_bits = cols_10_2_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_408_io_deq_ready = cols_10_3_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_409_clock = clock;
  assign q_409_reset = reset;
  assign q_409_io_enq_valid = cols_10_3_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_409_io_enq_bits = cols_10_3_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_409_io_deq_ready = cols_10_4_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_410_clock = clock;
  assign q_410_reset = reset;
  assign q_410_io_enq_valid = cols_10_4_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_410_io_enq_bits = cols_10_4_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_410_io_deq_ready = cols_10_5_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_411_clock = clock;
  assign q_411_reset = reset;
  assign q_411_io_enq_valid = cols_10_5_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_411_io_enq_bits = cols_10_5_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_411_io_deq_ready = cols_10_6_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_412_clock = clock;
  assign q_412_reset = reset;
  assign q_412_io_enq_valid = cols_10_6_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_412_io_enq_bits = cols_10_6_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_412_io_deq_ready = cols_10_7_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_413_clock = clock;
  assign q_413_reset = reset;
  assign q_413_io_enq_valid = cols_10_7_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_413_io_enq_bits = cols_10_7_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_413_io_deq_ready = cols_10_8_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_414_clock = clock;
  assign q_414_reset = reset;
  assign q_414_io_enq_valid = cols_10_8_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_414_io_enq_bits = cols_10_8_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_414_io_deq_ready = cols_10_9_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_415_clock = clock;
  assign q_415_reset = reset;
  assign q_415_io_enq_valid = cols_10_9_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_415_io_enq_bits = cols_10_9_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_415_io_deq_ready = cols_10_10_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_416_clock = clock;
  assign q_416_reset = reset;
  assign q_416_io_enq_valid = cols_10_10_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_416_io_enq_bits = cols_10_10_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_416_io_deq_ready = cols_10_11_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_417_clock = clock;
  assign q_417_reset = reset;
  assign q_417_io_enq_valid = cols_10_11_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_417_io_enq_bits = cols_10_11_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_417_io_deq_ready = cols_10_12_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_418_clock = clock;
  assign q_418_reset = reset;
  assign q_418_io_enq_valid = cols_10_12_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_418_io_enq_bits = cols_10_12_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_418_io_deq_ready = cols_10_13_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_419_clock = clock;
  assign q_419_reset = reset;
  assign q_419_io_enq_valid = cols_10_13_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_419_io_enq_bits = cols_10_13_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_419_io_deq_ready = cols_10_14_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_420_clock = clock;
  assign q_420_reset = reset;
  assign q_420_io_enq_valid = cols_10_14_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_420_io_enq_bits = cols_10_14_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_420_io_deq_ready = cols_10_15_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_421_clock = clock;
  assign q_421_reset = reset;
  assign q_421_io_enq_valid = cols_11_0_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_421_io_enq_bits = cols_11_0_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_421_io_deq_ready = cols_11_1_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_422_clock = clock;
  assign q_422_reset = reset;
  assign q_422_io_enq_valid = cols_11_1_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_422_io_enq_bits = cols_11_1_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_422_io_deq_ready = cols_11_2_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_423_clock = clock;
  assign q_423_reset = reset;
  assign q_423_io_enq_valid = cols_11_2_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_423_io_enq_bits = cols_11_2_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_423_io_deq_ready = cols_11_3_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_424_clock = clock;
  assign q_424_reset = reset;
  assign q_424_io_enq_valid = cols_11_3_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_424_io_enq_bits = cols_11_3_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_424_io_deq_ready = cols_11_4_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_425_clock = clock;
  assign q_425_reset = reset;
  assign q_425_io_enq_valid = cols_11_4_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_425_io_enq_bits = cols_11_4_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_425_io_deq_ready = cols_11_5_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_426_clock = clock;
  assign q_426_reset = reset;
  assign q_426_io_enq_valid = cols_11_5_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_426_io_enq_bits = cols_11_5_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_426_io_deq_ready = cols_11_6_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_427_clock = clock;
  assign q_427_reset = reset;
  assign q_427_io_enq_valid = cols_11_6_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_427_io_enq_bits = cols_11_6_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_427_io_deq_ready = cols_11_7_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_428_clock = clock;
  assign q_428_reset = reset;
  assign q_428_io_enq_valid = cols_11_7_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_428_io_enq_bits = cols_11_7_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_428_io_deq_ready = cols_11_8_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_429_clock = clock;
  assign q_429_reset = reset;
  assign q_429_io_enq_valid = cols_11_8_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_429_io_enq_bits = cols_11_8_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_429_io_deq_ready = cols_11_9_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_430_clock = clock;
  assign q_430_reset = reset;
  assign q_430_io_enq_valid = cols_11_9_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_430_io_enq_bits = cols_11_9_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_430_io_deq_ready = cols_11_10_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_431_clock = clock;
  assign q_431_reset = reset;
  assign q_431_io_enq_valid = cols_11_10_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_431_io_enq_bits = cols_11_10_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_431_io_deq_ready = cols_11_11_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_432_clock = clock;
  assign q_432_reset = reset;
  assign q_432_io_enq_valid = cols_11_11_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_432_io_enq_bits = cols_11_11_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_432_io_deq_ready = cols_11_12_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_433_clock = clock;
  assign q_433_reset = reset;
  assign q_433_io_enq_valid = cols_11_12_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_433_io_enq_bits = cols_11_12_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_433_io_deq_ready = cols_11_13_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_434_clock = clock;
  assign q_434_reset = reset;
  assign q_434_io_enq_valid = cols_11_13_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_434_io_enq_bits = cols_11_13_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_434_io_deq_ready = cols_11_14_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_435_clock = clock;
  assign q_435_reset = reset;
  assign q_435_io_enq_valid = cols_11_14_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_435_io_enq_bits = cols_11_14_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_435_io_deq_ready = cols_11_15_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_436_clock = clock;
  assign q_436_reset = reset;
  assign q_436_io_enq_valid = cols_12_0_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_436_io_enq_bits = cols_12_0_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_436_io_deq_ready = cols_12_1_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_437_clock = clock;
  assign q_437_reset = reset;
  assign q_437_io_enq_valid = cols_12_1_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_437_io_enq_bits = cols_12_1_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_437_io_deq_ready = cols_12_2_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_438_clock = clock;
  assign q_438_reset = reset;
  assign q_438_io_enq_valid = cols_12_2_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_438_io_enq_bits = cols_12_2_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_438_io_deq_ready = cols_12_3_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_439_clock = clock;
  assign q_439_reset = reset;
  assign q_439_io_enq_valid = cols_12_3_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_439_io_enq_bits = cols_12_3_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_439_io_deq_ready = cols_12_4_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_440_clock = clock;
  assign q_440_reset = reset;
  assign q_440_io_enq_valid = cols_12_4_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_440_io_enq_bits = cols_12_4_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_440_io_deq_ready = cols_12_5_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_441_clock = clock;
  assign q_441_reset = reset;
  assign q_441_io_enq_valid = cols_12_5_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_441_io_enq_bits = cols_12_5_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_441_io_deq_ready = cols_12_6_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_442_clock = clock;
  assign q_442_reset = reset;
  assign q_442_io_enq_valid = cols_12_6_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_442_io_enq_bits = cols_12_6_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_442_io_deq_ready = cols_12_7_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_443_clock = clock;
  assign q_443_reset = reset;
  assign q_443_io_enq_valid = cols_12_7_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_443_io_enq_bits = cols_12_7_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_443_io_deq_ready = cols_12_8_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_444_clock = clock;
  assign q_444_reset = reset;
  assign q_444_io_enq_valid = cols_12_8_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_444_io_enq_bits = cols_12_8_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_444_io_deq_ready = cols_12_9_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_445_clock = clock;
  assign q_445_reset = reset;
  assign q_445_io_enq_valid = cols_12_9_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_445_io_enq_bits = cols_12_9_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_445_io_deq_ready = cols_12_10_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_446_clock = clock;
  assign q_446_reset = reset;
  assign q_446_io_enq_valid = cols_12_10_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_446_io_enq_bits = cols_12_10_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_446_io_deq_ready = cols_12_11_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_447_clock = clock;
  assign q_447_reset = reset;
  assign q_447_io_enq_valid = cols_12_11_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_447_io_enq_bits = cols_12_11_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_447_io_deq_ready = cols_12_12_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_448_clock = clock;
  assign q_448_reset = reset;
  assign q_448_io_enq_valid = cols_12_12_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_448_io_enq_bits = cols_12_12_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_448_io_deq_ready = cols_12_13_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_449_clock = clock;
  assign q_449_reset = reset;
  assign q_449_io_enq_valid = cols_12_13_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_449_io_enq_bits = cols_12_13_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_449_io_deq_ready = cols_12_14_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_450_clock = clock;
  assign q_450_reset = reset;
  assign q_450_io_enq_valid = cols_12_14_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_450_io_enq_bits = cols_12_14_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_450_io_deq_ready = cols_12_15_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_451_clock = clock;
  assign q_451_reset = reset;
  assign q_451_io_enq_valid = cols_13_0_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_451_io_enq_bits = cols_13_0_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_451_io_deq_ready = cols_13_1_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_452_clock = clock;
  assign q_452_reset = reset;
  assign q_452_io_enq_valid = cols_13_1_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_452_io_enq_bits = cols_13_1_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_452_io_deq_ready = cols_13_2_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_453_clock = clock;
  assign q_453_reset = reset;
  assign q_453_io_enq_valid = cols_13_2_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_453_io_enq_bits = cols_13_2_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_453_io_deq_ready = cols_13_3_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_454_clock = clock;
  assign q_454_reset = reset;
  assign q_454_io_enq_valid = cols_13_3_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_454_io_enq_bits = cols_13_3_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_454_io_deq_ready = cols_13_4_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_455_clock = clock;
  assign q_455_reset = reset;
  assign q_455_io_enq_valid = cols_13_4_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_455_io_enq_bits = cols_13_4_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_455_io_deq_ready = cols_13_5_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_456_clock = clock;
  assign q_456_reset = reset;
  assign q_456_io_enq_valid = cols_13_5_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_456_io_enq_bits = cols_13_5_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_456_io_deq_ready = cols_13_6_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_457_clock = clock;
  assign q_457_reset = reset;
  assign q_457_io_enq_valid = cols_13_6_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_457_io_enq_bits = cols_13_6_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_457_io_deq_ready = cols_13_7_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_458_clock = clock;
  assign q_458_reset = reset;
  assign q_458_io_enq_valid = cols_13_7_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_458_io_enq_bits = cols_13_7_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_458_io_deq_ready = cols_13_8_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_459_clock = clock;
  assign q_459_reset = reset;
  assign q_459_io_enq_valid = cols_13_8_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_459_io_enq_bits = cols_13_8_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_459_io_deq_ready = cols_13_9_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_460_clock = clock;
  assign q_460_reset = reset;
  assign q_460_io_enq_valid = cols_13_9_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_460_io_enq_bits = cols_13_9_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_460_io_deq_ready = cols_13_10_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_461_clock = clock;
  assign q_461_reset = reset;
  assign q_461_io_enq_valid = cols_13_10_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_461_io_enq_bits = cols_13_10_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_461_io_deq_ready = cols_13_11_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_462_clock = clock;
  assign q_462_reset = reset;
  assign q_462_io_enq_valid = cols_13_11_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_462_io_enq_bits = cols_13_11_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_462_io_deq_ready = cols_13_12_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_463_clock = clock;
  assign q_463_reset = reset;
  assign q_463_io_enq_valid = cols_13_12_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_463_io_enq_bits = cols_13_12_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_463_io_deq_ready = cols_13_13_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_464_clock = clock;
  assign q_464_reset = reset;
  assign q_464_io_enq_valid = cols_13_13_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_464_io_enq_bits = cols_13_13_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_464_io_deq_ready = cols_13_14_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_465_clock = clock;
  assign q_465_reset = reset;
  assign q_465_io_enq_valid = cols_13_14_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_465_io_enq_bits = cols_13_14_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_465_io_deq_ready = cols_13_15_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_466_clock = clock;
  assign q_466_reset = reset;
  assign q_466_io_enq_valid = cols_14_0_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_466_io_enq_bits = cols_14_0_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_466_io_deq_ready = cols_14_1_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_467_clock = clock;
  assign q_467_reset = reset;
  assign q_467_io_enq_valid = cols_14_1_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_467_io_enq_bits = cols_14_1_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_467_io_deq_ready = cols_14_2_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_468_clock = clock;
  assign q_468_reset = reset;
  assign q_468_io_enq_valid = cols_14_2_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_468_io_enq_bits = cols_14_2_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_468_io_deq_ready = cols_14_3_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_469_clock = clock;
  assign q_469_reset = reset;
  assign q_469_io_enq_valid = cols_14_3_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_469_io_enq_bits = cols_14_3_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_469_io_deq_ready = cols_14_4_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_470_clock = clock;
  assign q_470_reset = reset;
  assign q_470_io_enq_valid = cols_14_4_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_470_io_enq_bits = cols_14_4_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_470_io_deq_ready = cols_14_5_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_471_clock = clock;
  assign q_471_reset = reset;
  assign q_471_io_enq_valid = cols_14_5_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_471_io_enq_bits = cols_14_5_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_471_io_deq_ready = cols_14_6_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_472_clock = clock;
  assign q_472_reset = reset;
  assign q_472_io_enq_valid = cols_14_6_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_472_io_enq_bits = cols_14_6_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_472_io_deq_ready = cols_14_7_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_473_clock = clock;
  assign q_473_reset = reset;
  assign q_473_io_enq_valid = cols_14_7_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_473_io_enq_bits = cols_14_7_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_473_io_deq_ready = cols_14_8_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_474_clock = clock;
  assign q_474_reset = reset;
  assign q_474_io_enq_valid = cols_14_8_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_474_io_enq_bits = cols_14_8_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_474_io_deq_ready = cols_14_9_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_475_clock = clock;
  assign q_475_reset = reset;
  assign q_475_io_enq_valid = cols_14_9_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_475_io_enq_bits = cols_14_9_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_475_io_deq_ready = cols_14_10_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_476_clock = clock;
  assign q_476_reset = reset;
  assign q_476_io_enq_valid = cols_14_10_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_476_io_enq_bits = cols_14_10_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_476_io_deq_ready = cols_14_11_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_477_clock = clock;
  assign q_477_reset = reset;
  assign q_477_io_enq_valid = cols_14_11_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_477_io_enq_bits = cols_14_11_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_477_io_deq_ready = cols_14_12_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_478_clock = clock;
  assign q_478_reset = reset;
  assign q_478_io_enq_valid = cols_14_12_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_478_io_enq_bits = cols_14_12_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_478_io_deq_ready = cols_14_13_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_479_clock = clock;
  assign q_479_reset = reset;
  assign q_479_io_enq_valid = cols_14_13_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_479_io_enq_bits = cols_14_13_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_479_io_deq_ready = cols_14_14_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_480_clock = clock;
  assign q_480_reset = reset;
  assign q_480_io_enq_valid = cols_14_14_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_480_io_enq_bits = cols_14_14_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_480_io_deq_ready = cols_14_15_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_481_clock = clock;
  assign q_481_reset = reset;
  assign q_481_io_enq_valid = cols_15_0_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_481_io_enq_bits = cols_15_0_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_481_io_deq_ready = cols_15_1_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_482_clock = clock;
  assign q_482_reset = reset;
  assign q_482_io_enq_valid = cols_15_1_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_482_io_enq_bits = cols_15_1_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_482_io_deq_ready = cols_15_2_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_483_clock = clock;
  assign q_483_reset = reset;
  assign q_483_io_enq_valid = cols_15_2_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_483_io_enq_bits = cols_15_2_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_483_io_deq_ready = cols_15_3_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_484_clock = clock;
  assign q_484_reset = reset;
  assign q_484_io_enq_valid = cols_15_3_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_484_io_enq_bits = cols_15_3_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_484_io_deq_ready = cols_15_4_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_485_clock = clock;
  assign q_485_reset = reset;
  assign q_485_io_enq_valid = cols_15_4_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_485_io_enq_bits = cols_15_4_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_485_io_deq_ready = cols_15_5_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_486_clock = clock;
  assign q_486_reset = reset;
  assign q_486_io_enq_valid = cols_15_5_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_486_io_enq_bits = cols_15_5_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_486_io_deq_ready = cols_15_6_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_487_clock = clock;
  assign q_487_reset = reset;
  assign q_487_io_enq_valid = cols_15_6_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_487_io_enq_bits = cols_15_6_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_487_io_deq_ready = cols_15_7_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_488_clock = clock;
  assign q_488_reset = reset;
  assign q_488_io_enq_valid = cols_15_7_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_488_io_enq_bits = cols_15_7_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_488_io_deq_ready = cols_15_8_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_489_clock = clock;
  assign q_489_reset = reset;
  assign q_489_io_enq_valid = cols_15_8_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_489_io_enq_bits = cols_15_8_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_489_io_deq_ready = cols_15_9_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_490_clock = clock;
  assign q_490_reset = reset;
  assign q_490_io_enq_valid = cols_15_9_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_490_io_enq_bits = cols_15_9_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_490_io_deq_ready = cols_15_10_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_491_clock = clock;
  assign q_491_reset = reset;
  assign q_491_io_enq_valid = cols_15_10_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_491_io_enq_bits = cols_15_10_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_491_io_deq_ready = cols_15_11_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_492_clock = clock;
  assign q_492_reset = reset;
  assign q_492_io_enq_valid = cols_15_11_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_492_io_enq_bits = cols_15_11_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_492_io_deq_ready = cols_15_12_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_493_clock = clock;
  assign q_493_reset = reset;
  assign q_493_io_enq_valid = cols_15_12_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_493_io_enq_bits = cols_15_12_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_493_io_deq_ready = cols_15_13_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_494_clock = clock;
  assign q_494_reset = reset;
  assign q_494_io_enq_valid = cols_15_13_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_494_io_enq_bits = cols_15_13_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_494_io_deq_ready = cols_15_14_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_495_clock = clock;
  assign q_495_reset = reset;
  assign q_495_io_enq_valid = cols_15_14_io_bottom_out_valid; // @[Decoupled.scala 363:22]
  assign q_495_io_enq_bits = cols_15_14_io_bottom_out_bits; // @[Decoupled.scala 364:21]
  assign q_495_io_deq_ready = cols_15_15_io_top_in_ready; // @[Stab.scala 97:70]
  assign q_496_clock = clock;
  assign q_496_reset = reset;
  assign q_496_io_enq_valid = io_value_in_0_valid; // @[Decoupled.scala 363:22]
  assign q_496_io_enq_bits = io_value_in_0_bits; // @[Decoupled.scala 364:21]
  assign q_496_io_deq_ready = cols_0_0_io_left_in_ready; // @[Stab.scala 100:101]
  assign q_497_clock = clock;
  assign q_497_reset = reset;
  assign q_497_io_enq_valid = io_value_in_1_valid; // @[Decoupled.scala 363:22]
  assign q_497_io_enq_bits = io_value_in_1_bits; // @[Decoupled.scala 364:21]
  assign q_497_io_deq_ready = cols_0_1_io_left_in_ready; // @[Stab.scala 100:101]
  assign q_498_clock = clock;
  assign q_498_reset = reset;
  assign q_498_io_enq_valid = io_value_in_2_valid; // @[Decoupled.scala 363:22]
  assign q_498_io_enq_bits = io_value_in_2_bits; // @[Decoupled.scala 364:21]
  assign q_498_io_deq_ready = cols_0_2_io_left_in_ready; // @[Stab.scala 100:101]
  assign q_499_clock = clock;
  assign q_499_reset = reset;
  assign q_499_io_enq_valid = io_value_in_3_valid; // @[Decoupled.scala 363:22]
  assign q_499_io_enq_bits = io_value_in_3_bits; // @[Decoupled.scala 364:21]
  assign q_499_io_deq_ready = cols_0_3_io_left_in_ready; // @[Stab.scala 100:101]
  assign q_500_clock = clock;
  assign q_500_reset = reset;
  assign q_500_io_enq_valid = io_value_in_4_valid; // @[Decoupled.scala 363:22]
  assign q_500_io_enq_bits = io_value_in_4_bits; // @[Decoupled.scala 364:21]
  assign q_500_io_deq_ready = cols_0_4_io_left_in_ready; // @[Stab.scala 100:101]
  assign q_501_clock = clock;
  assign q_501_reset = reset;
  assign q_501_io_enq_valid = io_value_in_5_valid; // @[Decoupled.scala 363:22]
  assign q_501_io_enq_bits = io_value_in_5_bits; // @[Decoupled.scala 364:21]
  assign q_501_io_deq_ready = cols_0_5_io_left_in_ready; // @[Stab.scala 100:101]
  assign q_502_clock = clock;
  assign q_502_reset = reset;
  assign q_502_io_enq_valid = io_value_in_6_valid; // @[Decoupled.scala 363:22]
  assign q_502_io_enq_bits = io_value_in_6_bits; // @[Decoupled.scala 364:21]
  assign q_502_io_deq_ready = cols_0_6_io_left_in_ready; // @[Stab.scala 100:101]
  assign q_503_clock = clock;
  assign q_503_reset = reset;
  assign q_503_io_enq_valid = io_value_in_7_valid; // @[Decoupled.scala 363:22]
  assign q_503_io_enq_bits = io_value_in_7_bits; // @[Decoupled.scala 364:21]
  assign q_503_io_deq_ready = cols_0_7_io_left_in_ready; // @[Stab.scala 100:101]
  assign q_504_clock = clock;
  assign q_504_reset = reset;
  assign q_504_io_enq_valid = io_value_in_8_valid; // @[Decoupled.scala 363:22]
  assign q_504_io_enq_bits = io_value_in_8_bits; // @[Decoupled.scala 364:21]
  assign q_504_io_deq_ready = cols_0_8_io_left_in_ready; // @[Stab.scala 100:101]
  assign q_505_clock = clock;
  assign q_505_reset = reset;
  assign q_505_io_enq_valid = io_value_in_9_valid; // @[Decoupled.scala 363:22]
  assign q_505_io_enq_bits = io_value_in_9_bits; // @[Decoupled.scala 364:21]
  assign q_505_io_deq_ready = cols_0_9_io_left_in_ready; // @[Stab.scala 100:101]
  assign q_506_clock = clock;
  assign q_506_reset = reset;
  assign q_506_io_enq_valid = io_value_in_10_valid; // @[Decoupled.scala 363:22]
  assign q_506_io_enq_bits = io_value_in_10_bits; // @[Decoupled.scala 364:21]
  assign q_506_io_deq_ready = cols_0_10_io_left_in_ready; // @[Stab.scala 100:101]
  assign q_507_clock = clock;
  assign q_507_reset = reset;
  assign q_507_io_enq_valid = io_value_in_11_valid; // @[Decoupled.scala 363:22]
  assign q_507_io_enq_bits = io_value_in_11_bits; // @[Decoupled.scala 364:21]
  assign q_507_io_deq_ready = cols_0_11_io_left_in_ready; // @[Stab.scala 100:101]
  assign q_508_clock = clock;
  assign q_508_reset = reset;
  assign q_508_io_enq_valid = io_value_in_12_valid; // @[Decoupled.scala 363:22]
  assign q_508_io_enq_bits = io_value_in_12_bits; // @[Decoupled.scala 364:21]
  assign q_508_io_deq_ready = cols_0_12_io_left_in_ready; // @[Stab.scala 100:101]
  assign q_509_clock = clock;
  assign q_509_reset = reset;
  assign q_509_io_enq_valid = io_value_in_13_valid; // @[Decoupled.scala 363:22]
  assign q_509_io_enq_bits = io_value_in_13_bits; // @[Decoupled.scala 364:21]
  assign q_509_io_deq_ready = cols_0_13_io_left_in_ready; // @[Stab.scala 100:101]
  assign q_510_clock = clock;
  assign q_510_reset = reset;
  assign q_510_io_enq_valid = io_value_in_14_valid; // @[Decoupled.scala 363:22]
  assign q_510_io_enq_bits = io_value_in_14_bits; // @[Decoupled.scala 364:21]
  assign q_510_io_deq_ready = cols_0_14_io_left_in_ready; // @[Stab.scala 100:101]
  assign q_511_clock = clock;
  assign q_511_reset = reset;
  assign q_511_io_enq_valid = io_value_in_15_valid; // @[Decoupled.scala 363:22]
  assign q_511_io_enq_bits = io_value_in_15_bits; // @[Decoupled.scala 364:21]
  assign q_511_io_deq_ready = cols_0_15_io_left_in_ready; // @[Stab.scala 100:101]
  assign q_512_clock = clock;
  assign q_512_reset = reset;
  assign q_512_io_enq_valid = cols_0_0_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_512_io_enq_bits = cols_0_0_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_512_io_deq_ready = io_value_out_0_0_ready; // @[Stab.scala 104:101]
  assign q_513_clock = clock;
  assign q_513_reset = reset;
  assign q_513_io_enq_valid = cols_1_0_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_513_io_enq_bits = cols_1_0_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_513_io_deq_ready = io_value_out_0_1_ready; // @[Stab.scala 104:101]
  assign q_514_clock = clock;
  assign q_514_reset = reset;
  assign q_514_io_enq_valid = cols_2_0_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_514_io_enq_bits = cols_2_0_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_514_io_deq_ready = io_value_out_0_2_ready; // @[Stab.scala 104:101]
  assign q_515_clock = clock;
  assign q_515_reset = reset;
  assign q_515_io_enq_valid = cols_3_0_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_515_io_enq_bits = cols_3_0_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_515_io_deq_ready = io_value_out_0_3_ready; // @[Stab.scala 104:101]
  assign q_516_clock = clock;
  assign q_516_reset = reset;
  assign q_516_io_enq_valid = cols_4_0_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_516_io_enq_bits = cols_4_0_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_516_io_deq_ready = io_value_out_0_4_ready; // @[Stab.scala 104:101]
  assign q_517_clock = clock;
  assign q_517_reset = reset;
  assign q_517_io_enq_valid = cols_5_0_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_517_io_enq_bits = cols_5_0_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_517_io_deq_ready = io_value_out_0_5_ready; // @[Stab.scala 104:101]
  assign q_518_clock = clock;
  assign q_518_reset = reset;
  assign q_518_io_enq_valid = cols_6_0_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_518_io_enq_bits = cols_6_0_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_518_io_deq_ready = io_value_out_0_6_ready; // @[Stab.scala 104:101]
  assign q_519_clock = clock;
  assign q_519_reset = reset;
  assign q_519_io_enq_valid = cols_7_0_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_519_io_enq_bits = cols_7_0_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_519_io_deq_ready = io_value_out_0_7_ready; // @[Stab.scala 104:101]
  assign q_520_clock = clock;
  assign q_520_reset = reset;
  assign q_520_io_enq_valid = cols_8_0_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_520_io_enq_bits = cols_8_0_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_520_io_deq_ready = io_value_out_0_8_ready; // @[Stab.scala 104:101]
  assign q_521_clock = clock;
  assign q_521_reset = reset;
  assign q_521_io_enq_valid = cols_9_0_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_521_io_enq_bits = cols_9_0_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_521_io_deq_ready = io_value_out_0_9_ready; // @[Stab.scala 104:101]
  assign q_522_clock = clock;
  assign q_522_reset = reset;
  assign q_522_io_enq_valid = cols_10_0_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_522_io_enq_bits = cols_10_0_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_522_io_deq_ready = io_value_out_0_10_ready; // @[Stab.scala 104:101]
  assign q_523_clock = clock;
  assign q_523_reset = reset;
  assign q_523_io_enq_valid = cols_11_0_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_523_io_enq_bits = cols_11_0_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_523_io_deq_ready = io_value_out_0_11_ready; // @[Stab.scala 104:101]
  assign q_524_clock = clock;
  assign q_524_reset = reset;
  assign q_524_io_enq_valid = cols_12_0_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_524_io_enq_bits = cols_12_0_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_524_io_deq_ready = io_value_out_0_12_ready; // @[Stab.scala 104:101]
  assign q_525_clock = clock;
  assign q_525_reset = reset;
  assign q_525_io_enq_valid = cols_13_0_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_525_io_enq_bits = cols_13_0_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_525_io_deq_ready = io_value_out_0_13_ready; // @[Stab.scala 104:101]
  assign q_526_clock = clock;
  assign q_526_reset = reset;
  assign q_526_io_enq_valid = cols_14_0_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_526_io_enq_bits = cols_14_0_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_526_io_deq_ready = io_value_out_0_14_ready; // @[Stab.scala 104:101]
  assign q_527_clock = clock;
  assign q_527_reset = reset;
  assign q_527_io_enq_valid = cols_15_0_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_527_io_enq_bits = cols_15_0_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_527_io_deq_ready = io_value_out_0_15_ready; // @[Stab.scala 104:101]
  assign q_528_clock = clock;
  assign q_528_reset = reset;
  assign q_528_io_enq_valid = cols_0_1_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_528_io_enq_bits = cols_0_1_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_528_io_deq_ready = io_value_out_1_0_ready; // @[Stab.scala 104:101]
  assign q_529_clock = clock;
  assign q_529_reset = reset;
  assign q_529_io_enq_valid = cols_1_1_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_529_io_enq_bits = cols_1_1_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_529_io_deq_ready = io_value_out_1_1_ready; // @[Stab.scala 104:101]
  assign q_530_clock = clock;
  assign q_530_reset = reset;
  assign q_530_io_enq_valid = cols_2_1_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_530_io_enq_bits = cols_2_1_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_530_io_deq_ready = io_value_out_1_2_ready; // @[Stab.scala 104:101]
  assign q_531_clock = clock;
  assign q_531_reset = reset;
  assign q_531_io_enq_valid = cols_3_1_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_531_io_enq_bits = cols_3_1_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_531_io_deq_ready = io_value_out_1_3_ready; // @[Stab.scala 104:101]
  assign q_532_clock = clock;
  assign q_532_reset = reset;
  assign q_532_io_enq_valid = cols_4_1_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_532_io_enq_bits = cols_4_1_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_532_io_deq_ready = io_value_out_1_4_ready; // @[Stab.scala 104:101]
  assign q_533_clock = clock;
  assign q_533_reset = reset;
  assign q_533_io_enq_valid = cols_5_1_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_533_io_enq_bits = cols_5_1_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_533_io_deq_ready = io_value_out_1_5_ready; // @[Stab.scala 104:101]
  assign q_534_clock = clock;
  assign q_534_reset = reset;
  assign q_534_io_enq_valid = cols_6_1_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_534_io_enq_bits = cols_6_1_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_534_io_deq_ready = io_value_out_1_6_ready; // @[Stab.scala 104:101]
  assign q_535_clock = clock;
  assign q_535_reset = reset;
  assign q_535_io_enq_valid = cols_7_1_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_535_io_enq_bits = cols_7_1_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_535_io_deq_ready = io_value_out_1_7_ready; // @[Stab.scala 104:101]
  assign q_536_clock = clock;
  assign q_536_reset = reset;
  assign q_536_io_enq_valid = cols_8_1_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_536_io_enq_bits = cols_8_1_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_536_io_deq_ready = io_value_out_1_8_ready; // @[Stab.scala 104:101]
  assign q_537_clock = clock;
  assign q_537_reset = reset;
  assign q_537_io_enq_valid = cols_9_1_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_537_io_enq_bits = cols_9_1_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_537_io_deq_ready = io_value_out_1_9_ready; // @[Stab.scala 104:101]
  assign q_538_clock = clock;
  assign q_538_reset = reset;
  assign q_538_io_enq_valid = cols_10_1_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_538_io_enq_bits = cols_10_1_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_538_io_deq_ready = io_value_out_1_10_ready; // @[Stab.scala 104:101]
  assign q_539_clock = clock;
  assign q_539_reset = reset;
  assign q_539_io_enq_valid = cols_11_1_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_539_io_enq_bits = cols_11_1_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_539_io_deq_ready = io_value_out_1_11_ready; // @[Stab.scala 104:101]
  assign q_540_clock = clock;
  assign q_540_reset = reset;
  assign q_540_io_enq_valid = cols_12_1_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_540_io_enq_bits = cols_12_1_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_540_io_deq_ready = io_value_out_1_12_ready; // @[Stab.scala 104:101]
  assign q_541_clock = clock;
  assign q_541_reset = reset;
  assign q_541_io_enq_valid = cols_13_1_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_541_io_enq_bits = cols_13_1_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_541_io_deq_ready = io_value_out_1_13_ready; // @[Stab.scala 104:101]
  assign q_542_clock = clock;
  assign q_542_reset = reset;
  assign q_542_io_enq_valid = cols_14_1_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_542_io_enq_bits = cols_14_1_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_542_io_deq_ready = io_value_out_1_14_ready; // @[Stab.scala 104:101]
  assign q_543_clock = clock;
  assign q_543_reset = reset;
  assign q_543_io_enq_valid = cols_15_1_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_543_io_enq_bits = cols_15_1_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_543_io_deq_ready = io_value_out_1_15_ready; // @[Stab.scala 104:101]
  assign q_544_clock = clock;
  assign q_544_reset = reset;
  assign q_544_io_enq_valid = cols_0_2_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_544_io_enq_bits = cols_0_2_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_544_io_deq_ready = io_value_out_2_0_ready; // @[Stab.scala 104:101]
  assign q_545_clock = clock;
  assign q_545_reset = reset;
  assign q_545_io_enq_valid = cols_1_2_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_545_io_enq_bits = cols_1_2_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_545_io_deq_ready = io_value_out_2_1_ready; // @[Stab.scala 104:101]
  assign q_546_clock = clock;
  assign q_546_reset = reset;
  assign q_546_io_enq_valid = cols_2_2_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_546_io_enq_bits = cols_2_2_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_546_io_deq_ready = io_value_out_2_2_ready; // @[Stab.scala 104:101]
  assign q_547_clock = clock;
  assign q_547_reset = reset;
  assign q_547_io_enq_valid = cols_3_2_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_547_io_enq_bits = cols_3_2_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_547_io_deq_ready = io_value_out_2_3_ready; // @[Stab.scala 104:101]
  assign q_548_clock = clock;
  assign q_548_reset = reset;
  assign q_548_io_enq_valid = cols_4_2_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_548_io_enq_bits = cols_4_2_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_548_io_deq_ready = io_value_out_2_4_ready; // @[Stab.scala 104:101]
  assign q_549_clock = clock;
  assign q_549_reset = reset;
  assign q_549_io_enq_valid = cols_5_2_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_549_io_enq_bits = cols_5_2_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_549_io_deq_ready = io_value_out_2_5_ready; // @[Stab.scala 104:101]
  assign q_550_clock = clock;
  assign q_550_reset = reset;
  assign q_550_io_enq_valid = cols_6_2_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_550_io_enq_bits = cols_6_2_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_550_io_deq_ready = io_value_out_2_6_ready; // @[Stab.scala 104:101]
  assign q_551_clock = clock;
  assign q_551_reset = reset;
  assign q_551_io_enq_valid = cols_7_2_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_551_io_enq_bits = cols_7_2_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_551_io_deq_ready = io_value_out_2_7_ready; // @[Stab.scala 104:101]
  assign q_552_clock = clock;
  assign q_552_reset = reset;
  assign q_552_io_enq_valid = cols_8_2_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_552_io_enq_bits = cols_8_2_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_552_io_deq_ready = io_value_out_2_8_ready; // @[Stab.scala 104:101]
  assign q_553_clock = clock;
  assign q_553_reset = reset;
  assign q_553_io_enq_valid = cols_9_2_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_553_io_enq_bits = cols_9_2_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_553_io_deq_ready = io_value_out_2_9_ready; // @[Stab.scala 104:101]
  assign q_554_clock = clock;
  assign q_554_reset = reset;
  assign q_554_io_enq_valid = cols_10_2_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_554_io_enq_bits = cols_10_2_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_554_io_deq_ready = io_value_out_2_10_ready; // @[Stab.scala 104:101]
  assign q_555_clock = clock;
  assign q_555_reset = reset;
  assign q_555_io_enq_valid = cols_11_2_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_555_io_enq_bits = cols_11_2_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_555_io_deq_ready = io_value_out_2_11_ready; // @[Stab.scala 104:101]
  assign q_556_clock = clock;
  assign q_556_reset = reset;
  assign q_556_io_enq_valid = cols_12_2_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_556_io_enq_bits = cols_12_2_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_556_io_deq_ready = io_value_out_2_12_ready; // @[Stab.scala 104:101]
  assign q_557_clock = clock;
  assign q_557_reset = reset;
  assign q_557_io_enq_valid = cols_13_2_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_557_io_enq_bits = cols_13_2_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_557_io_deq_ready = io_value_out_2_13_ready; // @[Stab.scala 104:101]
  assign q_558_clock = clock;
  assign q_558_reset = reset;
  assign q_558_io_enq_valid = cols_14_2_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_558_io_enq_bits = cols_14_2_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_558_io_deq_ready = io_value_out_2_14_ready; // @[Stab.scala 104:101]
  assign q_559_clock = clock;
  assign q_559_reset = reset;
  assign q_559_io_enq_valid = cols_15_2_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_559_io_enq_bits = cols_15_2_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_559_io_deq_ready = io_value_out_2_15_ready; // @[Stab.scala 104:101]
  assign q_560_clock = clock;
  assign q_560_reset = reset;
  assign q_560_io_enq_valid = cols_0_3_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_560_io_enq_bits = cols_0_3_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_560_io_deq_ready = io_value_out_3_0_ready; // @[Stab.scala 104:101]
  assign q_561_clock = clock;
  assign q_561_reset = reset;
  assign q_561_io_enq_valid = cols_1_3_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_561_io_enq_bits = cols_1_3_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_561_io_deq_ready = io_value_out_3_1_ready; // @[Stab.scala 104:101]
  assign q_562_clock = clock;
  assign q_562_reset = reset;
  assign q_562_io_enq_valid = cols_2_3_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_562_io_enq_bits = cols_2_3_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_562_io_deq_ready = io_value_out_3_2_ready; // @[Stab.scala 104:101]
  assign q_563_clock = clock;
  assign q_563_reset = reset;
  assign q_563_io_enq_valid = cols_3_3_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_563_io_enq_bits = cols_3_3_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_563_io_deq_ready = io_value_out_3_3_ready; // @[Stab.scala 104:101]
  assign q_564_clock = clock;
  assign q_564_reset = reset;
  assign q_564_io_enq_valid = cols_4_3_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_564_io_enq_bits = cols_4_3_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_564_io_deq_ready = io_value_out_3_4_ready; // @[Stab.scala 104:101]
  assign q_565_clock = clock;
  assign q_565_reset = reset;
  assign q_565_io_enq_valid = cols_5_3_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_565_io_enq_bits = cols_5_3_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_565_io_deq_ready = io_value_out_3_5_ready; // @[Stab.scala 104:101]
  assign q_566_clock = clock;
  assign q_566_reset = reset;
  assign q_566_io_enq_valid = cols_6_3_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_566_io_enq_bits = cols_6_3_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_566_io_deq_ready = io_value_out_3_6_ready; // @[Stab.scala 104:101]
  assign q_567_clock = clock;
  assign q_567_reset = reset;
  assign q_567_io_enq_valid = cols_7_3_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_567_io_enq_bits = cols_7_3_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_567_io_deq_ready = io_value_out_3_7_ready; // @[Stab.scala 104:101]
  assign q_568_clock = clock;
  assign q_568_reset = reset;
  assign q_568_io_enq_valid = cols_8_3_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_568_io_enq_bits = cols_8_3_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_568_io_deq_ready = io_value_out_3_8_ready; // @[Stab.scala 104:101]
  assign q_569_clock = clock;
  assign q_569_reset = reset;
  assign q_569_io_enq_valid = cols_9_3_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_569_io_enq_bits = cols_9_3_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_569_io_deq_ready = io_value_out_3_9_ready; // @[Stab.scala 104:101]
  assign q_570_clock = clock;
  assign q_570_reset = reset;
  assign q_570_io_enq_valid = cols_10_3_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_570_io_enq_bits = cols_10_3_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_570_io_deq_ready = io_value_out_3_10_ready; // @[Stab.scala 104:101]
  assign q_571_clock = clock;
  assign q_571_reset = reset;
  assign q_571_io_enq_valid = cols_11_3_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_571_io_enq_bits = cols_11_3_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_571_io_deq_ready = io_value_out_3_11_ready; // @[Stab.scala 104:101]
  assign q_572_clock = clock;
  assign q_572_reset = reset;
  assign q_572_io_enq_valid = cols_12_3_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_572_io_enq_bits = cols_12_3_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_572_io_deq_ready = io_value_out_3_12_ready; // @[Stab.scala 104:101]
  assign q_573_clock = clock;
  assign q_573_reset = reset;
  assign q_573_io_enq_valid = cols_13_3_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_573_io_enq_bits = cols_13_3_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_573_io_deq_ready = io_value_out_3_13_ready; // @[Stab.scala 104:101]
  assign q_574_clock = clock;
  assign q_574_reset = reset;
  assign q_574_io_enq_valid = cols_14_3_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_574_io_enq_bits = cols_14_3_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_574_io_deq_ready = io_value_out_3_14_ready; // @[Stab.scala 104:101]
  assign q_575_clock = clock;
  assign q_575_reset = reset;
  assign q_575_io_enq_valid = cols_15_3_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_575_io_enq_bits = cols_15_3_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_575_io_deq_ready = io_value_out_3_15_ready; // @[Stab.scala 104:101]
  assign q_576_clock = clock;
  assign q_576_reset = reset;
  assign q_576_io_enq_valid = cols_0_4_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_576_io_enq_bits = cols_0_4_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_576_io_deq_ready = io_value_out_4_0_ready; // @[Stab.scala 104:101]
  assign q_577_clock = clock;
  assign q_577_reset = reset;
  assign q_577_io_enq_valid = cols_1_4_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_577_io_enq_bits = cols_1_4_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_577_io_deq_ready = io_value_out_4_1_ready; // @[Stab.scala 104:101]
  assign q_578_clock = clock;
  assign q_578_reset = reset;
  assign q_578_io_enq_valid = cols_2_4_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_578_io_enq_bits = cols_2_4_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_578_io_deq_ready = io_value_out_4_2_ready; // @[Stab.scala 104:101]
  assign q_579_clock = clock;
  assign q_579_reset = reset;
  assign q_579_io_enq_valid = cols_3_4_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_579_io_enq_bits = cols_3_4_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_579_io_deq_ready = io_value_out_4_3_ready; // @[Stab.scala 104:101]
  assign q_580_clock = clock;
  assign q_580_reset = reset;
  assign q_580_io_enq_valid = cols_4_4_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_580_io_enq_bits = cols_4_4_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_580_io_deq_ready = io_value_out_4_4_ready; // @[Stab.scala 104:101]
  assign q_581_clock = clock;
  assign q_581_reset = reset;
  assign q_581_io_enq_valid = cols_5_4_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_581_io_enq_bits = cols_5_4_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_581_io_deq_ready = io_value_out_4_5_ready; // @[Stab.scala 104:101]
  assign q_582_clock = clock;
  assign q_582_reset = reset;
  assign q_582_io_enq_valid = cols_6_4_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_582_io_enq_bits = cols_6_4_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_582_io_deq_ready = io_value_out_4_6_ready; // @[Stab.scala 104:101]
  assign q_583_clock = clock;
  assign q_583_reset = reset;
  assign q_583_io_enq_valid = cols_7_4_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_583_io_enq_bits = cols_7_4_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_583_io_deq_ready = io_value_out_4_7_ready; // @[Stab.scala 104:101]
  assign q_584_clock = clock;
  assign q_584_reset = reset;
  assign q_584_io_enq_valid = cols_8_4_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_584_io_enq_bits = cols_8_4_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_584_io_deq_ready = io_value_out_4_8_ready; // @[Stab.scala 104:101]
  assign q_585_clock = clock;
  assign q_585_reset = reset;
  assign q_585_io_enq_valid = cols_9_4_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_585_io_enq_bits = cols_9_4_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_585_io_deq_ready = io_value_out_4_9_ready; // @[Stab.scala 104:101]
  assign q_586_clock = clock;
  assign q_586_reset = reset;
  assign q_586_io_enq_valid = cols_10_4_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_586_io_enq_bits = cols_10_4_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_586_io_deq_ready = io_value_out_4_10_ready; // @[Stab.scala 104:101]
  assign q_587_clock = clock;
  assign q_587_reset = reset;
  assign q_587_io_enq_valid = cols_11_4_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_587_io_enq_bits = cols_11_4_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_587_io_deq_ready = io_value_out_4_11_ready; // @[Stab.scala 104:101]
  assign q_588_clock = clock;
  assign q_588_reset = reset;
  assign q_588_io_enq_valid = cols_12_4_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_588_io_enq_bits = cols_12_4_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_588_io_deq_ready = io_value_out_4_12_ready; // @[Stab.scala 104:101]
  assign q_589_clock = clock;
  assign q_589_reset = reset;
  assign q_589_io_enq_valid = cols_13_4_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_589_io_enq_bits = cols_13_4_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_589_io_deq_ready = io_value_out_4_13_ready; // @[Stab.scala 104:101]
  assign q_590_clock = clock;
  assign q_590_reset = reset;
  assign q_590_io_enq_valid = cols_14_4_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_590_io_enq_bits = cols_14_4_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_590_io_deq_ready = io_value_out_4_14_ready; // @[Stab.scala 104:101]
  assign q_591_clock = clock;
  assign q_591_reset = reset;
  assign q_591_io_enq_valid = cols_15_4_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_591_io_enq_bits = cols_15_4_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_591_io_deq_ready = io_value_out_4_15_ready; // @[Stab.scala 104:101]
  assign q_592_clock = clock;
  assign q_592_reset = reset;
  assign q_592_io_enq_valid = cols_0_5_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_592_io_enq_bits = cols_0_5_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_592_io_deq_ready = io_value_out_5_0_ready; // @[Stab.scala 104:101]
  assign q_593_clock = clock;
  assign q_593_reset = reset;
  assign q_593_io_enq_valid = cols_1_5_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_593_io_enq_bits = cols_1_5_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_593_io_deq_ready = io_value_out_5_1_ready; // @[Stab.scala 104:101]
  assign q_594_clock = clock;
  assign q_594_reset = reset;
  assign q_594_io_enq_valid = cols_2_5_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_594_io_enq_bits = cols_2_5_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_594_io_deq_ready = io_value_out_5_2_ready; // @[Stab.scala 104:101]
  assign q_595_clock = clock;
  assign q_595_reset = reset;
  assign q_595_io_enq_valid = cols_3_5_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_595_io_enq_bits = cols_3_5_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_595_io_deq_ready = io_value_out_5_3_ready; // @[Stab.scala 104:101]
  assign q_596_clock = clock;
  assign q_596_reset = reset;
  assign q_596_io_enq_valid = cols_4_5_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_596_io_enq_bits = cols_4_5_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_596_io_deq_ready = io_value_out_5_4_ready; // @[Stab.scala 104:101]
  assign q_597_clock = clock;
  assign q_597_reset = reset;
  assign q_597_io_enq_valid = cols_5_5_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_597_io_enq_bits = cols_5_5_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_597_io_deq_ready = io_value_out_5_5_ready; // @[Stab.scala 104:101]
  assign q_598_clock = clock;
  assign q_598_reset = reset;
  assign q_598_io_enq_valid = cols_6_5_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_598_io_enq_bits = cols_6_5_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_598_io_deq_ready = io_value_out_5_6_ready; // @[Stab.scala 104:101]
  assign q_599_clock = clock;
  assign q_599_reset = reset;
  assign q_599_io_enq_valid = cols_7_5_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_599_io_enq_bits = cols_7_5_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_599_io_deq_ready = io_value_out_5_7_ready; // @[Stab.scala 104:101]
  assign q_600_clock = clock;
  assign q_600_reset = reset;
  assign q_600_io_enq_valid = cols_8_5_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_600_io_enq_bits = cols_8_5_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_600_io_deq_ready = io_value_out_5_8_ready; // @[Stab.scala 104:101]
  assign q_601_clock = clock;
  assign q_601_reset = reset;
  assign q_601_io_enq_valid = cols_9_5_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_601_io_enq_bits = cols_9_5_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_601_io_deq_ready = io_value_out_5_9_ready; // @[Stab.scala 104:101]
  assign q_602_clock = clock;
  assign q_602_reset = reset;
  assign q_602_io_enq_valid = cols_10_5_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_602_io_enq_bits = cols_10_5_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_602_io_deq_ready = io_value_out_5_10_ready; // @[Stab.scala 104:101]
  assign q_603_clock = clock;
  assign q_603_reset = reset;
  assign q_603_io_enq_valid = cols_11_5_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_603_io_enq_bits = cols_11_5_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_603_io_deq_ready = io_value_out_5_11_ready; // @[Stab.scala 104:101]
  assign q_604_clock = clock;
  assign q_604_reset = reset;
  assign q_604_io_enq_valid = cols_12_5_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_604_io_enq_bits = cols_12_5_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_604_io_deq_ready = io_value_out_5_12_ready; // @[Stab.scala 104:101]
  assign q_605_clock = clock;
  assign q_605_reset = reset;
  assign q_605_io_enq_valid = cols_13_5_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_605_io_enq_bits = cols_13_5_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_605_io_deq_ready = io_value_out_5_13_ready; // @[Stab.scala 104:101]
  assign q_606_clock = clock;
  assign q_606_reset = reset;
  assign q_606_io_enq_valid = cols_14_5_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_606_io_enq_bits = cols_14_5_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_606_io_deq_ready = io_value_out_5_14_ready; // @[Stab.scala 104:101]
  assign q_607_clock = clock;
  assign q_607_reset = reset;
  assign q_607_io_enq_valid = cols_15_5_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_607_io_enq_bits = cols_15_5_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_607_io_deq_ready = io_value_out_5_15_ready; // @[Stab.scala 104:101]
  assign q_608_clock = clock;
  assign q_608_reset = reset;
  assign q_608_io_enq_valid = cols_0_6_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_608_io_enq_bits = cols_0_6_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_608_io_deq_ready = io_value_out_6_0_ready; // @[Stab.scala 104:101]
  assign q_609_clock = clock;
  assign q_609_reset = reset;
  assign q_609_io_enq_valid = cols_1_6_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_609_io_enq_bits = cols_1_6_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_609_io_deq_ready = io_value_out_6_1_ready; // @[Stab.scala 104:101]
  assign q_610_clock = clock;
  assign q_610_reset = reset;
  assign q_610_io_enq_valid = cols_2_6_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_610_io_enq_bits = cols_2_6_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_610_io_deq_ready = io_value_out_6_2_ready; // @[Stab.scala 104:101]
  assign q_611_clock = clock;
  assign q_611_reset = reset;
  assign q_611_io_enq_valid = cols_3_6_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_611_io_enq_bits = cols_3_6_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_611_io_deq_ready = io_value_out_6_3_ready; // @[Stab.scala 104:101]
  assign q_612_clock = clock;
  assign q_612_reset = reset;
  assign q_612_io_enq_valid = cols_4_6_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_612_io_enq_bits = cols_4_6_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_612_io_deq_ready = io_value_out_6_4_ready; // @[Stab.scala 104:101]
  assign q_613_clock = clock;
  assign q_613_reset = reset;
  assign q_613_io_enq_valid = cols_5_6_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_613_io_enq_bits = cols_5_6_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_613_io_deq_ready = io_value_out_6_5_ready; // @[Stab.scala 104:101]
  assign q_614_clock = clock;
  assign q_614_reset = reset;
  assign q_614_io_enq_valid = cols_6_6_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_614_io_enq_bits = cols_6_6_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_614_io_deq_ready = io_value_out_6_6_ready; // @[Stab.scala 104:101]
  assign q_615_clock = clock;
  assign q_615_reset = reset;
  assign q_615_io_enq_valid = cols_7_6_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_615_io_enq_bits = cols_7_6_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_615_io_deq_ready = io_value_out_6_7_ready; // @[Stab.scala 104:101]
  assign q_616_clock = clock;
  assign q_616_reset = reset;
  assign q_616_io_enq_valid = cols_8_6_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_616_io_enq_bits = cols_8_6_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_616_io_deq_ready = io_value_out_6_8_ready; // @[Stab.scala 104:101]
  assign q_617_clock = clock;
  assign q_617_reset = reset;
  assign q_617_io_enq_valid = cols_9_6_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_617_io_enq_bits = cols_9_6_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_617_io_deq_ready = io_value_out_6_9_ready; // @[Stab.scala 104:101]
  assign q_618_clock = clock;
  assign q_618_reset = reset;
  assign q_618_io_enq_valid = cols_10_6_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_618_io_enq_bits = cols_10_6_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_618_io_deq_ready = io_value_out_6_10_ready; // @[Stab.scala 104:101]
  assign q_619_clock = clock;
  assign q_619_reset = reset;
  assign q_619_io_enq_valid = cols_11_6_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_619_io_enq_bits = cols_11_6_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_619_io_deq_ready = io_value_out_6_11_ready; // @[Stab.scala 104:101]
  assign q_620_clock = clock;
  assign q_620_reset = reset;
  assign q_620_io_enq_valid = cols_12_6_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_620_io_enq_bits = cols_12_6_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_620_io_deq_ready = io_value_out_6_12_ready; // @[Stab.scala 104:101]
  assign q_621_clock = clock;
  assign q_621_reset = reset;
  assign q_621_io_enq_valid = cols_13_6_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_621_io_enq_bits = cols_13_6_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_621_io_deq_ready = io_value_out_6_13_ready; // @[Stab.scala 104:101]
  assign q_622_clock = clock;
  assign q_622_reset = reset;
  assign q_622_io_enq_valid = cols_14_6_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_622_io_enq_bits = cols_14_6_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_622_io_deq_ready = io_value_out_6_14_ready; // @[Stab.scala 104:101]
  assign q_623_clock = clock;
  assign q_623_reset = reset;
  assign q_623_io_enq_valid = cols_15_6_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_623_io_enq_bits = cols_15_6_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_623_io_deq_ready = io_value_out_6_15_ready; // @[Stab.scala 104:101]
  assign q_624_clock = clock;
  assign q_624_reset = reset;
  assign q_624_io_enq_valid = cols_0_7_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_624_io_enq_bits = cols_0_7_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_624_io_deq_ready = io_value_out_7_0_ready; // @[Stab.scala 104:101]
  assign q_625_clock = clock;
  assign q_625_reset = reset;
  assign q_625_io_enq_valid = cols_1_7_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_625_io_enq_bits = cols_1_7_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_625_io_deq_ready = io_value_out_7_1_ready; // @[Stab.scala 104:101]
  assign q_626_clock = clock;
  assign q_626_reset = reset;
  assign q_626_io_enq_valid = cols_2_7_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_626_io_enq_bits = cols_2_7_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_626_io_deq_ready = io_value_out_7_2_ready; // @[Stab.scala 104:101]
  assign q_627_clock = clock;
  assign q_627_reset = reset;
  assign q_627_io_enq_valid = cols_3_7_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_627_io_enq_bits = cols_3_7_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_627_io_deq_ready = io_value_out_7_3_ready; // @[Stab.scala 104:101]
  assign q_628_clock = clock;
  assign q_628_reset = reset;
  assign q_628_io_enq_valid = cols_4_7_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_628_io_enq_bits = cols_4_7_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_628_io_deq_ready = io_value_out_7_4_ready; // @[Stab.scala 104:101]
  assign q_629_clock = clock;
  assign q_629_reset = reset;
  assign q_629_io_enq_valid = cols_5_7_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_629_io_enq_bits = cols_5_7_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_629_io_deq_ready = io_value_out_7_5_ready; // @[Stab.scala 104:101]
  assign q_630_clock = clock;
  assign q_630_reset = reset;
  assign q_630_io_enq_valid = cols_6_7_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_630_io_enq_bits = cols_6_7_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_630_io_deq_ready = io_value_out_7_6_ready; // @[Stab.scala 104:101]
  assign q_631_clock = clock;
  assign q_631_reset = reset;
  assign q_631_io_enq_valid = cols_7_7_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_631_io_enq_bits = cols_7_7_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_631_io_deq_ready = io_value_out_7_7_ready; // @[Stab.scala 104:101]
  assign q_632_clock = clock;
  assign q_632_reset = reset;
  assign q_632_io_enq_valid = cols_8_7_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_632_io_enq_bits = cols_8_7_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_632_io_deq_ready = io_value_out_7_8_ready; // @[Stab.scala 104:101]
  assign q_633_clock = clock;
  assign q_633_reset = reset;
  assign q_633_io_enq_valid = cols_9_7_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_633_io_enq_bits = cols_9_7_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_633_io_deq_ready = io_value_out_7_9_ready; // @[Stab.scala 104:101]
  assign q_634_clock = clock;
  assign q_634_reset = reset;
  assign q_634_io_enq_valid = cols_10_7_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_634_io_enq_bits = cols_10_7_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_634_io_deq_ready = io_value_out_7_10_ready; // @[Stab.scala 104:101]
  assign q_635_clock = clock;
  assign q_635_reset = reset;
  assign q_635_io_enq_valid = cols_11_7_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_635_io_enq_bits = cols_11_7_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_635_io_deq_ready = io_value_out_7_11_ready; // @[Stab.scala 104:101]
  assign q_636_clock = clock;
  assign q_636_reset = reset;
  assign q_636_io_enq_valid = cols_12_7_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_636_io_enq_bits = cols_12_7_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_636_io_deq_ready = io_value_out_7_12_ready; // @[Stab.scala 104:101]
  assign q_637_clock = clock;
  assign q_637_reset = reset;
  assign q_637_io_enq_valid = cols_13_7_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_637_io_enq_bits = cols_13_7_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_637_io_deq_ready = io_value_out_7_13_ready; // @[Stab.scala 104:101]
  assign q_638_clock = clock;
  assign q_638_reset = reset;
  assign q_638_io_enq_valid = cols_14_7_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_638_io_enq_bits = cols_14_7_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_638_io_deq_ready = io_value_out_7_14_ready; // @[Stab.scala 104:101]
  assign q_639_clock = clock;
  assign q_639_reset = reset;
  assign q_639_io_enq_valid = cols_15_7_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_639_io_enq_bits = cols_15_7_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_639_io_deq_ready = io_value_out_7_15_ready; // @[Stab.scala 104:101]
  assign q_640_clock = clock;
  assign q_640_reset = reset;
  assign q_640_io_enq_valid = cols_0_8_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_640_io_enq_bits = cols_0_8_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_640_io_deq_ready = io_value_out_8_0_ready; // @[Stab.scala 104:101]
  assign q_641_clock = clock;
  assign q_641_reset = reset;
  assign q_641_io_enq_valid = cols_1_8_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_641_io_enq_bits = cols_1_8_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_641_io_deq_ready = io_value_out_8_1_ready; // @[Stab.scala 104:101]
  assign q_642_clock = clock;
  assign q_642_reset = reset;
  assign q_642_io_enq_valid = cols_2_8_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_642_io_enq_bits = cols_2_8_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_642_io_deq_ready = io_value_out_8_2_ready; // @[Stab.scala 104:101]
  assign q_643_clock = clock;
  assign q_643_reset = reset;
  assign q_643_io_enq_valid = cols_3_8_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_643_io_enq_bits = cols_3_8_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_643_io_deq_ready = io_value_out_8_3_ready; // @[Stab.scala 104:101]
  assign q_644_clock = clock;
  assign q_644_reset = reset;
  assign q_644_io_enq_valid = cols_4_8_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_644_io_enq_bits = cols_4_8_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_644_io_deq_ready = io_value_out_8_4_ready; // @[Stab.scala 104:101]
  assign q_645_clock = clock;
  assign q_645_reset = reset;
  assign q_645_io_enq_valid = cols_5_8_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_645_io_enq_bits = cols_5_8_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_645_io_deq_ready = io_value_out_8_5_ready; // @[Stab.scala 104:101]
  assign q_646_clock = clock;
  assign q_646_reset = reset;
  assign q_646_io_enq_valid = cols_6_8_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_646_io_enq_bits = cols_6_8_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_646_io_deq_ready = io_value_out_8_6_ready; // @[Stab.scala 104:101]
  assign q_647_clock = clock;
  assign q_647_reset = reset;
  assign q_647_io_enq_valid = cols_7_8_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_647_io_enq_bits = cols_7_8_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_647_io_deq_ready = io_value_out_8_7_ready; // @[Stab.scala 104:101]
  assign q_648_clock = clock;
  assign q_648_reset = reset;
  assign q_648_io_enq_valid = cols_8_8_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_648_io_enq_bits = cols_8_8_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_648_io_deq_ready = io_value_out_8_8_ready; // @[Stab.scala 104:101]
  assign q_649_clock = clock;
  assign q_649_reset = reset;
  assign q_649_io_enq_valid = cols_9_8_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_649_io_enq_bits = cols_9_8_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_649_io_deq_ready = io_value_out_8_9_ready; // @[Stab.scala 104:101]
  assign q_650_clock = clock;
  assign q_650_reset = reset;
  assign q_650_io_enq_valid = cols_10_8_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_650_io_enq_bits = cols_10_8_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_650_io_deq_ready = io_value_out_8_10_ready; // @[Stab.scala 104:101]
  assign q_651_clock = clock;
  assign q_651_reset = reset;
  assign q_651_io_enq_valid = cols_11_8_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_651_io_enq_bits = cols_11_8_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_651_io_deq_ready = io_value_out_8_11_ready; // @[Stab.scala 104:101]
  assign q_652_clock = clock;
  assign q_652_reset = reset;
  assign q_652_io_enq_valid = cols_12_8_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_652_io_enq_bits = cols_12_8_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_652_io_deq_ready = io_value_out_8_12_ready; // @[Stab.scala 104:101]
  assign q_653_clock = clock;
  assign q_653_reset = reset;
  assign q_653_io_enq_valid = cols_13_8_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_653_io_enq_bits = cols_13_8_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_653_io_deq_ready = io_value_out_8_13_ready; // @[Stab.scala 104:101]
  assign q_654_clock = clock;
  assign q_654_reset = reset;
  assign q_654_io_enq_valid = cols_14_8_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_654_io_enq_bits = cols_14_8_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_654_io_deq_ready = io_value_out_8_14_ready; // @[Stab.scala 104:101]
  assign q_655_clock = clock;
  assign q_655_reset = reset;
  assign q_655_io_enq_valid = cols_15_8_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_655_io_enq_bits = cols_15_8_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_655_io_deq_ready = io_value_out_8_15_ready; // @[Stab.scala 104:101]
  assign q_656_clock = clock;
  assign q_656_reset = reset;
  assign q_656_io_enq_valid = cols_0_9_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_656_io_enq_bits = cols_0_9_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_656_io_deq_ready = io_value_out_9_0_ready; // @[Stab.scala 104:101]
  assign q_657_clock = clock;
  assign q_657_reset = reset;
  assign q_657_io_enq_valid = cols_1_9_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_657_io_enq_bits = cols_1_9_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_657_io_deq_ready = io_value_out_9_1_ready; // @[Stab.scala 104:101]
  assign q_658_clock = clock;
  assign q_658_reset = reset;
  assign q_658_io_enq_valid = cols_2_9_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_658_io_enq_bits = cols_2_9_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_658_io_deq_ready = io_value_out_9_2_ready; // @[Stab.scala 104:101]
  assign q_659_clock = clock;
  assign q_659_reset = reset;
  assign q_659_io_enq_valid = cols_3_9_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_659_io_enq_bits = cols_3_9_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_659_io_deq_ready = io_value_out_9_3_ready; // @[Stab.scala 104:101]
  assign q_660_clock = clock;
  assign q_660_reset = reset;
  assign q_660_io_enq_valid = cols_4_9_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_660_io_enq_bits = cols_4_9_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_660_io_deq_ready = io_value_out_9_4_ready; // @[Stab.scala 104:101]
  assign q_661_clock = clock;
  assign q_661_reset = reset;
  assign q_661_io_enq_valid = cols_5_9_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_661_io_enq_bits = cols_5_9_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_661_io_deq_ready = io_value_out_9_5_ready; // @[Stab.scala 104:101]
  assign q_662_clock = clock;
  assign q_662_reset = reset;
  assign q_662_io_enq_valid = cols_6_9_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_662_io_enq_bits = cols_6_9_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_662_io_deq_ready = io_value_out_9_6_ready; // @[Stab.scala 104:101]
  assign q_663_clock = clock;
  assign q_663_reset = reset;
  assign q_663_io_enq_valid = cols_7_9_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_663_io_enq_bits = cols_7_9_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_663_io_deq_ready = io_value_out_9_7_ready; // @[Stab.scala 104:101]
  assign q_664_clock = clock;
  assign q_664_reset = reset;
  assign q_664_io_enq_valid = cols_8_9_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_664_io_enq_bits = cols_8_9_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_664_io_deq_ready = io_value_out_9_8_ready; // @[Stab.scala 104:101]
  assign q_665_clock = clock;
  assign q_665_reset = reset;
  assign q_665_io_enq_valid = cols_9_9_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_665_io_enq_bits = cols_9_9_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_665_io_deq_ready = io_value_out_9_9_ready; // @[Stab.scala 104:101]
  assign q_666_clock = clock;
  assign q_666_reset = reset;
  assign q_666_io_enq_valid = cols_10_9_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_666_io_enq_bits = cols_10_9_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_666_io_deq_ready = io_value_out_9_10_ready; // @[Stab.scala 104:101]
  assign q_667_clock = clock;
  assign q_667_reset = reset;
  assign q_667_io_enq_valid = cols_11_9_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_667_io_enq_bits = cols_11_9_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_667_io_deq_ready = io_value_out_9_11_ready; // @[Stab.scala 104:101]
  assign q_668_clock = clock;
  assign q_668_reset = reset;
  assign q_668_io_enq_valid = cols_12_9_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_668_io_enq_bits = cols_12_9_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_668_io_deq_ready = io_value_out_9_12_ready; // @[Stab.scala 104:101]
  assign q_669_clock = clock;
  assign q_669_reset = reset;
  assign q_669_io_enq_valid = cols_13_9_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_669_io_enq_bits = cols_13_9_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_669_io_deq_ready = io_value_out_9_13_ready; // @[Stab.scala 104:101]
  assign q_670_clock = clock;
  assign q_670_reset = reset;
  assign q_670_io_enq_valid = cols_14_9_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_670_io_enq_bits = cols_14_9_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_670_io_deq_ready = io_value_out_9_14_ready; // @[Stab.scala 104:101]
  assign q_671_clock = clock;
  assign q_671_reset = reset;
  assign q_671_io_enq_valid = cols_15_9_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_671_io_enq_bits = cols_15_9_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_671_io_deq_ready = io_value_out_9_15_ready; // @[Stab.scala 104:101]
  assign q_672_clock = clock;
  assign q_672_reset = reset;
  assign q_672_io_enq_valid = cols_0_10_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_672_io_enq_bits = cols_0_10_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_672_io_deq_ready = io_value_out_10_0_ready; // @[Stab.scala 104:101]
  assign q_673_clock = clock;
  assign q_673_reset = reset;
  assign q_673_io_enq_valid = cols_1_10_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_673_io_enq_bits = cols_1_10_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_673_io_deq_ready = io_value_out_10_1_ready; // @[Stab.scala 104:101]
  assign q_674_clock = clock;
  assign q_674_reset = reset;
  assign q_674_io_enq_valid = cols_2_10_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_674_io_enq_bits = cols_2_10_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_674_io_deq_ready = io_value_out_10_2_ready; // @[Stab.scala 104:101]
  assign q_675_clock = clock;
  assign q_675_reset = reset;
  assign q_675_io_enq_valid = cols_3_10_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_675_io_enq_bits = cols_3_10_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_675_io_deq_ready = io_value_out_10_3_ready; // @[Stab.scala 104:101]
  assign q_676_clock = clock;
  assign q_676_reset = reset;
  assign q_676_io_enq_valid = cols_4_10_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_676_io_enq_bits = cols_4_10_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_676_io_deq_ready = io_value_out_10_4_ready; // @[Stab.scala 104:101]
  assign q_677_clock = clock;
  assign q_677_reset = reset;
  assign q_677_io_enq_valid = cols_5_10_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_677_io_enq_bits = cols_5_10_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_677_io_deq_ready = io_value_out_10_5_ready; // @[Stab.scala 104:101]
  assign q_678_clock = clock;
  assign q_678_reset = reset;
  assign q_678_io_enq_valid = cols_6_10_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_678_io_enq_bits = cols_6_10_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_678_io_deq_ready = io_value_out_10_6_ready; // @[Stab.scala 104:101]
  assign q_679_clock = clock;
  assign q_679_reset = reset;
  assign q_679_io_enq_valid = cols_7_10_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_679_io_enq_bits = cols_7_10_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_679_io_deq_ready = io_value_out_10_7_ready; // @[Stab.scala 104:101]
  assign q_680_clock = clock;
  assign q_680_reset = reset;
  assign q_680_io_enq_valid = cols_8_10_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_680_io_enq_bits = cols_8_10_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_680_io_deq_ready = io_value_out_10_8_ready; // @[Stab.scala 104:101]
  assign q_681_clock = clock;
  assign q_681_reset = reset;
  assign q_681_io_enq_valid = cols_9_10_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_681_io_enq_bits = cols_9_10_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_681_io_deq_ready = io_value_out_10_9_ready; // @[Stab.scala 104:101]
  assign q_682_clock = clock;
  assign q_682_reset = reset;
  assign q_682_io_enq_valid = cols_10_10_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_682_io_enq_bits = cols_10_10_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_682_io_deq_ready = io_value_out_10_10_ready; // @[Stab.scala 104:101]
  assign q_683_clock = clock;
  assign q_683_reset = reset;
  assign q_683_io_enq_valid = cols_11_10_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_683_io_enq_bits = cols_11_10_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_683_io_deq_ready = io_value_out_10_11_ready; // @[Stab.scala 104:101]
  assign q_684_clock = clock;
  assign q_684_reset = reset;
  assign q_684_io_enq_valid = cols_12_10_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_684_io_enq_bits = cols_12_10_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_684_io_deq_ready = io_value_out_10_12_ready; // @[Stab.scala 104:101]
  assign q_685_clock = clock;
  assign q_685_reset = reset;
  assign q_685_io_enq_valid = cols_13_10_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_685_io_enq_bits = cols_13_10_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_685_io_deq_ready = io_value_out_10_13_ready; // @[Stab.scala 104:101]
  assign q_686_clock = clock;
  assign q_686_reset = reset;
  assign q_686_io_enq_valid = cols_14_10_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_686_io_enq_bits = cols_14_10_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_686_io_deq_ready = io_value_out_10_14_ready; // @[Stab.scala 104:101]
  assign q_687_clock = clock;
  assign q_687_reset = reset;
  assign q_687_io_enq_valid = cols_15_10_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_687_io_enq_bits = cols_15_10_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_687_io_deq_ready = io_value_out_10_15_ready; // @[Stab.scala 104:101]
  assign q_688_clock = clock;
  assign q_688_reset = reset;
  assign q_688_io_enq_valid = cols_0_11_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_688_io_enq_bits = cols_0_11_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_688_io_deq_ready = io_value_out_11_0_ready; // @[Stab.scala 104:101]
  assign q_689_clock = clock;
  assign q_689_reset = reset;
  assign q_689_io_enq_valid = cols_1_11_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_689_io_enq_bits = cols_1_11_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_689_io_deq_ready = io_value_out_11_1_ready; // @[Stab.scala 104:101]
  assign q_690_clock = clock;
  assign q_690_reset = reset;
  assign q_690_io_enq_valid = cols_2_11_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_690_io_enq_bits = cols_2_11_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_690_io_deq_ready = io_value_out_11_2_ready; // @[Stab.scala 104:101]
  assign q_691_clock = clock;
  assign q_691_reset = reset;
  assign q_691_io_enq_valid = cols_3_11_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_691_io_enq_bits = cols_3_11_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_691_io_deq_ready = io_value_out_11_3_ready; // @[Stab.scala 104:101]
  assign q_692_clock = clock;
  assign q_692_reset = reset;
  assign q_692_io_enq_valid = cols_4_11_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_692_io_enq_bits = cols_4_11_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_692_io_deq_ready = io_value_out_11_4_ready; // @[Stab.scala 104:101]
  assign q_693_clock = clock;
  assign q_693_reset = reset;
  assign q_693_io_enq_valid = cols_5_11_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_693_io_enq_bits = cols_5_11_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_693_io_deq_ready = io_value_out_11_5_ready; // @[Stab.scala 104:101]
  assign q_694_clock = clock;
  assign q_694_reset = reset;
  assign q_694_io_enq_valid = cols_6_11_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_694_io_enq_bits = cols_6_11_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_694_io_deq_ready = io_value_out_11_6_ready; // @[Stab.scala 104:101]
  assign q_695_clock = clock;
  assign q_695_reset = reset;
  assign q_695_io_enq_valid = cols_7_11_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_695_io_enq_bits = cols_7_11_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_695_io_deq_ready = io_value_out_11_7_ready; // @[Stab.scala 104:101]
  assign q_696_clock = clock;
  assign q_696_reset = reset;
  assign q_696_io_enq_valid = cols_8_11_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_696_io_enq_bits = cols_8_11_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_696_io_deq_ready = io_value_out_11_8_ready; // @[Stab.scala 104:101]
  assign q_697_clock = clock;
  assign q_697_reset = reset;
  assign q_697_io_enq_valid = cols_9_11_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_697_io_enq_bits = cols_9_11_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_697_io_deq_ready = io_value_out_11_9_ready; // @[Stab.scala 104:101]
  assign q_698_clock = clock;
  assign q_698_reset = reset;
  assign q_698_io_enq_valid = cols_10_11_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_698_io_enq_bits = cols_10_11_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_698_io_deq_ready = io_value_out_11_10_ready; // @[Stab.scala 104:101]
  assign q_699_clock = clock;
  assign q_699_reset = reset;
  assign q_699_io_enq_valid = cols_11_11_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_699_io_enq_bits = cols_11_11_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_699_io_deq_ready = io_value_out_11_11_ready; // @[Stab.scala 104:101]
  assign q_700_clock = clock;
  assign q_700_reset = reset;
  assign q_700_io_enq_valid = cols_12_11_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_700_io_enq_bits = cols_12_11_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_700_io_deq_ready = io_value_out_11_12_ready; // @[Stab.scala 104:101]
  assign q_701_clock = clock;
  assign q_701_reset = reset;
  assign q_701_io_enq_valid = cols_13_11_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_701_io_enq_bits = cols_13_11_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_701_io_deq_ready = io_value_out_11_13_ready; // @[Stab.scala 104:101]
  assign q_702_clock = clock;
  assign q_702_reset = reset;
  assign q_702_io_enq_valid = cols_14_11_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_702_io_enq_bits = cols_14_11_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_702_io_deq_ready = io_value_out_11_14_ready; // @[Stab.scala 104:101]
  assign q_703_clock = clock;
  assign q_703_reset = reset;
  assign q_703_io_enq_valid = cols_15_11_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_703_io_enq_bits = cols_15_11_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_703_io_deq_ready = io_value_out_11_15_ready; // @[Stab.scala 104:101]
  assign q_704_clock = clock;
  assign q_704_reset = reset;
  assign q_704_io_enq_valid = cols_0_12_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_704_io_enq_bits = cols_0_12_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_704_io_deq_ready = io_value_out_12_0_ready; // @[Stab.scala 104:101]
  assign q_705_clock = clock;
  assign q_705_reset = reset;
  assign q_705_io_enq_valid = cols_1_12_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_705_io_enq_bits = cols_1_12_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_705_io_deq_ready = io_value_out_12_1_ready; // @[Stab.scala 104:101]
  assign q_706_clock = clock;
  assign q_706_reset = reset;
  assign q_706_io_enq_valid = cols_2_12_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_706_io_enq_bits = cols_2_12_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_706_io_deq_ready = io_value_out_12_2_ready; // @[Stab.scala 104:101]
  assign q_707_clock = clock;
  assign q_707_reset = reset;
  assign q_707_io_enq_valid = cols_3_12_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_707_io_enq_bits = cols_3_12_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_707_io_deq_ready = io_value_out_12_3_ready; // @[Stab.scala 104:101]
  assign q_708_clock = clock;
  assign q_708_reset = reset;
  assign q_708_io_enq_valid = cols_4_12_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_708_io_enq_bits = cols_4_12_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_708_io_deq_ready = io_value_out_12_4_ready; // @[Stab.scala 104:101]
  assign q_709_clock = clock;
  assign q_709_reset = reset;
  assign q_709_io_enq_valid = cols_5_12_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_709_io_enq_bits = cols_5_12_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_709_io_deq_ready = io_value_out_12_5_ready; // @[Stab.scala 104:101]
  assign q_710_clock = clock;
  assign q_710_reset = reset;
  assign q_710_io_enq_valid = cols_6_12_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_710_io_enq_bits = cols_6_12_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_710_io_deq_ready = io_value_out_12_6_ready; // @[Stab.scala 104:101]
  assign q_711_clock = clock;
  assign q_711_reset = reset;
  assign q_711_io_enq_valid = cols_7_12_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_711_io_enq_bits = cols_7_12_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_711_io_deq_ready = io_value_out_12_7_ready; // @[Stab.scala 104:101]
  assign q_712_clock = clock;
  assign q_712_reset = reset;
  assign q_712_io_enq_valid = cols_8_12_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_712_io_enq_bits = cols_8_12_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_712_io_deq_ready = io_value_out_12_8_ready; // @[Stab.scala 104:101]
  assign q_713_clock = clock;
  assign q_713_reset = reset;
  assign q_713_io_enq_valid = cols_9_12_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_713_io_enq_bits = cols_9_12_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_713_io_deq_ready = io_value_out_12_9_ready; // @[Stab.scala 104:101]
  assign q_714_clock = clock;
  assign q_714_reset = reset;
  assign q_714_io_enq_valid = cols_10_12_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_714_io_enq_bits = cols_10_12_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_714_io_deq_ready = io_value_out_12_10_ready; // @[Stab.scala 104:101]
  assign q_715_clock = clock;
  assign q_715_reset = reset;
  assign q_715_io_enq_valid = cols_11_12_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_715_io_enq_bits = cols_11_12_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_715_io_deq_ready = io_value_out_12_11_ready; // @[Stab.scala 104:101]
  assign q_716_clock = clock;
  assign q_716_reset = reset;
  assign q_716_io_enq_valid = cols_12_12_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_716_io_enq_bits = cols_12_12_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_716_io_deq_ready = io_value_out_12_12_ready; // @[Stab.scala 104:101]
  assign q_717_clock = clock;
  assign q_717_reset = reset;
  assign q_717_io_enq_valid = cols_13_12_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_717_io_enq_bits = cols_13_12_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_717_io_deq_ready = io_value_out_12_13_ready; // @[Stab.scala 104:101]
  assign q_718_clock = clock;
  assign q_718_reset = reset;
  assign q_718_io_enq_valid = cols_14_12_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_718_io_enq_bits = cols_14_12_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_718_io_deq_ready = io_value_out_12_14_ready; // @[Stab.scala 104:101]
  assign q_719_clock = clock;
  assign q_719_reset = reset;
  assign q_719_io_enq_valid = cols_15_12_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_719_io_enq_bits = cols_15_12_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_719_io_deq_ready = io_value_out_12_15_ready; // @[Stab.scala 104:101]
  assign q_720_clock = clock;
  assign q_720_reset = reset;
  assign q_720_io_enq_valid = cols_0_13_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_720_io_enq_bits = cols_0_13_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_720_io_deq_ready = io_value_out_13_0_ready; // @[Stab.scala 104:101]
  assign q_721_clock = clock;
  assign q_721_reset = reset;
  assign q_721_io_enq_valid = cols_1_13_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_721_io_enq_bits = cols_1_13_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_721_io_deq_ready = io_value_out_13_1_ready; // @[Stab.scala 104:101]
  assign q_722_clock = clock;
  assign q_722_reset = reset;
  assign q_722_io_enq_valid = cols_2_13_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_722_io_enq_bits = cols_2_13_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_722_io_deq_ready = io_value_out_13_2_ready; // @[Stab.scala 104:101]
  assign q_723_clock = clock;
  assign q_723_reset = reset;
  assign q_723_io_enq_valid = cols_3_13_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_723_io_enq_bits = cols_3_13_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_723_io_deq_ready = io_value_out_13_3_ready; // @[Stab.scala 104:101]
  assign q_724_clock = clock;
  assign q_724_reset = reset;
  assign q_724_io_enq_valid = cols_4_13_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_724_io_enq_bits = cols_4_13_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_724_io_deq_ready = io_value_out_13_4_ready; // @[Stab.scala 104:101]
  assign q_725_clock = clock;
  assign q_725_reset = reset;
  assign q_725_io_enq_valid = cols_5_13_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_725_io_enq_bits = cols_5_13_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_725_io_deq_ready = io_value_out_13_5_ready; // @[Stab.scala 104:101]
  assign q_726_clock = clock;
  assign q_726_reset = reset;
  assign q_726_io_enq_valid = cols_6_13_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_726_io_enq_bits = cols_6_13_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_726_io_deq_ready = io_value_out_13_6_ready; // @[Stab.scala 104:101]
  assign q_727_clock = clock;
  assign q_727_reset = reset;
  assign q_727_io_enq_valid = cols_7_13_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_727_io_enq_bits = cols_7_13_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_727_io_deq_ready = io_value_out_13_7_ready; // @[Stab.scala 104:101]
  assign q_728_clock = clock;
  assign q_728_reset = reset;
  assign q_728_io_enq_valid = cols_8_13_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_728_io_enq_bits = cols_8_13_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_728_io_deq_ready = io_value_out_13_8_ready; // @[Stab.scala 104:101]
  assign q_729_clock = clock;
  assign q_729_reset = reset;
  assign q_729_io_enq_valid = cols_9_13_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_729_io_enq_bits = cols_9_13_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_729_io_deq_ready = io_value_out_13_9_ready; // @[Stab.scala 104:101]
  assign q_730_clock = clock;
  assign q_730_reset = reset;
  assign q_730_io_enq_valid = cols_10_13_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_730_io_enq_bits = cols_10_13_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_730_io_deq_ready = io_value_out_13_10_ready; // @[Stab.scala 104:101]
  assign q_731_clock = clock;
  assign q_731_reset = reset;
  assign q_731_io_enq_valid = cols_11_13_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_731_io_enq_bits = cols_11_13_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_731_io_deq_ready = io_value_out_13_11_ready; // @[Stab.scala 104:101]
  assign q_732_clock = clock;
  assign q_732_reset = reset;
  assign q_732_io_enq_valid = cols_12_13_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_732_io_enq_bits = cols_12_13_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_732_io_deq_ready = io_value_out_13_12_ready; // @[Stab.scala 104:101]
  assign q_733_clock = clock;
  assign q_733_reset = reset;
  assign q_733_io_enq_valid = cols_13_13_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_733_io_enq_bits = cols_13_13_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_733_io_deq_ready = io_value_out_13_13_ready; // @[Stab.scala 104:101]
  assign q_734_clock = clock;
  assign q_734_reset = reset;
  assign q_734_io_enq_valid = cols_14_13_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_734_io_enq_bits = cols_14_13_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_734_io_deq_ready = io_value_out_13_14_ready; // @[Stab.scala 104:101]
  assign q_735_clock = clock;
  assign q_735_reset = reset;
  assign q_735_io_enq_valid = cols_15_13_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_735_io_enq_bits = cols_15_13_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_735_io_deq_ready = io_value_out_13_15_ready; // @[Stab.scala 104:101]
  assign q_736_clock = clock;
  assign q_736_reset = reset;
  assign q_736_io_enq_valid = cols_0_14_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_736_io_enq_bits = cols_0_14_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_736_io_deq_ready = io_value_out_14_0_ready; // @[Stab.scala 104:101]
  assign q_737_clock = clock;
  assign q_737_reset = reset;
  assign q_737_io_enq_valid = cols_1_14_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_737_io_enq_bits = cols_1_14_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_737_io_deq_ready = io_value_out_14_1_ready; // @[Stab.scala 104:101]
  assign q_738_clock = clock;
  assign q_738_reset = reset;
  assign q_738_io_enq_valid = cols_2_14_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_738_io_enq_bits = cols_2_14_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_738_io_deq_ready = io_value_out_14_2_ready; // @[Stab.scala 104:101]
  assign q_739_clock = clock;
  assign q_739_reset = reset;
  assign q_739_io_enq_valid = cols_3_14_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_739_io_enq_bits = cols_3_14_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_739_io_deq_ready = io_value_out_14_3_ready; // @[Stab.scala 104:101]
  assign q_740_clock = clock;
  assign q_740_reset = reset;
  assign q_740_io_enq_valid = cols_4_14_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_740_io_enq_bits = cols_4_14_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_740_io_deq_ready = io_value_out_14_4_ready; // @[Stab.scala 104:101]
  assign q_741_clock = clock;
  assign q_741_reset = reset;
  assign q_741_io_enq_valid = cols_5_14_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_741_io_enq_bits = cols_5_14_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_741_io_deq_ready = io_value_out_14_5_ready; // @[Stab.scala 104:101]
  assign q_742_clock = clock;
  assign q_742_reset = reset;
  assign q_742_io_enq_valid = cols_6_14_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_742_io_enq_bits = cols_6_14_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_742_io_deq_ready = io_value_out_14_6_ready; // @[Stab.scala 104:101]
  assign q_743_clock = clock;
  assign q_743_reset = reset;
  assign q_743_io_enq_valid = cols_7_14_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_743_io_enq_bits = cols_7_14_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_743_io_deq_ready = io_value_out_14_7_ready; // @[Stab.scala 104:101]
  assign q_744_clock = clock;
  assign q_744_reset = reset;
  assign q_744_io_enq_valid = cols_8_14_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_744_io_enq_bits = cols_8_14_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_744_io_deq_ready = io_value_out_14_8_ready; // @[Stab.scala 104:101]
  assign q_745_clock = clock;
  assign q_745_reset = reset;
  assign q_745_io_enq_valid = cols_9_14_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_745_io_enq_bits = cols_9_14_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_745_io_deq_ready = io_value_out_14_9_ready; // @[Stab.scala 104:101]
  assign q_746_clock = clock;
  assign q_746_reset = reset;
  assign q_746_io_enq_valid = cols_10_14_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_746_io_enq_bits = cols_10_14_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_746_io_deq_ready = io_value_out_14_10_ready; // @[Stab.scala 104:101]
  assign q_747_clock = clock;
  assign q_747_reset = reset;
  assign q_747_io_enq_valid = cols_11_14_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_747_io_enq_bits = cols_11_14_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_747_io_deq_ready = io_value_out_14_11_ready; // @[Stab.scala 104:101]
  assign q_748_clock = clock;
  assign q_748_reset = reset;
  assign q_748_io_enq_valid = cols_12_14_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_748_io_enq_bits = cols_12_14_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_748_io_deq_ready = io_value_out_14_12_ready; // @[Stab.scala 104:101]
  assign q_749_clock = clock;
  assign q_749_reset = reset;
  assign q_749_io_enq_valid = cols_13_14_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_749_io_enq_bits = cols_13_14_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_749_io_deq_ready = io_value_out_14_13_ready; // @[Stab.scala 104:101]
  assign q_750_clock = clock;
  assign q_750_reset = reset;
  assign q_750_io_enq_valid = cols_14_14_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_750_io_enq_bits = cols_14_14_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_750_io_deq_ready = io_value_out_14_14_ready; // @[Stab.scala 104:101]
  assign q_751_clock = clock;
  assign q_751_reset = reset;
  assign q_751_io_enq_valid = cols_15_14_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_751_io_enq_bits = cols_15_14_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_751_io_deq_ready = io_value_out_14_15_ready; // @[Stab.scala 104:101]
  assign q_752_clock = clock;
  assign q_752_reset = reset;
  assign q_752_io_enq_valid = cols_0_15_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_752_io_enq_bits = cols_0_15_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_752_io_deq_ready = io_value_out_15_0_ready; // @[Stab.scala 104:101]
  assign q_753_clock = clock;
  assign q_753_reset = reset;
  assign q_753_io_enq_valid = cols_1_15_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_753_io_enq_bits = cols_1_15_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_753_io_deq_ready = io_value_out_15_1_ready; // @[Stab.scala 104:101]
  assign q_754_clock = clock;
  assign q_754_reset = reset;
  assign q_754_io_enq_valid = cols_2_15_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_754_io_enq_bits = cols_2_15_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_754_io_deq_ready = io_value_out_15_2_ready; // @[Stab.scala 104:101]
  assign q_755_clock = clock;
  assign q_755_reset = reset;
  assign q_755_io_enq_valid = cols_3_15_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_755_io_enq_bits = cols_3_15_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_755_io_deq_ready = io_value_out_15_3_ready; // @[Stab.scala 104:101]
  assign q_756_clock = clock;
  assign q_756_reset = reset;
  assign q_756_io_enq_valid = cols_4_15_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_756_io_enq_bits = cols_4_15_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_756_io_deq_ready = io_value_out_15_4_ready; // @[Stab.scala 104:101]
  assign q_757_clock = clock;
  assign q_757_reset = reset;
  assign q_757_io_enq_valid = cols_5_15_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_757_io_enq_bits = cols_5_15_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_757_io_deq_ready = io_value_out_15_5_ready; // @[Stab.scala 104:101]
  assign q_758_clock = clock;
  assign q_758_reset = reset;
  assign q_758_io_enq_valid = cols_6_15_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_758_io_enq_bits = cols_6_15_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_758_io_deq_ready = io_value_out_15_6_ready; // @[Stab.scala 104:101]
  assign q_759_clock = clock;
  assign q_759_reset = reset;
  assign q_759_io_enq_valid = cols_7_15_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_759_io_enq_bits = cols_7_15_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_759_io_deq_ready = io_value_out_15_7_ready; // @[Stab.scala 104:101]
  assign q_760_clock = clock;
  assign q_760_reset = reset;
  assign q_760_io_enq_valid = cols_8_15_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_760_io_enq_bits = cols_8_15_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_760_io_deq_ready = io_value_out_15_8_ready; // @[Stab.scala 104:101]
  assign q_761_clock = clock;
  assign q_761_reset = reset;
  assign q_761_io_enq_valid = cols_9_15_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_761_io_enq_bits = cols_9_15_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_761_io_deq_ready = io_value_out_15_9_ready; // @[Stab.scala 104:101]
  assign q_762_clock = clock;
  assign q_762_reset = reset;
  assign q_762_io_enq_valid = cols_10_15_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_762_io_enq_bits = cols_10_15_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_762_io_deq_ready = io_value_out_15_10_ready; // @[Stab.scala 104:101]
  assign q_763_clock = clock;
  assign q_763_reset = reset;
  assign q_763_io_enq_valid = cols_11_15_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_763_io_enq_bits = cols_11_15_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_763_io_deq_ready = io_value_out_15_11_ready; // @[Stab.scala 104:101]
  assign q_764_clock = clock;
  assign q_764_reset = reset;
  assign q_764_io_enq_valid = cols_12_15_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_764_io_enq_bits = cols_12_15_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_764_io_deq_ready = io_value_out_15_12_ready; // @[Stab.scala 104:101]
  assign q_765_clock = clock;
  assign q_765_reset = reset;
  assign q_765_io_enq_valid = cols_13_15_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_765_io_enq_bits = cols_13_15_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_765_io_deq_ready = io_value_out_15_13_ready; // @[Stab.scala 104:101]
  assign q_766_clock = clock;
  assign q_766_reset = reset;
  assign q_766_io_enq_valid = cols_14_15_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_766_io_enq_bits = cols_14_15_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_766_io_deq_ready = io_value_out_15_14_ready; // @[Stab.scala 104:101]
  assign q_767_clock = clock;
  assign q_767_reset = reset;
  assign q_767_io_enq_valid = cols_15_15_io_sum_valid; // @[Decoupled.scala 363:22]
  assign q_767_io_enq_bits = cols_15_15_io_sum_bits; // @[Decoupled.scala 364:21]
  assign q_767_io_deq_ready = io_value_out_15_15_ready; // @[Stab.scala 104:101]
endmodule
module StreamSplitterBinaryTree(
  output        io_stream_in_ready,
  input         io_stream_in_valid,
  input  [31:0] io_stream_in_bits,
  input         io_stream_out_0_ready,
  output        io_stream_out_0_valid,
  output [31:0] io_stream_out_0_bits
);
  assign io_stream_in_ready = io_stream_out_0_ready; // @[Stab.scala 214:17]
  assign io_stream_out_0_valid = io_stream_in_valid; // @[Stab.scala 214:17]
  assign io_stream_out_0_bits = io_stream_in_bits; // @[Stab.scala 214:17]
endmodule
module StreamTranspose(
  input         clock,
  input         reset,
  output        io_stream_in_ready,
  input         io_stream_in_valid,
  input  [31:0] io_stream_in_bits,
  input         io_stream_out_0_ready,
  output        io_stream_out_0_valid,
  output [31:0] io_stream_out_0_bits,
  input         io_stream_out_1_ready,
  output        io_stream_out_1_valid,
  output [31:0] io_stream_out_1_bits,
  input         io_stream_out_2_ready,
  output        io_stream_out_2_valid,
  output [31:0] io_stream_out_2_bits,
  input         io_stream_out_3_ready,
  output        io_stream_out_3_valid,
  output [31:0] io_stream_out_3_bits,
  input         io_stream_out_4_ready,
  output        io_stream_out_4_valid,
  output [31:0] io_stream_out_4_bits,
  input         io_stream_out_5_ready,
  output        io_stream_out_5_valid,
  output [31:0] io_stream_out_5_bits,
  input         io_stream_out_6_ready,
  output        io_stream_out_6_valid,
  output [31:0] io_stream_out_6_bits,
  input         io_stream_out_7_ready,
  output        io_stream_out_7_valid,
  output [31:0] io_stream_out_7_bits,
  input         io_stream_out_8_ready,
  output        io_stream_out_8_valid,
  output [31:0] io_stream_out_8_bits,
  input         io_stream_out_9_ready,
  output        io_stream_out_9_valid,
  output [31:0] io_stream_out_9_bits,
  input         io_stream_out_10_ready,
  output        io_stream_out_10_valid,
  output [31:0] io_stream_out_10_bits,
  input         io_stream_out_11_ready,
  output        io_stream_out_11_valid,
  output [31:0] io_stream_out_11_bits,
  input         io_stream_out_12_ready,
  output        io_stream_out_12_valid,
  output [31:0] io_stream_out_12_bits,
  input         io_stream_out_13_ready,
  output        io_stream_out_13_valid,
  output [31:0] io_stream_out_13_bits,
  input         io_stream_out_14_ready,
  output        io_stream_out_14_valid,
  output [31:0] io_stream_out_14_bits,
  input         io_stream_out_15_ready,
  output        io_stream_out_15_valid,
  output [31:0] io_stream_out_15_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  splitters_0_io_stream_in_ready; // @[Stab.scala 230:46]
  wire  splitters_0_io_stream_in_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_0_io_stream_in_bits; // @[Stab.scala 230:46]
  wire  splitters_0_io_stream_out_0_ready; // @[Stab.scala 230:46]
  wire  splitters_0_io_stream_out_0_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_0_io_stream_out_0_bits; // @[Stab.scala 230:46]
  wire  splitters_1_io_stream_in_ready; // @[Stab.scala 230:46]
  wire  splitters_1_io_stream_in_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_1_io_stream_in_bits; // @[Stab.scala 230:46]
  wire  splitters_1_io_stream_out_0_ready; // @[Stab.scala 230:46]
  wire  splitters_1_io_stream_out_0_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_1_io_stream_out_0_bits; // @[Stab.scala 230:46]
  wire  splitters_2_io_stream_in_ready; // @[Stab.scala 230:46]
  wire  splitters_2_io_stream_in_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_2_io_stream_in_bits; // @[Stab.scala 230:46]
  wire  splitters_2_io_stream_out_0_ready; // @[Stab.scala 230:46]
  wire  splitters_2_io_stream_out_0_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_2_io_stream_out_0_bits; // @[Stab.scala 230:46]
  wire  splitters_3_io_stream_in_ready; // @[Stab.scala 230:46]
  wire  splitters_3_io_stream_in_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_3_io_stream_in_bits; // @[Stab.scala 230:46]
  wire  splitters_3_io_stream_out_0_ready; // @[Stab.scala 230:46]
  wire  splitters_3_io_stream_out_0_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_3_io_stream_out_0_bits; // @[Stab.scala 230:46]
  wire  splitters_4_io_stream_in_ready; // @[Stab.scala 230:46]
  wire  splitters_4_io_stream_in_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_4_io_stream_in_bits; // @[Stab.scala 230:46]
  wire  splitters_4_io_stream_out_0_ready; // @[Stab.scala 230:46]
  wire  splitters_4_io_stream_out_0_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_4_io_stream_out_0_bits; // @[Stab.scala 230:46]
  wire  splitters_5_io_stream_in_ready; // @[Stab.scala 230:46]
  wire  splitters_5_io_stream_in_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_5_io_stream_in_bits; // @[Stab.scala 230:46]
  wire  splitters_5_io_stream_out_0_ready; // @[Stab.scala 230:46]
  wire  splitters_5_io_stream_out_0_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_5_io_stream_out_0_bits; // @[Stab.scala 230:46]
  wire  splitters_6_io_stream_in_ready; // @[Stab.scala 230:46]
  wire  splitters_6_io_stream_in_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_6_io_stream_in_bits; // @[Stab.scala 230:46]
  wire  splitters_6_io_stream_out_0_ready; // @[Stab.scala 230:46]
  wire  splitters_6_io_stream_out_0_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_6_io_stream_out_0_bits; // @[Stab.scala 230:46]
  wire  splitters_7_io_stream_in_ready; // @[Stab.scala 230:46]
  wire  splitters_7_io_stream_in_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_7_io_stream_in_bits; // @[Stab.scala 230:46]
  wire  splitters_7_io_stream_out_0_ready; // @[Stab.scala 230:46]
  wire  splitters_7_io_stream_out_0_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_7_io_stream_out_0_bits; // @[Stab.scala 230:46]
  wire  splitters_8_io_stream_in_ready; // @[Stab.scala 230:46]
  wire  splitters_8_io_stream_in_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_8_io_stream_in_bits; // @[Stab.scala 230:46]
  wire  splitters_8_io_stream_out_0_ready; // @[Stab.scala 230:46]
  wire  splitters_8_io_stream_out_0_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_8_io_stream_out_0_bits; // @[Stab.scala 230:46]
  wire  splitters_9_io_stream_in_ready; // @[Stab.scala 230:46]
  wire  splitters_9_io_stream_in_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_9_io_stream_in_bits; // @[Stab.scala 230:46]
  wire  splitters_9_io_stream_out_0_ready; // @[Stab.scala 230:46]
  wire  splitters_9_io_stream_out_0_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_9_io_stream_out_0_bits; // @[Stab.scala 230:46]
  wire  splitters_10_io_stream_in_ready; // @[Stab.scala 230:46]
  wire  splitters_10_io_stream_in_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_10_io_stream_in_bits; // @[Stab.scala 230:46]
  wire  splitters_10_io_stream_out_0_ready; // @[Stab.scala 230:46]
  wire  splitters_10_io_stream_out_0_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_10_io_stream_out_0_bits; // @[Stab.scala 230:46]
  wire  splitters_11_io_stream_in_ready; // @[Stab.scala 230:46]
  wire  splitters_11_io_stream_in_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_11_io_stream_in_bits; // @[Stab.scala 230:46]
  wire  splitters_11_io_stream_out_0_ready; // @[Stab.scala 230:46]
  wire  splitters_11_io_stream_out_0_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_11_io_stream_out_0_bits; // @[Stab.scala 230:46]
  wire  splitters_12_io_stream_in_ready; // @[Stab.scala 230:46]
  wire  splitters_12_io_stream_in_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_12_io_stream_in_bits; // @[Stab.scala 230:46]
  wire  splitters_12_io_stream_out_0_ready; // @[Stab.scala 230:46]
  wire  splitters_12_io_stream_out_0_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_12_io_stream_out_0_bits; // @[Stab.scala 230:46]
  wire  splitters_13_io_stream_in_ready; // @[Stab.scala 230:46]
  wire  splitters_13_io_stream_in_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_13_io_stream_in_bits; // @[Stab.scala 230:46]
  wire  splitters_13_io_stream_out_0_ready; // @[Stab.scala 230:46]
  wire  splitters_13_io_stream_out_0_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_13_io_stream_out_0_bits; // @[Stab.scala 230:46]
  wire  splitters_14_io_stream_in_ready; // @[Stab.scala 230:46]
  wire  splitters_14_io_stream_in_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_14_io_stream_in_bits; // @[Stab.scala 230:46]
  wire  splitters_14_io_stream_out_0_ready; // @[Stab.scala 230:46]
  wire  splitters_14_io_stream_out_0_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_14_io_stream_out_0_bits; // @[Stab.scala 230:46]
  wire  splitters_15_io_stream_in_ready; // @[Stab.scala 230:46]
  wire  splitters_15_io_stream_in_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_15_io_stream_in_bits; // @[Stab.scala 230:46]
  wire  splitters_15_io_stream_out_0_ready; // @[Stab.scala 230:46]
  wire  splitters_15_io_stream_out_0_valid; // @[Stab.scala 230:46]
  wire [31:0] splitters_15_io_stream_out_0_bits; // @[Stab.scala 230:46]
  wire  _turn_T = io_stream_in_ready & io_stream_in_valid; // @[Decoupled.scala 50:35]
  reg [3:0] turn; // @[Counter.scala 62:40]
  wire  turn_wrap_wrap = turn == 4'hf; // @[Counter.scala 74:24]
  wire [3:0] _turn_wrap_value_T_1 = turn + 4'h1; // @[Counter.scala 78:24]
  wire  _splitters_0_io_stream_in_valid_T = turn == 4'h0; // @[Stab.scala 238:41]
  wire  _GEN_2 = _splitters_0_io_stream_in_valid_T & splitters_0_io_stream_in_ready; // @[Stab.scala 235:22 240:25 241:26]
  wire  _splitters_1_io_stream_in_valid_T = turn == 4'h1; // @[Stab.scala 238:41]
  wire  _GEN_3 = _splitters_1_io_stream_in_valid_T ? splitters_1_io_stream_in_ready : _GEN_2; // @[Stab.scala 240:25 241:26]
  wire  _splitters_2_io_stream_in_valid_T = turn == 4'h2; // @[Stab.scala 238:41]
  wire  _GEN_4 = _splitters_2_io_stream_in_valid_T ? splitters_2_io_stream_in_ready : _GEN_3; // @[Stab.scala 240:25 241:26]
  wire  _splitters_3_io_stream_in_valid_T = turn == 4'h3; // @[Stab.scala 238:41]
  wire  _GEN_5 = _splitters_3_io_stream_in_valid_T ? splitters_3_io_stream_in_ready : _GEN_4; // @[Stab.scala 240:25 241:26]
  wire  _splitters_4_io_stream_in_valid_T = turn == 4'h4; // @[Stab.scala 238:41]
  wire  _GEN_6 = _splitters_4_io_stream_in_valid_T ? splitters_4_io_stream_in_ready : _GEN_5; // @[Stab.scala 240:25 241:26]
  wire  _splitters_5_io_stream_in_valid_T = turn == 4'h5; // @[Stab.scala 238:41]
  wire  _GEN_7 = _splitters_5_io_stream_in_valid_T ? splitters_5_io_stream_in_ready : _GEN_6; // @[Stab.scala 240:25 241:26]
  wire  _splitters_6_io_stream_in_valid_T = turn == 4'h6; // @[Stab.scala 238:41]
  wire  _GEN_8 = _splitters_6_io_stream_in_valid_T ? splitters_6_io_stream_in_ready : _GEN_7; // @[Stab.scala 240:25 241:26]
  wire  _splitters_7_io_stream_in_valid_T = turn == 4'h7; // @[Stab.scala 238:41]
  wire  _GEN_9 = _splitters_7_io_stream_in_valid_T ? splitters_7_io_stream_in_ready : _GEN_8; // @[Stab.scala 240:25 241:26]
  wire  _splitters_8_io_stream_in_valid_T = turn == 4'h8; // @[Stab.scala 238:41]
  wire  _GEN_10 = _splitters_8_io_stream_in_valid_T ? splitters_8_io_stream_in_ready : _GEN_9; // @[Stab.scala 240:25 241:26]
  wire  _splitters_9_io_stream_in_valid_T = turn == 4'h9; // @[Stab.scala 238:41]
  wire  _GEN_11 = _splitters_9_io_stream_in_valid_T ? splitters_9_io_stream_in_ready : _GEN_10; // @[Stab.scala 240:25 241:26]
  wire  _splitters_10_io_stream_in_valid_T = turn == 4'ha; // @[Stab.scala 238:41]
  wire  _GEN_12 = _splitters_10_io_stream_in_valid_T ? splitters_10_io_stream_in_ready : _GEN_11; // @[Stab.scala 240:25 241:26]
  wire  _splitters_11_io_stream_in_valid_T = turn == 4'hb; // @[Stab.scala 238:41]
  wire  _GEN_13 = _splitters_11_io_stream_in_valid_T ? splitters_11_io_stream_in_ready : _GEN_12; // @[Stab.scala 240:25 241:26]
  wire  _splitters_12_io_stream_in_valid_T = turn == 4'hc; // @[Stab.scala 238:41]
  wire  _GEN_14 = _splitters_12_io_stream_in_valid_T ? splitters_12_io_stream_in_ready : _GEN_13; // @[Stab.scala 240:25 241:26]
  wire  _splitters_13_io_stream_in_valid_T = turn == 4'hd; // @[Stab.scala 238:41]
  wire  _GEN_15 = _splitters_13_io_stream_in_valid_T ? splitters_13_io_stream_in_ready : _GEN_14; // @[Stab.scala 240:25 241:26]
  wire  _splitters_14_io_stream_in_valid_T = turn == 4'he; // @[Stab.scala 238:41]
  wire  _GEN_16 = _splitters_14_io_stream_in_valid_T ? splitters_14_io_stream_in_ready : _GEN_15; // @[Stab.scala 240:25 241:26]
  StreamSplitterBinaryTree splitters_0 ( // @[Stab.scala 230:46]
    .io_stream_in_ready(splitters_0_io_stream_in_ready),
    .io_stream_in_valid(splitters_0_io_stream_in_valid),
    .io_stream_in_bits(splitters_0_io_stream_in_bits),
    .io_stream_out_0_ready(splitters_0_io_stream_out_0_ready),
    .io_stream_out_0_valid(splitters_0_io_stream_out_0_valid),
    .io_stream_out_0_bits(splitters_0_io_stream_out_0_bits)
  );
  StreamSplitterBinaryTree splitters_1 ( // @[Stab.scala 230:46]
    .io_stream_in_ready(splitters_1_io_stream_in_ready),
    .io_stream_in_valid(splitters_1_io_stream_in_valid),
    .io_stream_in_bits(splitters_1_io_stream_in_bits),
    .io_stream_out_0_ready(splitters_1_io_stream_out_0_ready),
    .io_stream_out_0_valid(splitters_1_io_stream_out_0_valid),
    .io_stream_out_0_bits(splitters_1_io_stream_out_0_bits)
  );
  StreamSplitterBinaryTree splitters_2 ( // @[Stab.scala 230:46]
    .io_stream_in_ready(splitters_2_io_stream_in_ready),
    .io_stream_in_valid(splitters_2_io_stream_in_valid),
    .io_stream_in_bits(splitters_2_io_stream_in_bits),
    .io_stream_out_0_ready(splitters_2_io_stream_out_0_ready),
    .io_stream_out_0_valid(splitters_2_io_stream_out_0_valid),
    .io_stream_out_0_bits(splitters_2_io_stream_out_0_bits)
  );
  StreamSplitterBinaryTree splitters_3 ( // @[Stab.scala 230:46]
    .io_stream_in_ready(splitters_3_io_stream_in_ready),
    .io_stream_in_valid(splitters_3_io_stream_in_valid),
    .io_stream_in_bits(splitters_3_io_stream_in_bits),
    .io_stream_out_0_ready(splitters_3_io_stream_out_0_ready),
    .io_stream_out_0_valid(splitters_3_io_stream_out_0_valid),
    .io_stream_out_0_bits(splitters_3_io_stream_out_0_bits)
  );
  StreamSplitterBinaryTree splitters_4 ( // @[Stab.scala 230:46]
    .io_stream_in_ready(splitters_4_io_stream_in_ready),
    .io_stream_in_valid(splitters_4_io_stream_in_valid),
    .io_stream_in_bits(splitters_4_io_stream_in_bits),
    .io_stream_out_0_ready(splitters_4_io_stream_out_0_ready),
    .io_stream_out_0_valid(splitters_4_io_stream_out_0_valid),
    .io_stream_out_0_bits(splitters_4_io_stream_out_0_bits)
  );
  StreamSplitterBinaryTree splitters_5 ( // @[Stab.scala 230:46]
    .io_stream_in_ready(splitters_5_io_stream_in_ready),
    .io_stream_in_valid(splitters_5_io_stream_in_valid),
    .io_stream_in_bits(splitters_5_io_stream_in_bits),
    .io_stream_out_0_ready(splitters_5_io_stream_out_0_ready),
    .io_stream_out_0_valid(splitters_5_io_stream_out_0_valid),
    .io_stream_out_0_bits(splitters_5_io_stream_out_0_bits)
  );
  StreamSplitterBinaryTree splitters_6 ( // @[Stab.scala 230:46]
    .io_stream_in_ready(splitters_6_io_stream_in_ready),
    .io_stream_in_valid(splitters_6_io_stream_in_valid),
    .io_stream_in_bits(splitters_6_io_stream_in_bits),
    .io_stream_out_0_ready(splitters_6_io_stream_out_0_ready),
    .io_stream_out_0_valid(splitters_6_io_stream_out_0_valid),
    .io_stream_out_0_bits(splitters_6_io_stream_out_0_bits)
  );
  StreamSplitterBinaryTree splitters_7 ( // @[Stab.scala 230:46]
    .io_stream_in_ready(splitters_7_io_stream_in_ready),
    .io_stream_in_valid(splitters_7_io_stream_in_valid),
    .io_stream_in_bits(splitters_7_io_stream_in_bits),
    .io_stream_out_0_ready(splitters_7_io_stream_out_0_ready),
    .io_stream_out_0_valid(splitters_7_io_stream_out_0_valid),
    .io_stream_out_0_bits(splitters_7_io_stream_out_0_bits)
  );
  StreamSplitterBinaryTree splitters_8 ( // @[Stab.scala 230:46]
    .io_stream_in_ready(splitters_8_io_stream_in_ready),
    .io_stream_in_valid(splitters_8_io_stream_in_valid),
    .io_stream_in_bits(splitters_8_io_stream_in_bits),
    .io_stream_out_0_ready(splitters_8_io_stream_out_0_ready),
    .io_stream_out_0_valid(splitters_8_io_stream_out_0_valid),
    .io_stream_out_0_bits(splitters_8_io_stream_out_0_bits)
  );
  StreamSplitterBinaryTree splitters_9 ( // @[Stab.scala 230:46]
    .io_stream_in_ready(splitters_9_io_stream_in_ready),
    .io_stream_in_valid(splitters_9_io_stream_in_valid),
    .io_stream_in_bits(splitters_9_io_stream_in_bits),
    .io_stream_out_0_ready(splitters_9_io_stream_out_0_ready),
    .io_stream_out_0_valid(splitters_9_io_stream_out_0_valid),
    .io_stream_out_0_bits(splitters_9_io_stream_out_0_bits)
  );
  StreamSplitterBinaryTree splitters_10 ( // @[Stab.scala 230:46]
    .io_stream_in_ready(splitters_10_io_stream_in_ready),
    .io_stream_in_valid(splitters_10_io_stream_in_valid),
    .io_stream_in_bits(splitters_10_io_stream_in_bits),
    .io_stream_out_0_ready(splitters_10_io_stream_out_0_ready),
    .io_stream_out_0_valid(splitters_10_io_stream_out_0_valid),
    .io_stream_out_0_bits(splitters_10_io_stream_out_0_bits)
  );
  StreamSplitterBinaryTree splitters_11 ( // @[Stab.scala 230:46]
    .io_stream_in_ready(splitters_11_io_stream_in_ready),
    .io_stream_in_valid(splitters_11_io_stream_in_valid),
    .io_stream_in_bits(splitters_11_io_stream_in_bits),
    .io_stream_out_0_ready(splitters_11_io_stream_out_0_ready),
    .io_stream_out_0_valid(splitters_11_io_stream_out_0_valid),
    .io_stream_out_0_bits(splitters_11_io_stream_out_0_bits)
  );
  StreamSplitterBinaryTree splitters_12 ( // @[Stab.scala 230:46]
    .io_stream_in_ready(splitters_12_io_stream_in_ready),
    .io_stream_in_valid(splitters_12_io_stream_in_valid),
    .io_stream_in_bits(splitters_12_io_stream_in_bits),
    .io_stream_out_0_ready(splitters_12_io_stream_out_0_ready),
    .io_stream_out_0_valid(splitters_12_io_stream_out_0_valid),
    .io_stream_out_0_bits(splitters_12_io_stream_out_0_bits)
  );
  StreamSplitterBinaryTree splitters_13 ( // @[Stab.scala 230:46]
    .io_stream_in_ready(splitters_13_io_stream_in_ready),
    .io_stream_in_valid(splitters_13_io_stream_in_valid),
    .io_stream_in_bits(splitters_13_io_stream_in_bits),
    .io_stream_out_0_ready(splitters_13_io_stream_out_0_ready),
    .io_stream_out_0_valid(splitters_13_io_stream_out_0_valid),
    .io_stream_out_0_bits(splitters_13_io_stream_out_0_bits)
  );
  StreamSplitterBinaryTree splitters_14 ( // @[Stab.scala 230:46]
    .io_stream_in_ready(splitters_14_io_stream_in_ready),
    .io_stream_in_valid(splitters_14_io_stream_in_valid),
    .io_stream_in_bits(splitters_14_io_stream_in_bits),
    .io_stream_out_0_ready(splitters_14_io_stream_out_0_ready),
    .io_stream_out_0_valid(splitters_14_io_stream_out_0_valid),
    .io_stream_out_0_bits(splitters_14_io_stream_out_0_bits)
  );
  StreamSplitterBinaryTree splitters_15 ( // @[Stab.scala 230:46]
    .io_stream_in_ready(splitters_15_io_stream_in_ready),
    .io_stream_in_valid(splitters_15_io_stream_in_valid),
    .io_stream_in_bits(splitters_15_io_stream_in_bits),
    .io_stream_out_0_ready(splitters_15_io_stream_out_0_ready),
    .io_stream_out_0_valid(splitters_15_io_stream_out_0_valid),
    .io_stream_out_0_bits(splitters_15_io_stream_out_0_bits)
  );
  assign io_stream_in_ready = turn_wrap_wrap ? splitters_15_io_stream_in_ready : _GEN_16; // @[Stab.scala 240:25 241:26]
  assign io_stream_out_0_valid = splitters_0_io_stream_out_0_valid; // @[Stab.scala 234:17]
  assign io_stream_out_0_bits = splitters_0_io_stream_out_0_bits; // @[Stab.scala 234:17]
  assign io_stream_out_1_valid = splitters_1_io_stream_out_0_valid; // @[Stab.scala 234:17]
  assign io_stream_out_1_bits = splitters_1_io_stream_out_0_bits; // @[Stab.scala 234:17]
  assign io_stream_out_2_valid = splitters_2_io_stream_out_0_valid; // @[Stab.scala 234:17]
  assign io_stream_out_2_bits = splitters_2_io_stream_out_0_bits; // @[Stab.scala 234:17]
  assign io_stream_out_3_valid = splitters_3_io_stream_out_0_valid; // @[Stab.scala 234:17]
  assign io_stream_out_3_bits = splitters_3_io_stream_out_0_bits; // @[Stab.scala 234:17]
  assign io_stream_out_4_valid = splitters_4_io_stream_out_0_valid; // @[Stab.scala 234:17]
  assign io_stream_out_4_bits = splitters_4_io_stream_out_0_bits; // @[Stab.scala 234:17]
  assign io_stream_out_5_valid = splitters_5_io_stream_out_0_valid; // @[Stab.scala 234:17]
  assign io_stream_out_5_bits = splitters_5_io_stream_out_0_bits; // @[Stab.scala 234:17]
  assign io_stream_out_6_valid = splitters_6_io_stream_out_0_valid; // @[Stab.scala 234:17]
  assign io_stream_out_6_bits = splitters_6_io_stream_out_0_bits; // @[Stab.scala 234:17]
  assign io_stream_out_7_valid = splitters_7_io_stream_out_0_valid; // @[Stab.scala 234:17]
  assign io_stream_out_7_bits = splitters_7_io_stream_out_0_bits; // @[Stab.scala 234:17]
  assign io_stream_out_8_valid = splitters_8_io_stream_out_0_valid; // @[Stab.scala 234:17]
  assign io_stream_out_8_bits = splitters_8_io_stream_out_0_bits; // @[Stab.scala 234:17]
  assign io_stream_out_9_valid = splitters_9_io_stream_out_0_valid; // @[Stab.scala 234:17]
  assign io_stream_out_9_bits = splitters_9_io_stream_out_0_bits; // @[Stab.scala 234:17]
  assign io_stream_out_10_valid = splitters_10_io_stream_out_0_valid; // @[Stab.scala 234:17]
  assign io_stream_out_10_bits = splitters_10_io_stream_out_0_bits; // @[Stab.scala 234:17]
  assign io_stream_out_11_valid = splitters_11_io_stream_out_0_valid; // @[Stab.scala 234:17]
  assign io_stream_out_11_bits = splitters_11_io_stream_out_0_bits; // @[Stab.scala 234:17]
  assign io_stream_out_12_valid = splitters_12_io_stream_out_0_valid; // @[Stab.scala 234:17]
  assign io_stream_out_12_bits = splitters_12_io_stream_out_0_bits; // @[Stab.scala 234:17]
  assign io_stream_out_13_valid = splitters_13_io_stream_out_0_valid; // @[Stab.scala 234:17]
  assign io_stream_out_13_bits = splitters_13_io_stream_out_0_bits; // @[Stab.scala 234:17]
  assign io_stream_out_14_valid = splitters_14_io_stream_out_0_valid; // @[Stab.scala 234:17]
  assign io_stream_out_14_bits = splitters_14_io_stream_out_0_bits; // @[Stab.scala 234:17]
  assign io_stream_out_15_valid = splitters_15_io_stream_out_0_valid; // @[Stab.scala 234:17]
  assign io_stream_out_15_bits = splitters_15_io_stream_out_0_bits; // @[Stab.scala 234:17]
  assign splitters_0_io_stream_in_valid = turn == 4'h0 & io_stream_in_valid; // @[Stab.scala 238:35]
  assign splitters_0_io_stream_in_bits = io_stream_in_bits; // @[Stab.scala 239:29]
  assign splitters_0_io_stream_out_0_ready = io_stream_out_0_ready; // @[Stab.scala 234:17]
  assign splitters_1_io_stream_in_valid = turn == 4'h1 & io_stream_in_valid; // @[Stab.scala 238:35]
  assign splitters_1_io_stream_in_bits = io_stream_in_bits; // @[Stab.scala 239:29]
  assign splitters_1_io_stream_out_0_ready = io_stream_out_1_ready; // @[Stab.scala 234:17]
  assign splitters_2_io_stream_in_valid = turn == 4'h2 & io_stream_in_valid; // @[Stab.scala 238:35]
  assign splitters_2_io_stream_in_bits = io_stream_in_bits; // @[Stab.scala 239:29]
  assign splitters_2_io_stream_out_0_ready = io_stream_out_2_ready; // @[Stab.scala 234:17]
  assign splitters_3_io_stream_in_valid = turn == 4'h3 & io_stream_in_valid; // @[Stab.scala 238:35]
  assign splitters_3_io_stream_in_bits = io_stream_in_bits; // @[Stab.scala 239:29]
  assign splitters_3_io_stream_out_0_ready = io_stream_out_3_ready; // @[Stab.scala 234:17]
  assign splitters_4_io_stream_in_valid = turn == 4'h4 & io_stream_in_valid; // @[Stab.scala 238:35]
  assign splitters_4_io_stream_in_bits = io_stream_in_bits; // @[Stab.scala 239:29]
  assign splitters_4_io_stream_out_0_ready = io_stream_out_4_ready; // @[Stab.scala 234:17]
  assign splitters_5_io_stream_in_valid = turn == 4'h5 & io_stream_in_valid; // @[Stab.scala 238:35]
  assign splitters_5_io_stream_in_bits = io_stream_in_bits; // @[Stab.scala 239:29]
  assign splitters_5_io_stream_out_0_ready = io_stream_out_5_ready; // @[Stab.scala 234:17]
  assign splitters_6_io_stream_in_valid = turn == 4'h6 & io_stream_in_valid; // @[Stab.scala 238:35]
  assign splitters_6_io_stream_in_bits = io_stream_in_bits; // @[Stab.scala 239:29]
  assign splitters_6_io_stream_out_0_ready = io_stream_out_6_ready; // @[Stab.scala 234:17]
  assign splitters_7_io_stream_in_valid = turn == 4'h7 & io_stream_in_valid; // @[Stab.scala 238:35]
  assign splitters_7_io_stream_in_bits = io_stream_in_bits; // @[Stab.scala 239:29]
  assign splitters_7_io_stream_out_0_ready = io_stream_out_7_ready; // @[Stab.scala 234:17]
  assign splitters_8_io_stream_in_valid = turn == 4'h8 & io_stream_in_valid; // @[Stab.scala 238:35]
  assign splitters_8_io_stream_in_bits = io_stream_in_bits; // @[Stab.scala 239:29]
  assign splitters_8_io_stream_out_0_ready = io_stream_out_8_ready; // @[Stab.scala 234:17]
  assign splitters_9_io_stream_in_valid = turn == 4'h9 & io_stream_in_valid; // @[Stab.scala 238:35]
  assign splitters_9_io_stream_in_bits = io_stream_in_bits; // @[Stab.scala 239:29]
  assign splitters_9_io_stream_out_0_ready = io_stream_out_9_ready; // @[Stab.scala 234:17]
  assign splitters_10_io_stream_in_valid = turn == 4'ha & io_stream_in_valid; // @[Stab.scala 238:35]
  assign splitters_10_io_stream_in_bits = io_stream_in_bits; // @[Stab.scala 239:29]
  assign splitters_10_io_stream_out_0_ready = io_stream_out_10_ready; // @[Stab.scala 234:17]
  assign splitters_11_io_stream_in_valid = turn == 4'hb & io_stream_in_valid; // @[Stab.scala 238:35]
  assign splitters_11_io_stream_in_bits = io_stream_in_bits; // @[Stab.scala 239:29]
  assign splitters_11_io_stream_out_0_ready = io_stream_out_11_ready; // @[Stab.scala 234:17]
  assign splitters_12_io_stream_in_valid = turn == 4'hc & io_stream_in_valid; // @[Stab.scala 238:35]
  assign splitters_12_io_stream_in_bits = io_stream_in_bits; // @[Stab.scala 239:29]
  assign splitters_12_io_stream_out_0_ready = io_stream_out_12_ready; // @[Stab.scala 234:17]
  assign splitters_13_io_stream_in_valid = turn == 4'hd & io_stream_in_valid; // @[Stab.scala 238:35]
  assign splitters_13_io_stream_in_bits = io_stream_in_bits; // @[Stab.scala 239:29]
  assign splitters_13_io_stream_out_0_ready = io_stream_out_13_ready; // @[Stab.scala 234:17]
  assign splitters_14_io_stream_in_valid = turn == 4'he & io_stream_in_valid; // @[Stab.scala 238:35]
  assign splitters_14_io_stream_in_bits = io_stream_in_bits; // @[Stab.scala 239:29]
  assign splitters_14_io_stream_out_0_ready = io_stream_out_14_ready; // @[Stab.scala 234:17]
  assign splitters_15_io_stream_in_valid = turn_wrap_wrap & io_stream_in_valid; // @[Stab.scala 238:35]
  assign splitters_15_io_stream_in_bits = io_stream_in_bits; // @[Stab.scala 239:29]
  assign splitters_15_io_stream_out_0_ready = io_stream_out_15_ready; // @[Stab.scala 234:17]
  always @(posedge clock) begin
    if (reset) begin // @[Counter.scala 62:40]
      turn <= 4'h0; // @[Counter.scala 62:40]
    end else if (_turn_T) begin // @[Counter.scala 120:16]
      turn <= _turn_wrap_value_T_1; // @[Counter.scala 78:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  turn = _RAND_0[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  wrap1 = ~use2 & _T_1; // @[Stab.scala 142:41]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_2 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_3 = _T & wrap1 | _GEN_2; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_3;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_1(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg  counter1; // @[Counter.scala 62:40]
  wire  wrap1 = _T_2 & counter1; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_3 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_4 = _T & wrap1 | _GEN_3; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_4;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 1'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      counter1 <= counter1 + 1'h1; // @[Counter.scala 78:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_2(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [1:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 2'h2; // @[Counter.scala 74:24]
  wire [1:0] _wrap_value_T_1 = counter1 + 2'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 2'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 2'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_3(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [1:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 2'h3; // @[Counter.scala 74:24]
  wire [1:0] _wrap_value_T_1 = counter1 + 2'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_3 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_4 = _T & wrap1 | _GEN_3; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_4;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 2'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_4(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [2:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 3'h4; // @[Counter.scala 74:24]
  wire [2:0] _wrap_value_T_1 = counter1 + 3'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 3'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 3'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_5(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [2:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 3'h5; // @[Counter.scala 74:24]
  wire [2:0] _wrap_value_T_1 = counter1 + 3'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 3'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 3'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_6(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [2:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 3'h6; // @[Counter.scala 74:24]
  wire [2:0] _wrap_value_T_1 = counter1 + 3'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 3'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 3'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_7(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [2:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 3'h7; // @[Counter.scala 74:24]
  wire [2:0] _wrap_value_T_1 = counter1 + 3'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_3 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_4 = _T & wrap1 | _GEN_3; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_4;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 3'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_8(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [3:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 4'h8; // @[Counter.scala 74:24]
  wire [3:0] _wrap_value_T_1 = counter1 + 4'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 4'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 4'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_9(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [3:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 4'h9; // @[Counter.scala 74:24]
  wire [3:0] _wrap_value_T_1 = counter1 + 4'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 4'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 4'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_10(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [3:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 4'ha; // @[Counter.scala 74:24]
  wire [3:0] _wrap_value_T_1 = counter1 + 4'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 4'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 4'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_11(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [3:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 4'hb; // @[Counter.scala 74:24]
  wire [3:0] _wrap_value_T_1 = counter1 + 4'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 4'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 4'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_12(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [3:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 4'hc; // @[Counter.scala 74:24]
  wire [3:0] _wrap_value_T_1 = counter1 + 4'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 4'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 4'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_13(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [3:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 4'hd; // @[Counter.scala 74:24]
  wire [3:0] _wrap_value_T_1 = counter1 + 4'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 4'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 4'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_14(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [3:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 4'he; // @[Counter.scala 74:24]
  wire [3:0] _wrap_value_T_1 = counter1 + 4'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 4'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 4'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_15(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [3:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 4'hf; // @[Counter.scala 74:24]
  wire [3:0] _wrap_value_T_1 = counter1 + 4'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_3 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_4 = _T & wrap1 | _GEN_3; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_4;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 4'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_16(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [4:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 5'h10; // @[Counter.scala 74:24]
  wire [4:0] _wrap_value_T_1 = counter1 + 5'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 5'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_17(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [4:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 5'h11; // @[Counter.scala 74:24]
  wire [4:0] _wrap_value_T_1 = counter1 + 5'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 5'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_18(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [4:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 5'h12; // @[Counter.scala 74:24]
  wire [4:0] _wrap_value_T_1 = counter1 + 5'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 5'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_19(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [4:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 5'h13; // @[Counter.scala 74:24]
  wire [4:0] _wrap_value_T_1 = counter1 + 5'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 5'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_20(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [4:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 5'h14; // @[Counter.scala 74:24]
  wire [4:0] _wrap_value_T_1 = counter1 + 5'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 5'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_21(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [4:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 5'h15; // @[Counter.scala 74:24]
  wire [4:0] _wrap_value_T_1 = counter1 + 5'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 5'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_22(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [4:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 5'h16; // @[Counter.scala 74:24]
  wire [4:0] _wrap_value_T_1 = counter1 + 5'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 5'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_23(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [4:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 5'h17; // @[Counter.scala 74:24]
  wire [4:0] _wrap_value_T_1 = counter1 + 5'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 5'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_24(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [4:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 5'h18; // @[Counter.scala 74:24]
  wire [4:0] _wrap_value_T_1 = counter1 + 5'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 5'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_25(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [4:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 5'h19; // @[Counter.scala 74:24]
  wire [4:0] _wrap_value_T_1 = counter1 + 5'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 5'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_26(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [4:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 5'h1a; // @[Counter.scala 74:24]
  wire [4:0] _wrap_value_T_1 = counter1 + 5'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 5'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_27(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [4:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 5'h1b; // @[Counter.scala 74:24]
  wire [4:0] _wrap_value_T_1 = counter1 + 5'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 5'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_28(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [4:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 5'h1c; // @[Counter.scala 74:24]
  wire [4:0] _wrap_value_T_1 = counter1 + 5'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 5'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_29(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [4:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 5'h1d; // @[Counter.scala 74:24]
  wire [4:0] _wrap_value_T_1 = counter1 + 5'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 5'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_30(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [4:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 5'h1e; // @[Counter.scala 74:24]
  wire [4:0] _wrap_value_T_1 = counter1 + 5'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 5'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_31(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [4:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 5'h1f; // @[Counter.scala 74:24]
  wire [4:0] _wrap_value_T_1 = counter1 + 5'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_3 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_4 = _T & wrap1 | _GEN_3; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_4;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 5'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_32(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h20; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_33(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h21; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_34(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h22; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_35(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h23; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_36(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h24; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_37(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h25; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_38(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h26; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_39(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h27; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_40(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h28; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_41(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h29; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_42(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h2a; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_43(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h2b; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_44(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h2c; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_45(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h2d; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_46(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h2e; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_47(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h2f; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_48(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h30; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_49(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h31; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_50(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h32; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_51(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h33; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_52(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h34; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_53(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h35; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_54(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h36; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_55(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h37; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_56(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h38; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_57(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h39; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_58(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h3a; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_59(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h3b; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_60(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h3c; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_61(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h3d; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_62(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h3e; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 6'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_63(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [5:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 6'h3f; // @[Counter.scala 74:24]
  wire [5:0] _wrap_value_T_1 = counter1 + 6'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_3 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_4 = _T & wrap1 | _GEN_3; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_4;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 6'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_64(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h40; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_65(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h41; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_66(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h42; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_67(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h43; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_68(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h44; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_69(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h45; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_70(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h46; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_71(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h47; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_72(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h48; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_73(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h49; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_74(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h4a; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_75(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h4b; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_76(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h4c; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_77(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h4d; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_78(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h4e; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_79(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h4f; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_80(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h50; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_81(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h51; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_82(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h52; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_83(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h53; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_84(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h54; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_85(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h55; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_86(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h56; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_87(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h57; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_88(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h58; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_89(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h59; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_90(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h5a; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_91(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h5b; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_92(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h5c; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_93(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h5d; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_94(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h5e; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_95(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h5f; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_96(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h60; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_97(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h61; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_98(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h62; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_99(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h63; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_100(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h64; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_101(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h65; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_102(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h66; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_103(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h67; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_104(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h68; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_105(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h69; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_106(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h6a; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_107(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h6b; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_108(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h6c; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_109(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h6d; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_110(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h6e; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_111(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h6f; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_112(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h70; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_113(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h71; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_114(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h72; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_115(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h73; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_116(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h74; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_117(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h75; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_118(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h76; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_119(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h77; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_120(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h78; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_121(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h79; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_122(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h7a; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_123(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h7b; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_124(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h7c; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_125(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h7d; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_126(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h7e; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 7'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_127(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [6:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 7'h7f; // @[Counter.scala 74:24]
  wire [6:0] _wrap_value_T_1 = counter1 + 7'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_3 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_4 = _T & wrap1 | _GEN_3; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_4;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 7'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_128(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h80; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_129(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h81; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_130(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h82; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_131(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h83; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_132(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h84; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_133(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h85; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_134(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h86; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_135(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h87; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_136(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h88; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_137(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h89; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_138(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h8a; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_139(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h8b; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_140(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h8c; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_141(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h8d; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_142(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h8e; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_143(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h8f; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_144(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h90; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_145(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h91; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_146(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h92; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_147(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h93; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_148(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h94; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_149(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h95; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_150(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h96; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_151(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h97; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_152(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h98; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_153(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h99; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_154(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h9a; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_155(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h9b; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_156(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h9c; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_157(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h9d; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_158(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h9e; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_159(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'h9f; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_160(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'ha0; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_161(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'ha1; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_162(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'ha2; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_163(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'ha3; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_164(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'ha4; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_165(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'ha5; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_166(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'ha6; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_167(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'ha7; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_168(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'ha8; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_169(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'ha9; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_170(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'haa; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_171(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hab; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_172(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hac; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_173(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'had; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_174(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hae; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_175(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'haf; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_176(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hb0; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_177(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hb1; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_178(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hb2; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_179(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hb3; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_180(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hb4; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_181(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hb5; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_182(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hb6; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_183(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hb7; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_184(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hb8; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_185(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hb9; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_186(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hba; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_187(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hbb; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_188(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hbc; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_189(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hbd; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_190(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hbe; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_191(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hbf; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_192(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hc0; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_193(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hc1; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_194(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hc2; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_195(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hc3; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_196(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hc4; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_197(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hc5; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_198(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hc6; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_199(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hc7; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_200(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hc8; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_201(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hc9; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_202(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hca; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_203(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hcb; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_204(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hcc; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_205(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hcd; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_206(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hce; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_207(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hcf; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_208(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hd0; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_209(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hd1; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_210(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hd2; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_211(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hd3; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_212(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hd4; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_213(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hd5; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_214(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hd6; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_215(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hd7; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_216(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hd8; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_217(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hd9; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_218(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hda; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_219(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hdb; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_220(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hdc; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_221(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hdd; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_222(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hde; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_223(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hdf; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_224(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'he0; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_225(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'he1; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_226(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'he2; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_227(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'he3; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_228(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'he4; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_229(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'he5; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_230(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'he6; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_231(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'he7; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_232(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'he8; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_233(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'he9; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_234(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hea; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_235(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'heb; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_236(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hec; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_237(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hed; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_238(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hee; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_239(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hef; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_240(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hf0; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_241(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hf1; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_242(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hf2; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_243(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hf3; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_244(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hf4; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_245(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hf5; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_246(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hf6; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_247(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hf7; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_248(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hf8; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_249(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hf9; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_250(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hfa; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_251(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hfb; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_252(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hfc; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_253(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hfd; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMerger_254(
  input         clock,
  input         reset,
  output        io_stream1_ready,
  input         io_stream1_valid,
  input  [31:0] io_stream1_bits,
  output        io_stream2_ready,
  input         io_stream2_valid,
  input  [31:0] io_stream2_bits,
  input         io_result_ready,
  output        io_result_valid,
  output [31:0] io_result_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg  use2; // @[Stab.scala 141:34]
  wire  _T = ~use2; // @[Stab.scala 142:35]
  wire  _T_1 = io_result_ready & io_result_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = ~use2 & _T_1; // @[Stab.scala 142:41]
  reg [7:0] counter1; // @[Counter.scala 62:40]
  wire  wrap_wrap = counter1 == 8'hfe; // @[Counter.scala 74:24]
  wire [7:0] _wrap_value_T_1 = counter1 + 8'h1; // @[Counter.scala 78:24]
  wire  wrap1 = _T_2 & wrap_wrap; // @[Counter.scala 120:{16,23}]
  wire  wrap2 = use2 & _T_1; // @[Stab.scala 143:40]
  wire  _GEN_4 = use2 & wrap2 ? 1'h0 : use2; // @[Stab.scala 145:23 146:10 141:34]
  wire  _GEN_5 = _T & wrap1 | _GEN_4; // @[Stab.scala 149:24 150:10]
  assign io_stream1_ready = _T & io_result_ready; // @[Stab.scala 155:15 156:15 152:20]
  assign io_stream2_ready = _T ? 1'h0 : io_result_ready; // @[Stab.scala 155:15 153:20 158:15]
  assign io_result_valid = _T ? io_stream1_valid : io_stream2_valid; // @[Stab.scala 155:15 156:15 158:15]
  assign io_result_bits = _T ? io_stream1_bits : io_stream2_bits; // @[Stab.scala 155:15 156:15 158:15]
  always @(posedge clock) begin
    if (reset) begin // @[Stab.scala 141:34]
      use2 <= 1'h0; // @[Stab.scala 141:34]
    end else begin
      use2 <= _GEN_5;
    end
    if (reset) begin // @[Counter.scala 62:40]
      counter1 <= 8'h0; // @[Counter.scala 62:40]
    end else if (_T_2) begin // @[Counter.scala 120:16]
      if (wrap_wrap) begin // @[Counter.scala 88:20]
        counter1 <= 8'h0; // @[Counter.scala 88:28]
      end else begin
        counter1 <= _wrap_value_T_1; // @[Counter.scala 78:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  use2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  counter1 = _RAND_1[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module StreamMergerTree(
  input         clock,
  input         reset,
  output        io_stream_in_0_ready,
  input         io_stream_in_0_valid,
  input  [31:0] io_stream_in_0_bits,
  output        io_stream_in_1_ready,
  input         io_stream_in_1_valid,
  input  [31:0] io_stream_in_1_bits,
  output        io_stream_in_2_ready,
  input         io_stream_in_2_valid,
  input  [31:0] io_stream_in_2_bits,
  output        io_stream_in_3_ready,
  input         io_stream_in_3_valid,
  input  [31:0] io_stream_in_3_bits,
  output        io_stream_in_4_ready,
  input         io_stream_in_4_valid,
  input  [31:0] io_stream_in_4_bits,
  output        io_stream_in_5_ready,
  input         io_stream_in_5_valid,
  input  [31:0] io_stream_in_5_bits,
  output        io_stream_in_6_ready,
  input         io_stream_in_6_valid,
  input  [31:0] io_stream_in_6_bits,
  output        io_stream_in_7_ready,
  input         io_stream_in_7_valid,
  input  [31:0] io_stream_in_7_bits,
  output        io_stream_in_8_ready,
  input         io_stream_in_8_valid,
  input  [31:0] io_stream_in_8_bits,
  output        io_stream_in_9_ready,
  input         io_stream_in_9_valid,
  input  [31:0] io_stream_in_9_bits,
  output        io_stream_in_10_ready,
  input         io_stream_in_10_valid,
  input  [31:0] io_stream_in_10_bits,
  output        io_stream_in_11_ready,
  input         io_stream_in_11_valid,
  input  [31:0] io_stream_in_11_bits,
  output        io_stream_in_12_ready,
  input         io_stream_in_12_valid,
  input  [31:0] io_stream_in_12_bits,
  output        io_stream_in_13_ready,
  input         io_stream_in_13_valid,
  input  [31:0] io_stream_in_13_bits,
  output        io_stream_in_14_ready,
  input         io_stream_in_14_valid,
  input  [31:0] io_stream_in_14_bits,
  output        io_stream_in_15_ready,
  input         io_stream_in_15_valid,
  input  [31:0] io_stream_in_15_bits,
  output        io_stream_in_16_ready,
  input         io_stream_in_16_valid,
  input  [31:0] io_stream_in_16_bits,
  output        io_stream_in_17_ready,
  input         io_stream_in_17_valid,
  input  [31:0] io_stream_in_17_bits,
  output        io_stream_in_18_ready,
  input         io_stream_in_18_valid,
  input  [31:0] io_stream_in_18_bits,
  output        io_stream_in_19_ready,
  input         io_stream_in_19_valid,
  input  [31:0] io_stream_in_19_bits,
  output        io_stream_in_20_ready,
  input         io_stream_in_20_valid,
  input  [31:0] io_stream_in_20_bits,
  output        io_stream_in_21_ready,
  input         io_stream_in_21_valid,
  input  [31:0] io_stream_in_21_bits,
  output        io_stream_in_22_ready,
  input         io_stream_in_22_valid,
  input  [31:0] io_stream_in_22_bits,
  output        io_stream_in_23_ready,
  input         io_stream_in_23_valid,
  input  [31:0] io_stream_in_23_bits,
  output        io_stream_in_24_ready,
  input         io_stream_in_24_valid,
  input  [31:0] io_stream_in_24_bits,
  output        io_stream_in_25_ready,
  input         io_stream_in_25_valid,
  input  [31:0] io_stream_in_25_bits,
  output        io_stream_in_26_ready,
  input         io_stream_in_26_valid,
  input  [31:0] io_stream_in_26_bits,
  output        io_stream_in_27_ready,
  input         io_stream_in_27_valid,
  input  [31:0] io_stream_in_27_bits,
  output        io_stream_in_28_ready,
  input         io_stream_in_28_valid,
  input  [31:0] io_stream_in_28_bits,
  output        io_stream_in_29_ready,
  input         io_stream_in_29_valid,
  input  [31:0] io_stream_in_29_bits,
  output        io_stream_in_30_ready,
  input         io_stream_in_30_valid,
  input  [31:0] io_stream_in_30_bits,
  output        io_stream_in_31_ready,
  input         io_stream_in_31_valid,
  input  [31:0] io_stream_in_31_bits,
  output        io_stream_in_32_ready,
  input         io_stream_in_32_valid,
  input  [31:0] io_stream_in_32_bits,
  output        io_stream_in_33_ready,
  input         io_stream_in_33_valid,
  input  [31:0] io_stream_in_33_bits,
  output        io_stream_in_34_ready,
  input         io_stream_in_34_valid,
  input  [31:0] io_stream_in_34_bits,
  output        io_stream_in_35_ready,
  input         io_stream_in_35_valid,
  input  [31:0] io_stream_in_35_bits,
  output        io_stream_in_36_ready,
  input         io_stream_in_36_valid,
  input  [31:0] io_stream_in_36_bits,
  output        io_stream_in_37_ready,
  input         io_stream_in_37_valid,
  input  [31:0] io_stream_in_37_bits,
  output        io_stream_in_38_ready,
  input         io_stream_in_38_valid,
  input  [31:0] io_stream_in_38_bits,
  output        io_stream_in_39_ready,
  input         io_stream_in_39_valid,
  input  [31:0] io_stream_in_39_bits,
  output        io_stream_in_40_ready,
  input         io_stream_in_40_valid,
  input  [31:0] io_stream_in_40_bits,
  output        io_stream_in_41_ready,
  input         io_stream_in_41_valid,
  input  [31:0] io_stream_in_41_bits,
  output        io_stream_in_42_ready,
  input         io_stream_in_42_valid,
  input  [31:0] io_stream_in_42_bits,
  output        io_stream_in_43_ready,
  input         io_stream_in_43_valid,
  input  [31:0] io_stream_in_43_bits,
  output        io_stream_in_44_ready,
  input         io_stream_in_44_valid,
  input  [31:0] io_stream_in_44_bits,
  output        io_stream_in_45_ready,
  input         io_stream_in_45_valid,
  input  [31:0] io_stream_in_45_bits,
  output        io_stream_in_46_ready,
  input         io_stream_in_46_valid,
  input  [31:0] io_stream_in_46_bits,
  output        io_stream_in_47_ready,
  input         io_stream_in_47_valid,
  input  [31:0] io_stream_in_47_bits,
  output        io_stream_in_48_ready,
  input         io_stream_in_48_valid,
  input  [31:0] io_stream_in_48_bits,
  output        io_stream_in_49_ready,
  input         io_stream_in_49_valid,
  input  [31:0] io_stream_in_49_bits,
  output        io_stream_in_50_ready,
  input         io_stream_in_50_valid,
  input  [31:0] io_stream_in_50_bits,
  output        io_stream_in_51_ready,
  input         io_stream_in_51_valid,
  input  [31:0] io_stream_in_51_bits,
  output        io_stream_in_52_ready,
  input         io_stream_in_52_valid,
  input  [31:0] io_stream_in_52_bits,
  output        io_stream_in_53_ready,
  input         io_stream_in_53_valid,
  input  [31:0] io_stream_in_53_bits,
  output        io_stream_in_54_ready,
  input         io_stream_in_54_valid,
  input  [31:0] io_stream_in_54_bits,
  output        io_stream_in_55_ready,
  input         io_stream_in_55_valid,
  input  [31:0] io_stream_in_55_bits,
  output        io_stream_in_56_ready,
  input         io_stream_in_56_valid,
  input  [31:0] io_stream_in_56_bits,
  output        io_stream_in_57_ready,
  input         io_stream_in_57_valid,
  input  [31:0] io_stream_in_57_bits,
  output        io_stream_in_58_ready,
  input         io_stream_in_58_valid,
  input  [31:0] io_stream_in_58_bits,
  output        io_stream_in_59_ready,
  input         io_stream_in_59_valid,
  input  [31:0] io_stream_in_59_bits,
  output        io_stream_in_60_ready,
  input         io_stream_in_60_valid,
  input  [31:0] io_stream_in_60_bits,
  output        io_stream_in_61_ready,
  input         io_stream_in_61_valid,
  input  [31:0] io_stream_in_61_bits,
  output        io_stream_in_62_ready,
  input         io_stream_in_62_valid,
  input  [31:0] io_stream_in_62_bits,
  output        io_stream_in_63_ready,
  input         io_stream_in_63_valid,
  input  [31:0] io_stream_in_63_bits,
  output        io_stream_in_64_ready,
  input         io_stream_in_64_valid,
  input  [31:0] io_stream_in_64_bits,
  output        io_stream_in_65_ready,
  input         io_stream_in_65_valid,
  input  [31:0] io_stream_in_65_bits,
  output        io_stream_in_66_ready,
  input         io_stream_in_66_valid,
  input  [31:0] io_stream_in_66_bits,
  output        io_stream_in_67_ready,
  input         io_stream_in_67_valid,
  input  [31:0] io_stream_in_67_bits,
  output        io_stream_in_68_ready,
  input         io_stream_in_68_valid,
  input  [31:0] io_stream_in_68_bits,
  output        io_stream_in_69_ready,
  input         io_stream_in_69_valid,
  input  [31:0] io_stream_in_69_bits,
  output        io_stream_in_70_ready,
  input         io_stream_in_70_valid,
  input  [31:0] io_stream_in_70_bits,
  output        io_stream_in_71_ready,
  input         io_stream_in_71_valid,
  input  [31:0] io_stream_in_71_bits,
  output        io_stream_in_72_ready,
  input         io_stream_in_72_valid,
  input  [31:0] io_stream_in_72_bits,
  output        io_stream_in_73_ready,
  input         io_stream_in_73_valid,
  input  [31:0] io_stream_in_73_bits,
  output        io_stream_in_74_ready,
  input         io_stream_in_74_valid,
  input  [31:0] io_stream_in_74_bits,
  output        io_stream_in_75_ready,
  input         io_stream_in_75_valid,
  input  [31:0] io_stream_in_75_bits,
  output        io_stream_in_76_ready,
  input         io_stream_in_76_valid,
  input  [31:0] io_stream_in_76_bits,
  output        io_stream_in_77_ready,
  input         io_stream_in_77_valid,
  input  [31:0] io_stream_in_77_bits,
  output        io_stream_in_78_ready,
  input         io_stream_in_78_valid,
  input  [31:0] io_stream_in_78_bits,
  output        io_stream_in_79_ready,
  input         io_stream_in_79_valid,
  input  [31:0] io_stream_in_79_bits,
  output        io_stream_in_80_ready,
  input         io_stream_in_80_valid,
  input  [31:0] io_stream_in_80_bits,
  output        io_stream_in_81_ready,
  input         io_stream_in_81_valid,
  input  [31:0] io_stream_in_81_bits,
  output        io_stream_in_82_ready,
  input         io_stream_in_82_valid,
  input  [31:0] io_stream_in_82_bits,
  output        io_stream_in_83_ready,
  input         io_stream_in_83_valid,
  input  [31:0] io_stream_in_83_bits,
  output        io_stream_in_84_ready,
  input         io_stream_in_84_valid,
  input  [31:0] io_stream_in_84_bits,
  output        io_stream_in_85_ready,
  input         io_stream_in_85_valid,
  input  [31:0] io_stream_in_85_bits,
  output        io_stream_in_86_ready,
  input         io_stream_in_86_valid,
  input  [31:0] io_stream_in_86_bits,
  output        io_stream_in_87_ready,
  input         io_stream_in_87_valid,
  input  [31:0] io_stream_in_87_bits,
  output        io_stream_in_88_ready,
  input         io_stream_in_88_valid,
  input  [31:0] io_stream_in_88_bits,
  output        io_stream_in_89_ready,
  input         io_stream_in_89_valid,
  input  [31:0] io_stream_in_89_bits,
  output        io_stream_in_90_ready,
  input         io_stream_in_90_valid,
  input  [31:0] io_stream_in_90_bits,
  output        io_stream_in_91_ready,
  input         io_stream_in_91_valid,
  input  [31:0] io_stream_in_91_bits,
  output        io_stream_in_92_ready,
  input         io_stream_in_92_valid,
  input  [31:0] io_stream_in_92_bits,
  output        io_stream_in_93_ready,
  input         io_stream_in_93_valid,
  input  [31:0] io_stream_in_93_bits,
  output        io_stream_in_94_ready,
  input         io_stream_in_94_valid,
  input  [31:0] io_stream_in_94_bits,
  output        io_stream_in_95_ready,
  input         io_stream_in_95_valid,
  input  [31:0] io_stream_in_95_bits,
  output        io_stream_in_96_ready,
  input         io_stream_in_96_valid,
  input  [31:0] io_stream_in_96_bits,
  output        io_stream_in_97_ready,
  input         io_stream_in_97_valid,
  input  [31:0] io_stream_in_97_bits,
  output        io_stream_in_98_ready,
  input         io_stream_in_98_valid,
  input  [31:0] io_stream_in_98_bits,
  output        io_stream_in_99_ready,
  input         io_stream_in_99_valid,
  input  [31:0] io_stream_in_99_bits,
  output        io_stream_in_100_ready,
  input         io_stream_in_100_valid,
  input  [31:0] io_stream_in_100_bits,
  output        io_stream_in_101_ready,
  input         io_stream_in_101_valid,
  input  [31:0] io_stream_in_101_bits,
  output        io_stream_in_102_ready,
  input         io_stream_in_102_valid,
  input  [31:0] io_stream_in_102_bits,
  output        io_stream_in_103_ready,
  input         io_stream_in_103_valid,
  input  [31:0] io_stream_in_103_bits,
  output        io_stream_in_104_ready,
  input         io_stream_in_104_valid,
  input  [31:0] io_stream_in_104_bits,
  output        io_stream_in_105_ready,
  input         io_stream_in_105_valid,
  input  [31:0] io_stream_in_105_bits,
  output        io_stream_in_106_ready,
  input         io_stream_in_106_valid,
  input  [31:0] io_stream_in_106_bits,
  output        io_stream_in_107_ready,
  input         io_stream_in_107_valid,
  input  [31:0] io_stream_in_107_bits,
  output        io_stream_in_108_ready,
  input         io_stream_in_108_valid,
  input  [31:0] io_stream_in_108_bits,
  output        io_stream_in_109_ready,
  input         io_stream_in_109_valid,
  input  [31:0] io_stream_in_109_bits,
  output        io_stream_in_110_ready,
  input         io_stream_in_110_valid,
  input  [31:0] io_stream_in_110_bits,
  output        io_stream_in_111_ready,
  input         io_stream_in_111_valid,
  input  [31:0] io_stream_in_111_bits,
  output        io_stream_in_112_ready,
  input         io_stream_in_112_valid,
  input  [31:0] io_stream_in_112_bits,
  output        io_stream_in_113_ready,
  input         io_stream_in_113_valid,
  input  [31:0] io_stream_in_113_bits,
  output        io_stream_in_114_ready,
  input         io_stream_in_114_valid,
  input  [31:0] io_stream_in_114_bits,
  output        io_stream_in_115_ready,
  input         io_stream_in_115_valid,
  input  [31:0] io_stream_in_115_bits,
  output        io_stream_in_116_ready,
  input         io_stream_in_116_valid,
  input  [31:0] io_stream_in_116_bits,
  output        io_stream_in_117_ready,
  input         io_stream_in_117_valid,
  input  [31:0] io_stream_in_117_bits,
  output        io_stream_in_118_ready,
  input         io_stream_in_118_valid,
  input  [31:0] io_stream_in_118_bits,
  output        io_stream_in_119_ready,
  input         io_stream_in_119_valid,
  input  [31:0] io_stream_in_119_bits,
  output        io_stream_in_120_ready,
  input         io_stream_in_120_valid,
  input  [31:0] io_stream_in_120_bits,
  output        io_stream_in_121_ready,
  input         io_stream_in_121_valid,
  input  [31:0] io_stream_in_121_bits,
  output        io_stream_in_122_ready,
  input         io_stream_in_122_valid,
  input  [31:0] io_stream_in_122_bits,
  output        io_stream_in_123_ready,
  input         io_stream_in_123_valid,
  input  [31:0] io_stream_in_123_bits,
  output        io_stream_in_124_ready,
  input         io_stream_in_124_valid,
  input  [31:0] io_stream_in_124_bits,
  output        io_stream_in_125_ready,
  input         io_stream_in_125_valid,
  input  [31:0] io_stream_in_125_bits,
  output        io_stream_in_126_ready,
  input         io_stream_in_126_valid,
  input  [31:0] io_stream_in_126_bits,
  output        io_stream_in_127_ready,
  input         io_stream_in_127_valid,
  input  [31:0] io_stream_in_127_bits,
  output        io_stream_in_128_ready,
  input         io_stream_in_128_valid,
  input  [31:0] io_stream_in_128_bits,
  output        io_stream_in_129_ready,
  input         io_stream_in_129_valid,
  input  [31:0] io_stream_in_129_bits,
  output        io_stream_in_130_ready,
  input         io_stream_in_130_valid,
  input  [31:0] io_stream_in_130_bits,
  output        io_stream_in_131_ready,
  input         io_stream_in_131_valid,
  input  [31:0] io_stream_in_131_bits,
  output        io_stream_in_132_ready,
  input         io_stream_in_132_valid,
  input  [31:0] io_stream_in_132_bits,
  output        io_stream_in_133_ready,
  input         io_stream_in_133_valid,
  input  [31:0] io_stream_in_133_bits,
  output        io_stream_in_134_ready,
  input         io_stream_in_134_valid,
  input  [31:0] io_stream_in_134_bits,
  output        io_stream_in_135_ready,
  input         io_stream_in_135_valid,
  input  [31:0] io_stream_in_135_bits,
  output        io_stream_in_136_ready,
  input         io_stream_in_136_valid,
  input  [31:0] io_stream_in_136_bits,
  output        io_stream_in_137_ready,
  input         io_stream_in_137_valid,
  input  [31:0] io_stream_in_137_bits,
  output        io_stream_in_138_ready,
  input         io_stream_in_138_valid,
  input  [31:0] io_stream_in_138_bits,
  output        io_stream_in_139_ready,
  input         io_stream_in_139_valid,
  input  [31:0] io_stream_in_139_bits,
  output        io_stream_in_140_ready,
  input         io_stream_in_140_valid,
  input  [31:0] io_stream_in_140_bits,
  output        io_stream_in_141_ready,
  input         io_stream_in_141_valid,
  input  [31:0] io_stream_in_141_bits,
  output        io_stream_in_142_ready,
  input         io_stream_in_142_valid,
  input  [31:0] io_stream_in_142_bits,
  output        io_stream_in_143_ready,
  input         io_stream_in_143_valid,
  input  [31:0] io_stream_in_143_bits,
  output        io_stream_in_144_ready,
  input         io_stream_in_144_valid,
  input  [31:0] io_stream_in_144_bits,
  output        io_stream_in_145_ready,
  input         io_stream_in_145_valid,
  input  [31:0] io_stream_in_145_bits,
  output        io_stream_in_146_ready,
  input         io_stream_in_146_valid,
  input  [31:0] io_stream_in_146_bits,
  output        io_stream_in_147_ready,
  input         io_stream_in_147_valid,
  input  [31:0] io_stream_in_147_bits,
  output        io_stream_in_148_ready,
  input         io_stream_in_148_valid,
  input  [31:0] io_stream_in_148_bits,
  output        io_stream_in_149_ready,
  input         io_stream_in_149_valid,
  input  [31:0] io_stream_in_149_bits,
  output        io_stream_in_150_ready,
  input         io_stream_in_150_valid,
  input  [31:0] io_stream_in_150_bits,
  output        io_stream_in_151_ready,
  input         io_stream_in_151_valid,
  input  [31:0] io_stream_in_151_bits,
  output        io_stream_in_152_ready,
  input         io_stream_in_152_valid,
  input  [31:0] io_stream_in_152_bits,
  output        io_stream_in_153_ready,
  input         io_stream_in_153_valid,
  input  [31:0] io_stream_in_153_bits,
  output        io_stream_in_154_ready,
  input         io_stream_in_154_valid,
  input  [31:0] io_stream_in_154_bits,
  output        io_stream_in_155_ready,
  input         io_stream_in_155_valid,
  input  [31:0] io_stream_in_155_bits,
  output        io_stream_in_156_ready,
  input         io_stream_in_156_valid,
  input  [31:0] io_stream_in_156_bits,
  output        io_stream_in_157_ready,
  input         io_stream_in_157_valid,
  input  [31:0] io_stream_in_157_bits,
  output        io_stream_in_158_ready,
  input         io_stream_in_158_valid,
  input  [31:0] io_stream_in_158_bits,
  output        io_stream_in_159_ready,
  input         io_stream_in_159_valid,
  input  [31:0] io_stream_in_159_bits,
  output        io_stream_in_160_ready,
  input         io_stream_in_160_valid,
  input  [31:0] io_stream_in_160_bits,
  output        io_stream_in_161_ready,
  input         io_stream_in_161_valid,
  input  [31:0] io_stream_in_161_bits,
  output        io_stream_in_162_ready,
  input         io_stream_in_162_valid,
  input  [31:0] io_stream_in_162_bits,
  output        io_stream_in_163_ready,
  input         io_stream_in_163_valid,
  input  [31:0] io_stream_in_163_bits,
  output        io_stream_in_164_ready,
  input         io_stream_in_164_valid,
  input  [31:0] io_stream_in_164_bits,
  output        io_stream_in_165_ready,
  input         io_stream_in_165_valid,
  input  [31:0] io_stream_in_165_bits,
  output        io_stream_in_166_ready,
  input         io_stream_in_166_valid,
  input  [31:0] io_stream_in_166_bits,
  output        io_stream_in_167_ready,
  input         io_stream_in_167_valid,
  input  [31:0] io_stream_in_167_bits,
  output        io_stream_in_168_ready,
  input         io_stream_in_168_valid,
  input  [31:0] io_stream_in_168_bits,
  output        io_stream_in_169_ready,
  input         io_stream_in_169_valid,
  input  [31:0] io_stream_in_169_bits,
  output        io_stream_in_170_ready,
  input         io_stream_in_170_valid,
  input  [31:0] io_stream_in_170_bits,
  output        io_stream_in_171_ready,
  input         io_stream_in_171_valid,
  input  [31:0] io_stream_in_171_bits,
  output        io_stream_in_172_ready,
  input         io_stream_in_172_valid,
  input  [31:0] io_stream_in_172_bits,
  output        io_stream_in_173_ready,
  input         io_stream_in_173_valid,
  input  [31:0] io_stream_in_173_bits,
  output        io_stream_in_174_ready,
  input         io_stream_in_174_valid,
  input  [31:0] io_stream_in_174_bits,
  output        io_stream_in_175_ready,
  input         io_stream_in_175_valid,
  input  [31:0] io_stream_in_175_bits,
  output        io_stream_in_176_ready,
  input         io_stream_in_176_valid,
  input  [31:0] io_stream_in_176_bits,
  output        io_stream_in_177_ready,
  input         io_stream_in_177_valid,
  input  [31:0] io_stream_in_177_bits,
  output        io_stream_in_178_ready,
  input         io_stream_in_178_valid,
  input  [31:0] io_stream_in_178_bits,
  output        io_stream_in_179_ready,
  input         io_stream_in_179_valid,
  input  [31:0] io_stream_in_179_bits,
  output        io_stream_in_180_ready,
  input         io_stream_in_180_valid,
  input  [31:0] io_stream_in_180_bits,
  output        io_stream_in_181_ready,
  input         io_stream_in_181_valid,
  input  [31:0] io_stream_in_181_bits,
  output        io_stream_in_182_ready,
  input         io_stream_in_182_valid,
  input  [31:0] io_stream_in_182_bits,
  output        io_stream_in_183_ready,
  input         io_stream_in_183_valid,
  input  [31:0] io_stream_in_183_bits,
  output        io_stream_in_184_ready,
  input         io_stream_in_184_valid,
  input  [31:0] io_stream_in_184_bits,
  output        io_stream_in_185_ready,
  input         io_stream_in_185_valid,
  input  [31:0] io_stream_in_185_bits,
  output        io_stream_in_186_ready,
  input         io_stream_in_186_valid,
  input  [31:0] io_stream_in_186_bits,
  output        io_stream_in_187_ready,
  input         io_stream_in_187_valid,
  input  [31:0] io_stream_in_187_bits,
  output        io_stream_in_188_ready,
  input         io_stream_in_188_valid,
  input  [31:0] io_stream_in_188_bits,
  output        io_stream_in_189_ready,
  input         io_stream_in_189_valid,
  input  [31:0] io_stream_in_189_bits,
  output        io_stream_in_190_ready,
  input         io_stream_in_190_valid,
  input  [31:0] io_stream_in_190_bits,
  output        io_stream_in_191_ready,
  input         io_stream_in_191_valid,
  input  [31:0] io_stream_in_191_bits,
  output        io_stream_in_192_ready,
  input         io_stream_in_192_valid,
  input  [31:0] io_stream_in_192_bits,
  output        io_stream_in_193_ready,
  input         io_stream_in_193_valid,
  input  [31:0] io_stream_in_193_bits,
  output        io_stream_in_194_ready,
  input         io_stream_in_194_valid,
  input  [31:0] io_stream_in_194_bits,
  output        io_stream_in_195_ready,
  input         io_stream_in_195_valid,
  input  [31:0] io_stream_in_195_bits,
  output        io_stream_in_196_ready,
  input         io_stream_in_196_valid,
  input  [31:0] io_stream_in_196_bits,
  output        io_stream_in_197_ready,
  input         io_stream_in_197_valid,
  input  [31:0] io_stream_in_197_bits,
  output        io_stream_in_198_ready,
  input         io_stream_in_198_valid,
  input  [31:0] io_stream_in_198_bits,
  output        io_stream_in_199_ready,
  input         io_stream_in_199_valid,
  input  [31:0] io_stream_in_199_bits,
  output        io_stream_in_200_ready,
  input         io_stream_in_200_valid,
  input  [31:0] io_stream_in_200_bits,
  output        io_stream_in_201_ready,
  input         io_stream_in_201_valid,
  input  [31:0] io_stream_in_201_bits,
  output        io_stream_in_202_ready,
  input         io_stream_in_202_valid,
  input  [31:0] io_stream_in_202_bits,
  output        io_stream_in_203_ready,
  input         io_stream_in_203_valid,
  input  [31:0] io_stream_in_203_bits,
  output        io_stream_in_204_ready,
  input         io_stream_in_204_valid,
  input  [31:0] io_stream_in_204_bits,
  output        io_stream_in_205_ready,
  input         io_stream_in_205_valid,
  input  [31:0] io_stream_in_205_bits,
  output        io_stream_in_206_ready,
  input         io_stream_in_206_valid,
  input  [31:0] io_stream_in_206_bits,
  output        io_stream_in_207_ready,
  input         io_stream_in_207_valid,
  input  [31:0] io_stream_in_207_bits,
  output        io_stream_in_208_ready,
  input         io_stream_in_208_valid,
  input  [31:0] io_stream_in_208_bits,
  output        io_stream_in_209_ready,
  input         io_stream_in_209_valid,
  input  [31:0] io_stream_in_209_bits,
  output        io_stream_in_210_ready,
  input         io_stream_in_210_valid,
  input  [31:0] io_stream_in_210_bits,
  output        io_stream_in_211_ready,
  input         io_stream_in_211_valid,
  input  [31:0] io_stream_in_211_bits,
  output        io_stream_in_212_ready,
  input         io_stream_in_212_valid,
  input  [31:0] io_stream_in_212_bits,
  output        io_stream_in_213_ready,
  input         io_stream_in_213_valid,
  input  [31:0] io_stream_in_213_bits,
  output        io_stream_in_214_ready,
  input         io_stream_in_214_valid,
  input  [31:0] io_stream_in_214_bits,
  output        io_stream_in_215_ready,
  input         io_stream_in_215_valid,
  input  [31:0] io_stream_in_215_bits,
  output        io_stream_in_216_ready,
  input         io_stream_in_216_valid,
  input  [31:0] io_stream_in_216_bits,
  output        io_stream_in_217_ready,
  input         io_stream_in_217_valid,
  input  [31:0] io_stream_in_217_bits,
  output        io_stream_in_218_ready,
  input         io_stream_in_218_valid,
  input  [31:0] io_stream_in_218_bits,
  output        io_stream_in_219_ready,
  input         io_stream_in_219_valid,
  input  [31:0] io_stream_in_219_bits,
  output        io_stream_in_220_ready,
  input         io_stream_in_220_valid,
  input  [31:0] io_stream_in_220_bits,
  output        io_stream_in_221_ready,
  input         io_stream_in_221_valid,
  input  [31:0] io_stream_in_221_bits,
  output        io_stream_in_222_ready,
  input         io_stream_in_222_valid,
  input  [31:0] io_stream_in_222_bits,
  output        io_stream_in_223_ready,
  input         io_stream_in_223_valid,
  input  [31:0] io_stream_in_223_bits,
  output        io_stream_in_224_ready,
  input         io_stream_in_224_valid,
  input  [31:0] io_stream_in_224_bits,
  output        io_stream_in_225_ready,
  input         io_stream_in_225_valid,
  input  [31:0] io_stream_in_225_bits,
  output        io_stream_in_226_ready,
  input         io_stream_in_226_valid,
  input  [31:0] io_stream_in_226_bits,
  output        io_stream_in_227_ready,
  input         io_stream_in_227_valid,
  input  [31:0] io_stream_in_227_bits,
  output        io_stream_in_228_ready,
  input         io_stream_in_228_valid,
  input  [31:0] io_stream_in_228_bits,
  output        io_stream_in_229_ready,
  input         io_stream_in_229_valid,
  input  [31:0] io_stream_in_229_bits,
  output        io_stream_in_230_ready,
  input         io_stream_in_230_valid,
  input  [31:0] io_stream_in_230_bits,
  output        io_stream_in_231_ready,
  input         io_stream_in_231_valid,
  input  [31:0] io_stream_in_231_bits,
  output        io_stream_in_232_ready,
  input         io_stream_in_232_valid,
  input  [31:0] io_stream_in_232_bits,
  output        io_stream_in_233_ready,
  input         io_stream_in_233_valid,
  input  [31:0] io_stream_in_233_bits,
  output        io_stream_in_234_ready,
  input         io_stream_in_234_valid,
  input  [31:0] io_stream_in_234_bits,
  output        io_stream_in_235_ready,
  input         io_stream_in_235_valid,
  input  [31:0] io_stream_in_235_bits,
  output        io_stream_in_236_ready,
  input         io_stream_in_236_valid,
  input  [31:0] io_stream_in_236_bits,
  output        io_stream_in_237_ready,
  input         io_stream_in_237_valid,
  input  [31:0] io_stream_in_237_bits,
  output        io_stream_in_238_ready,
  input         io_stream_in_238_valid,
  input  [31:0] io_stream_in_238_bits,
  output        io_stream_in_239_ready,
  input         io_stream_in_239_valid,
  input  [31:0] io_stream_in_239_bits,
  output        io_stream_in_240_ready,
  input         io_stream_in_240_valid,
  input  [31:0] io_stream_in_240_bits,
  output        io_stream_in_241_ready,
  input         io_stream_in_241_valid,
  input  [31:0] io_stream_in_241_bits,
  output        io_stream_in_242_ready,
  input         io_stream_in_242_valid,
  input  [31:0] io_stream_in_242_bits,
  output        io_stream_in_243_ready,
  input         io_stream_in_243_valid,
  input  [31:0] io_stream_in_243_bits,
  output        io_stream_in_244_ready,
  input         io_stream_in_244_valid,
  input  [31:0] io_stream_in_244_bits,
  output        io_stream_in_245_ready,
  input         io_stream_in_245_valid,
  input  [31:0] io_stream_in_245_bits,
  output        io_stream_in_246_ready,
  input         io_stream_in_246_valid,
  input  [31:0] io_stream_in_246_bits,
  output        io_stream_in_247_ready,
  input         io_stream_in_247_valid,
  input  [31:0] io_stream_in_247_bits,
  output        io_stream_in_248_ready,
  input         io_stream_in_248_valid,
  input  [31:0] io_stream_in_248_bits,
  output        io_stream_in_249_ready,
  input         io_stream_in_249_valid,
  input  [31:0] io_stream_in_249_bits,
  output        io_stream_in_250_ready,
  input         io_stream_in_250_valid,
  input  [31:0] io_stream_in_250_bits,
  output        io_stream_in_251_ready,
  input         io_stream_in_251_valid,
  input  [31:0] io_stream_in_251_bits,
  output        io_stream_in_252_ready,
  input         io_stream_in_252_valid,
  input  [31:0] io_stream_in_252_bits,
  output        io_stream_in_253_ready,
  input         io_stream_in_253_valid,
  input  [31:0] io_stream_in_253_bits,
  output        io_stream_in_254_ready,
  input         io_stream_in_254_valid,
  input  [31:0] io_stream_in_254_bits,
  output        io_stream_in_255_ready,
  input         io_stream_in_255_valid,
  input  [31:0] io_stream_in_255_bits,
  input         io_stream_out_ready,
  output        io_stream_out_valid,
  output [31:0] io_stream_out_bits
);
  wire  last_merger_clock; // @[Stab.scala 175:24]
  wire  last_merger_reset; // @[Stab.scala 175:24]
  wire  last_merger_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_clock; // @[Decoupled.scala 361:21]
  wire  last_q_reset; // @[Decoupled.scala 361:21]
  wire  last_q_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_1_clock; // @[Stab.scala 175:24]
  wire  last_merger_1_reset; // @[Stab.scala 175:24]
  wire  last_merger_1_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_1_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_1_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_1_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_1_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_1_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_1_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_1_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_1_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_1_clock; // @[Decoupled.scala 361:21]
  wire  last_q_1_reset; // @[Decoupled.scala 361:21]
  wire  last_q_1_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_1_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_1_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_1_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_1_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_1_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_2_clock; // @[Stab.scala 175:24]
  wire  last_merger_2_reset; // @[Stab.scala 175:24]
  wire  last_merger_2_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_2_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_2_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_2_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_2_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_2_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_2_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_2_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_2_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_2_clock; // @[Decoupled.scala 361:21]
  wire  last_q_2_reset; // @[Decoupled.scala 361:21]
  wire  last_q_2_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_2_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_2_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_2_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_2_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_2_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_3_clock; // @[Stab.scala 175:24]
  wire  last_merger_3_reset; // @[Stab.scala 175:24]
  wire  last_merger_3_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_3_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_3_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_3_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_3_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_3_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_3_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_3_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_3_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_3_clock; // @[Decoupled.scala 361:21]
  wire  last_q_3_reset; // @[Decoupled.scala 361:21]
  wire  last_q_3_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_3_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_3_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_3_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_3_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_3_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_4_clock; // @[Stab.scala 175:24]
  wire  last_merger_4_reset; // @[Stab.scala 175:24]
  wire  last_merger_4_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_4_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_4_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_4_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_4_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_4_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_4_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_4_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_4_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_4_clock; // @[Decoupled.scala 361:21]
  wire  last_q_4_reset; // @[Decoupled.scala 361:21]
  wire  last_q_4_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_4_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_4_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_4_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_4_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_4_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_5_clock; // @[Stab.scala 175:24]
  wire  last_merger_5_reset; // @[Stab.scala 175:24]
  wire  last_merger_5_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_5_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_5_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_5_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_5_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_5_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_5_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_5_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_5_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_5_clock; // @[Decoupled.scala 361:21]
  wire  last_q_5_reset; // @[Decoupled.scala 361:21]
  wire  last_q_5_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_5_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_5_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_5_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_5_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_5_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_6_clock; // @[Stab.scala 175:24]
  wire  last_merger_6_reset; // @[Stab.scala 175:24]
  wire  last_merger_6_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_6_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_6_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_6_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_6_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_6_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_6_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_6_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_6_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_6_clock; // @[Decoupled.scala 361:21]
  wire  last_q_6_reset; // @[Decoupled.scala 361:21]
  wire  last_q_6_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_6_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_6_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_6_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_6_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_6_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_7_clock; // @[Stab.scala 175:24]
  wire  last_merger_7_reset; // @[Stab.scala 175:24]
  wire  last_merger_7_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_7_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_7_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_7_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_7_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_7_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_7_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_7_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_7_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_7_clock; // @[Decoupled.scala 361:21]
  wire  last_q_7_reset; // @[Decoupled.scala 361:21]
  wire  last_q_7_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_7_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_7_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_7_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_7_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_7_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_8_clock; // @[Stab.scala 175:24]
  wire  last_merger_8_reset; // @[Stab.scala 175:24]
  wire  last_merger_8_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_8_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_8_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_8_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_8_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_8_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_8_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_8_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_8_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_8_clock; // @[Decoupled.scala 361:21]
  wire  last_q_8_reset; // @[Decoupled.scala 361:21]
  wire  last_q_8_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_8_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_8_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_8_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_8_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_8_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_9_clock; // @[Stab.scala 175:24]
  wire  last_merger_9_reset; // @[Stab.scala 175:24]
  wire  last_merger_9_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_9_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_9_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_9_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_9_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_9_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_9_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_9_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_9_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_9_clock; // @[Decoupled.scala 361:21]
  wire  last_q_9_reset; // @[Decoupled.scala 361:21]
  wire  last_q_9_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_9_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_9_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_9_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_9_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_9_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_10_clock; // @[Stab.scala 175:24]
  wire  last_merger_10_reset; // @[Stab.scala 175:24]
  wire  last_merger_10_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_10_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_10_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_10_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_10_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_10_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_10_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_10_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_10_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_10_clock; // @[Decoupled.scala 361:21]
  wire  last_q_10_reset; // @[Decoupled.scala 361:21]
  wire  last_q_10_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_10_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_10_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_10_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_10_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_10_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_11_clock; // @[Stab.scala 175:24]
  wire  last_merger_11_reset; // @[Stab.scala 175:24]
  wire  last_merger_11_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_11_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_11_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_11_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_11_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_11_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_11_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_11_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_11_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_11_clock; // @[Decoupled.scala 361:21]
  wire  last_q_11_reset; // @[Decoupled.scala 361:21]
  wire  last_q_11_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_11_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_11_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_11_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_11_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_11_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_12_clock; // @[Stab.scala 175:24]
  wire  last_merger_12_reset; // @[Stab.scala 175:24]
  wire  last_merger_12_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_12_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_12_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_12_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_12_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_12_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_12_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_12_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_12_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_12_clock; // @[Decoupled.scala 361:21]
  wire  last_q_12_reset; // @[Decoupled.scala 361:21]
  wire  last_q_12_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_12_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_12_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_12_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_12_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_12_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_13_clock; // @[Stab.scala 175:24]
  wire  last_merger_13_reset; // @[Stab.scala 175:24]
  wire  last_merger_13_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_13_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_13_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_13_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_13_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_13_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_13_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_13_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_13_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_13_clock; // @[Decoupled.scala 361:21]
  wire  last_q_13_reset; // @[Decoupled.scala 361:21]
  wire  last_q_13_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_13_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_13_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_13_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_13_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_13_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_14_clock; // @[Stab.scala 175:24]
  wire  last_merger_14_reset; // @[Stab.scala 175:24]
  wire  last_merger_14_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_14_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_14_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_14_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_14_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_14_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_14_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_14_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_14_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_14_clock; // @[Decoupled.scala 361:21]
  wire  last_q_14_reset; // @[Decoupled.scala 361:21]
  wire  last_q_14_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_14_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_14_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_14_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_14_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_14_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_15_clock; // @[Stab.scala 175:24]
  wire  last_merger_15_reset; // @[Stab.scala 175:24]
  wire  last_merger_15_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_15_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_15_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_15_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_15_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_15_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_15_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_15_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_15_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_15_clock; // @[Decoupled.scala 361:21]
  wire  last_q_15_reset; // @[Decoupled.scala 361:21]
  wire  last_q_15_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_15_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_15_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_15_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_15_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_15_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_16_clock; // @[Stab.scala 175:24]
  wire  last_merger_16_reset; // @[Stab.scala 175:24]
  wire  last_merger_16_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_16_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_16_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_16_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_16_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_16_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_16_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_16_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_16_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_16_clock; // @[Decoupled.scala 361:21]
  wire  last_q_16_reset; // @[Decoupled.scala 361:21]
  wire  last_q_16_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_16_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_16_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_16_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_16_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_16_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_17_clock; // @[Stab.scala 175:24]
  wire  last_merger_17_reset; // @[Stab.scala 175:24]
  wire  last_merger_17_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_17_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_17_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_17_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_17_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_17_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_17_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_17_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_17_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_17_clock; // @[Decoupled.scala 361:21]
  wire  last_q_17_reset; // @[Decoupled.scala 361:21]
  wire  last_q_17_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_17_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_17_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_17_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_17_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_17_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_18_clock; // @[Stab.scala 175:24]
  wire  last_merger_18_reset; // @[Stab.scala 175:24]
  wire  last_merger_18_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_18_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_18_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_18_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_18_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_18_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_18_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_18_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_18_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_18_clock; // @[Decoupled.scala 361:21]
  wire  last_q_18_reset; // @[Decoupled.scala 361:21]
  wire  last_q_18_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_18_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_18_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_18_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_18_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_18_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_19_clock; // @[Stab.scala 175:24]
  wire  last_merger_19_reset; // @[Stab.scala 175:24]
  wire  last_merger_19_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_19_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_19_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_19_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_19_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_19_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_19_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_19_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_19_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_19_clock; // @[Decoupled.scala 361:21]
  wire  last_q_19_reset; // @[Decoupled.scala 361:21]
  wire  last_q_19_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_19_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_19_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_19_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_19_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_19_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_20_clock; // @[Stab.scala 175:24]
  wire  last_merger_20_reset; // @[Stab.scala 175:24]
  wire  last_merger_20_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_20_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_20_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_20_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_20_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_20_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_20_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_20_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_20_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_20_clock; // @[Decoupled.scala 361:21]
  wire  last_q_20_reset; // @[Decoupled.scala 361:21]
  wire  last_q_20_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_20_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_20_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_20_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_20_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_20_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_21_clock; // @[Stab.scala 175:24]
  wire  last_merger_21_reset; // @[Stab.scala 175:24]
  wire  last_merger_21_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_21_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_21_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_21_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_21_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_21_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_21_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_21_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_21_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_21_clock; // @[Decoupled.scala 361:21]
  wire  last_q_21_reset; // @[Decoupled.scala 361:21]
  wire  last_q_21_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_21_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_21_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_21_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_21_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_21_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_22_clock; // @[Stab.scala 175:24]
  wire  last_merger_22_reset; // @[Stab.scala 175:24]
  wire  last_merger_22_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_22_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_22_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_22_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_22_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_22_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_22_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_22_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_22_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_22_clock; // @[Decoupled.scala 361:21]
  wire  last_q_22_reset; // @[Decoupled.scala 361:21]
  wire  last_q_22_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_22_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_22_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_22_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_22_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_22_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_23_clock; // @[Stab.scala 175:24]
  wire  last_merger_23_reset; // @[Stab.scala 175:24]
  wire  last_merger_23_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_23_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_23_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_23_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_23_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_23_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_23_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_23_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_23_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_23_clock; // @[Decoupled.scala 361:21]
  wire  last_q_23_reset; // @[Decoupled.scala 361:21]
  wire  last_q_23_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_23_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_23_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_23_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_23_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_23_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_24_clock; // @[Stab.scala 175:24]
  wire  last_merger_24_reset; // @[Stab.scala 175:24]
  wire  last_merger_24_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_24_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_24_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_24_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_24_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_24_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_24_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_24_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_24_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_24_clock; // @[Decoupled.scala 361:21]
  wire  last_q_24_reset; // @[Decoupled.scala 361:21]
  wire  last_q_24_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_24_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_24_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_24_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_24_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_24_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_25_clock; // @[Stab.scala 175:24]
  wire  last_merger_25_reset; // @[Stab.scala 175:24]
  wire  last_merger_25_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_25_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_25_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_25_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_25_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_25_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_25_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_25_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_25_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_25_clock; // @[Decoupled.scala 361:21]
  wire  last_q_25_reset; // @[Decoupled.scala 361:21]
  wire  last_q_25_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_25_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_25_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_25_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_25_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_25_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_26_clock; // @[Stab.scala 175:24]
  wire  last_merger_26_reset; // @[Stab.scala 175:24]
  wire  last_merger_26_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_26_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_26_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_26_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_26_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_26_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_26_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_26_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_26_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_26_clock; // @[Decoupled.scala 361:21]
  wire  last_q_26_reset; // @[Decoupled.scala 361:21]
  wire  last_q_26_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_26_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_26_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_26_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_26_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_26_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_27_clock; // @[Stab.scala 175:24]
  wire  last_merger_27_reset; // @[Stab.scala 175:24]
  wire  last_merger_27_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_27_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_27_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_27_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_27_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_27_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_27_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_27_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_27_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_27_clock; // @[Decoupled.scala 361:21]
  wire  last_q_27_reset; // @[Decoupled.scala 361:21]
  wire  last_q_27_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_27_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_27_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_27_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_27_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_27_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_28_clock; // @[Stab.scala 175:24]
  wire  last_merger_28_reset; // @[Stab.scala 175:24]
  wire  last_merger_28_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_28_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_28_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_28_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_28_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_28_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_28_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_28_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_28_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_28_clock; // @[Decoupled.scala 361:21]
  wire  last_q_28_reset; // @[Decoupled.scala 361:21]
  wire  last_q_28_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_28_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_28_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_28_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_28_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_28_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_29_clock; // @[Stab.scala 175:24]
  wire  last_merger_29_reset; // @[Stab.scala 175:24]
  wire  last_merger_29_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_29_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_29_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_29_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_29_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_29_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_29_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_29_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_29_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_29_clock; // @[Decoupled.scala 361:21]
  wire  last_q_29_reset; // @[Decoupled.scala 361:21]
  wire  last_q_29_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_29_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_29_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_29_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_29_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_29_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_30_clock; // @[Stab.scala 175:24]
  wire  last_merger_30_reset; // @[Stab.scala 175:24]
  wire  last_merger_30_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_30_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_30_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_30_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_30_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_30_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_30_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_30_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_30_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_30_clock; // @[Decoupled.scala 361:21]
  wire  last_q_30_reset; // @[Decoupled.scala 361:21]
  wire  last_q_30_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_30_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_30_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_30_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_30_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_30_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_31_clock; // @[Stab.scala 175:24]
  wire  last_merger_31_reset; // @[Stab.scala 175:24]
  wire  last_merger_31_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_31_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_31_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_31_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_31_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_31_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_31_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_31_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_31_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_31_clock; // @[Decoupled.scala 361:21]
  wire  last_q_31_reset; // @[Decoupled.scala 361:21]
  wire  last_q_31_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_31_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_31_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_31_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_31_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_31_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_32_clock; // @[Stab.scala 175:24]
  wire  last_merger_32_reset; // @[Stab.scala 175:24]
  wire  last_merger_32_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_32_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_32_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_32_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_32_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_32_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_32_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_32_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_32_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_32_clock; // @[Decoupled.scala 361:21]
  wire  last_q_32_reset; // @[Decoupled.scala 361:21]
  wire  last_q_32_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_32_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_32_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_32_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_32_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_32_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_33_clock; // @[Stab.scala 175:24]
  wire  last_merger_33_reset; // @[Stab.scala 175:24]
  wire  last_merger_33_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_33_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_33_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_33_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_33_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_33_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_33_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_33_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_33_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_33_clock; // @[Decoupled.scala 361:21]
  wire  last_q_33_reset; // @[Decoupled.scala 361:21]
  wire  last_q_33_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_33_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_33_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_33_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_33_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_33_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_34_clock; // @[Stab.scala 175:24]
  wire  last_merger_34_reset; // @[Stab.scala 175:24]
  wire  last_merger_34_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_34_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_34_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_34_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_34_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_34_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_34_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_34_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_34_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_34_clock; // @[Decoupled.scala 361:21]
  wire  last_q_34_reset; // @[Decoupled.scala 361:21]
  wire  last_q_34_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_34_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_34_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_34_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_34_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_34_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_35_clock; // @[Stab.scala 175:24]
  wire  last_merger_35_reset; // @[Stab.scala 175:24]
  wire  last_merger_35_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_35_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_35_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_35_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_35_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_35_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_35_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_35_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_35_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_35_clock; // @[Decoupled.scala 361:21]
  wire  last_q_35_reset; // @[Decoupled.scala 361:21]
  wire  last_q_35_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_35_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_35_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_35_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_35_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_35_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_36_clock; // @[Stab.scala 175:24]
  wire  last_merger_36_reset; // @[Stab.scala 175:24]
  wire  last_merger_36_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_36_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_36_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_36_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_36_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_36_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_36_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_36_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_36_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_36_clock; // @[Decoupled.scala 361:21]
  wire  last_q_36_reset; // @[Decoupled.scala 361:21]
  wire  last_q_36_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_36_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_36_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_36_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_36_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_36_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_37_clock; // @[Stab.scala 175:24]
  wire  last_merger_37_reset; // @[Stab.scala 175:24]
  wire  last_merger_37_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_37_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_37_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_37_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_37_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_37_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_37_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_37_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_37_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_37_clock; // @[Decoupled.scala 361:21]
  wire  last_q_37_reset; // @[Decoupled.scala 361:21]
  wire  last_q_37_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_37_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_37_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_37_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_37_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_37_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_38_clock; // @[Stab.scala 175:24]
  wire  last_merger_38_reset; // @[Stab.scala 175:24]
  wire  last_merger_38_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_38_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_38_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_38_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_38_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_38_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_38_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_38_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_38_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_38_clock; // @[Decoupled.scala 361:21]
  wire  last_q_38_reset; // @[Decoupled.scala 361:21]
  wire  last_q_38_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_38_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_38_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_38_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_38_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_38_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_39_clock; // @[Stab.scala 175:24]
  wire  last_merger_39_reset; // @[Stab.scala 175:24]
  wire  last_merger_39_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_39_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_39_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_39_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_39_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_39_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_39_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_39_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_39_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_39_clock; // @[Decoupled.scala 361:21]
  wire  last_q_39_reset; // @[Decoupled.scala 361:21]
  wire  last_q_39_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_39_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_39_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_39_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_39_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_39_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_40_clock; // @[Stab.scala 175:24]
  wire  last_merger_40_reset; // @[Stab.scala 175:24]
  wire  last_merger_40_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_40_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_40_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_40_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_40_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_40_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_40_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_40_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_40_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_40_clock; // @[Decoupled.scala 361:21]
  wire  last_q_40_reset; // @[Decoupled.scala 361:21]
  wire  last_q_40_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_40_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_40_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_40_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_40_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_40_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_41_clock; // @[Stab.scala 175:24]
  wire  last_merger_41_reset; // @[Stab.scala 175:24]
  wire  last_merger_41_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_41_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_41_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_41_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_41_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_41_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_41_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_41_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_41_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_41_clock; // @[Decoupled.scala 361:21]
  wire  last_q_41_reset; // @[Decoupled.scala 361:21]
  wire  last_q_41_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_41_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_41_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_41_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_41_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_41_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_42_clock; // @[Stab.scala 175:24]
  wire  last_merger_42_reset; // @[Stab.scala 175:24]
  wire  last_merger_42_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_42_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_42_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_42_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_42_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_42_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_42_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_42_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_42_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_42_clock; // @[Decoupled.scala 361:21]
  wire  last_q_42_reset; // @[Decoupled.scala 361:21]
  wire  last_q_42_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_42_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_42_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_42_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_42_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_42_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_43_clock; // @[Stab.scala 175:24]
  wire  last_merger_43_reset; // @[Stab.scala 175:24]
  wire  last_merger_43_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_43_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_43_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_43_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_43_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_43_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_43_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_43_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_43_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_43_clock; // @[Decoupled.scala 361:21]
  wire  last_q_43_reset; // @[Decoupled.scala 361:21]
  wire  last_q_43_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_43_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_43_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_43_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_43_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_43_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_44_clock; // @[Stab.scala 175:24]
  wire  last_merger_44_reset; // @[Stab.scala 175:24]
  wire  last_merger_44_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_44_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_44_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_44_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_44_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_44_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_44_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_44_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_44_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_44_clock; // @[Decoupled.scala 361:21]
  wire  last_q_44_reset; // @[Decoupled.scala 361:21]
  wire  last_q_44_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_44_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_44_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_44_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_44_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_44_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_45_clock; // @[Stab.scala 175:24]
  wire  last_merger_45_reset; // @[Stab.scala 175:24]
  wire  last_merger_45_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_45_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_45_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_45_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_45_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_45_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_45_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_45_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_45_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_45_clock; // @[Decoupled.scala 361:21]
  wire  last_q_45_reset; // @[Decoupled.scala 361:21]
  wire  last_q_45_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_45_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_45_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_45_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_45_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_45_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_46_clock; // @[Stab.scala 175:24]
  wire  last_merger_46_reset; // @[Stab.scala 175:24]
  wire  last_merger_46_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_46_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_46_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_46_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_46_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_46_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_46_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_46_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_46_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_46_clock; // @[Decoupled.scala 361:21]
  wire  last_q_46_reset; // @[Decoupled.scala 361:21]
  wire  last_q_46_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_46_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_46_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_46_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_46_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_46_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_47_clock; // @[Stab.scala 175:24]
  wire  last_merger_47_reset; // @[Stab.scala 175:24]
  wire  last_merger_47_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_47_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_47_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_47_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_47_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_47_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_47_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_47_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_47_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_47_clock; // @[Decoupled.scala 361:21]
  wire  last_q_47_reset; // @[Decoupled.scala 361:21]
  wire  last_q_47_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_47_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_47_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_47_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_47_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_47_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_48_clock; // @[Stab.scala 175:24]
  wire  last_merger_48_reset; // @[Stab.scala 175:24]
  wire  last_merger_48_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_48_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_48_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_48_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_48_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_48_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_48_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_48_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_48_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_48_clock; // @[Decoupled.scala 361:21]
  wire  last_q_48_reset; // @[Decoupled.scala 361:21]
  wire  last_q_48_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_48_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_48_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_48_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_48_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_48_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_49_clock; // @[Stab.scala 175:24]
  wire  last_merger_49_reset; // @[Stab.scala 175:24]
  wire  last_merger_49_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_49_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_49_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_49_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_49_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_49_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_49_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_49_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_49_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_49_clock; // @[Decoupled.scala 361:21]
  wire  last_q_49_reset; // @[Decoupled.scala 361:21]
  wire  last_q_49_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_49_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_49_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_49_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_49_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_49_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_50_clock; // @[Stab.scala 175:24]
  wire  last_merger_50_reset; // @[Stab.scala 175:24]
  wire  last_merger_50_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_50_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_50_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_50_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_50_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_50_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_50_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_50_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_50_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_50_clock; // @[Decoupled.scala 361:21]
  wire  last_q_50_reset; // @[Decoupled.scala 361:21]
  wire  last_q_50_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_50_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_50_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_50_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_50_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_50_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_51_clock; // @[Stab.scala 175:24]
  wire  last_merger_51_reset; // @[Stab.scala 175:24]
  wire  last_merger_51_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_51_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_51_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_51_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_51_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_51_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_51_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_51_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_51_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_51_clock; // @[Decoupled.scala 361:21]
  wire  last_q_51_reset; // @[Decoupled.scala 361:21]
  wire  last_q_51_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_51_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_51_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_51_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_51_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_51_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_52_clock; // @[Stab.scala 175:24]
  wire  last_merger_52_reset; // @[Stab.scala 175:24]
  wire  last_merger_52_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_52_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_52_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_52_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_52_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_52_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_52_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_52_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_52_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_52_clock; // @[Decoupled.scala 361:21]
  wire  last_q_52_reset; // @[Decoupled.scala 361:21]
  wire  last_q_52_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_52_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_52_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_52_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_52_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_52_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_53_clock; // @[Stab.scala 175:24]
  wire  last_merger_53_reset; // @[Stab.scala 175:24]
  wire  last_merger_53_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_53_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_53_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_53_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_53_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_53_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_53_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_53_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_53_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_53_clock; // @[Decoupled.scala 361:21]
  wire  last_q_53_reset; // @[Decoupled.scala 361:21]
  wire  last_q_53_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_53_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_53_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_53_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_53_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_53_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_54_clock; // @[Stab.scala 175:24]
  wire  last_merger_54_reset; // @[Stab.scala 175:24]
  wire  last_merger_54_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_54_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_54_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_54_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_54_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_54_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_54_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_54_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_54_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_54_clock; // @[Decoupled.scala 361:21]
  wire  last_q_54_reset; // @[Decoupled.scala 361:21]
  wire  last_q_54_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_54_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_54_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_54_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_54_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_54_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_55_clock; // @[Stab.scala 175:24]
  wire  last_merger_55_reset; // @[Stab.scala 175:24]
  wire  last_merger_55_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_55_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_55_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_55_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_55_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_55_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_55_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_55_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_55_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_55_clock; // @[Decoupled.scala 361:21]
  wire  last_q_55_reset; // @[Decoupled.scala 361:21]
  wire  last_q_55_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_55_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_55_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_55_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_55_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_55_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_56_clock; // @[Stab.scala 175:24]
  wire  last_merger_56_reset; // @[Stab.scala 175:24]
  wire  last_merger_56_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_56_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_56_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_56_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_56_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_56_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_56_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_56_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_56_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_56_clock; // @[Decoupled.scala 361:21]
  wire  last_q_56_reset; // @[Decoupled.scala 361:21]
  wire  last_q_56_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_56_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_56_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_56_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_56_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_56_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_57_clock; // @[Stab.scala 175:24]
  wire  last_merger_57_reset; // @[Stab.scala 175:24]
  wire  last_merger_57_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_57_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_57_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_57_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_57_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_57_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_57_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_57_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_57_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_57_clock; // @[Decoupled.scala 361:21]
  wire  last_q_57_reset; // @[Decoupled.scala 361:21]
  wire  last_q_57_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_57_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_57_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_57_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_57_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_57_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_58_clock; // @[Stab.scala 175:24]
  wire  last_merger_58_reset; // @[Stab.scala 175:24]
  wire  last_merger_58_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_58_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_58_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_58_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_58_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_58_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_58_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_58_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_58_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_58_clock; // @[Decoupled.scala 361:21]
  wire  last_q_58_reset; // @[Decoupled.scala 361:21]
  wire  last_q_58_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_58_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_58_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_58_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_58_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_58_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_59_clock; // @[Stab.scala 175:24]
  wire  last_merger_59_reset; // @[Stab.scala 175:24]
  wire  last_merger_59_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_59_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_59_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_59_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_59_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_59_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_59_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_59_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_59_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_59_clock; // @[Decoupled.scala 361:21]
  wire  last_q_59_reset; // @[Decoupled.scala 361:21]
  wire  last_q_59_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_59_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_59_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_59_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_59_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_59_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_60_clock; // @[Stab.scala 175:24]
  wire  last_merger_60_reset; // @[Stab.scala 175:24]
  wire  last_merger_60_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_60_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_60_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_60_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_60_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_60_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_60_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_60_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_60_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_60_clock; // @[Decoupled.scala 361:21]
  wire  last_q_60_reset; // @[Decoupled.scala 361:21]
  wire  last_q_60_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_60_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_60_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_60_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_60_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_60_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_61_clock; // @[Stab.scala 175:24]
  wire  last_merger_61_reset; // @[Stab.scala 175:24]
  wire  last_merger_61_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_61_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_61_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_61_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_61_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_61_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_61_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_61_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_61_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_61_clock; // @[Decoupled.scala 361:21]
  wire  last_q_61_reset; // @[Decoupled.scala 361:21]
  wire  last_q_61_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_61_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_61_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_61_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_61_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_61_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_62_clock; // @[Stab.scala 175:24]
  wire  last_merger_62_reset; // @[Stab.scala 175:24]
  wire  last_merger_62_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_62_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_62_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_62_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_62_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_62_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_62_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_62_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_62_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_62_clock; // @[Decoupled.scala 361:21]
  wire  last_q_62_reset; // @[Decoupled.scala 361:21]
  wire  last_q_62_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_62_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_62_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_62_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_62_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_62_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_63_clock; // @[Stab.scala 175:24]
  wire  last_merger_63_reset; // @[Stab.scala 175:24]
  wire  last_merger_63_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_63_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_63_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_63_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_63_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_63_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_63_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_63_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_63_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_63_clock; // @[Decoupled.scala 361:21]
  wire  last_q_63_reset; // @[Decoupled.scala 361:21]
  wire  last_q_63_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_63_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_63_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_63_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_63_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_63_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_64_clock; // @[Stab.scala 175:24]
  wire  last_merger_64_reset; // @[Stab.scala 175:24]
  wire  last_merger_64_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_64_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_64_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_64_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_64_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_64_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_64_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_64_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_64_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_64_clock; // @[Decoupled.scala 361:21]
  wire  last_q_64_reset; // @[Decoupled.scala 361:21]
  wire  last_q_64_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_64_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_64_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_64_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_64_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_64_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_65_clock; // @[Stab.scala 175:24]
  wire  last_merger_65_reset; // @[Stab.scala 175:24]
  wire  last_merger_65_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_65_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_65_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_65_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_65_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_65_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_65_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_65_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_65_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_65_clock; // @[Decoupled.scala 361:21]
  wire  last_q_65_reset; // @[Decoupled.scala 361:21]
  wire  last_q_65_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_65_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_65_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_65_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_65_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_65_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_66_clock; // @[Stab.scala 175:24]
  wire  last_merger_66_reset; // @[Stab.scala 175:24]
  wire  last_merger_66_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_66_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_66_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_66_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_66_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_66_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_66_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_66_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_66_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_66_clock; // @[Decoupled.scala 361:21]
  wire  last_q_66_reset; // @[Decoupled.scala 361:21]
  wire  last_q_66_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_66_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_66_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_66_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_66_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_66_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_67_clock; // @[Stab.scala 175:24]
  wire  last_merger_67_reset; // @[Stab.scala 175:24]
  wire  last_merger_67_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_67_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_67_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_67_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_67_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_67_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_67_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_67_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_67_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_67_clock; // @[Decoupled.scala 361:21]
  wire  last_q_67_reset; // @[Decoupled.scala 361:21]
  wire  last_q_67_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_67_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_67_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_67_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_67_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_67_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_68_clock; // @[Stab.scala 175:24]
  wire  last_merger_68_reset; // @[Stab.scala 175:24]
  wire  last_merger_68_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_68_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_68_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_68_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_68_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_68_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_68_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_68_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_68_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_68_clock; // @[Decoupled.scala 361:21]
  wire  last_q_68_reset; // @[Decoupled.scala 361:21]
  wire  last_q_68_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_68_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_68_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_68_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_68_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_68_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_69_clock; // @[Stab.scala 175:24]
  wire  last_merger_69_reset; // @[Stab.scala 175:24]
  wire  last_merger_69_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_69_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_69_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_69_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_69_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_69_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_69_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_69_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_69_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_69_clock; // @[Decoupled.scala 361:21]
  wire  last_q_69_reset; // @[Decoupled.scala 361:21]
  wire  last_q_69_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_69_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_69_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_69_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_69_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_69_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_70_clock; // @[Stab.scala 175:24]
  wire  last_merger_70_reset; // @[Stab.scala 175:24]
  wire  last_merger_70_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_70_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_70_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_70_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_70_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_70_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_70_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_70_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_70_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_70_clock; // @[Decoupled.scala 361:21]
  wire  last_q_70_reset; // @[Decoupled.scala 361:21]
  wire  last_q_70_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_70_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_70_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_70_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_70_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_70_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_71_clock; // @[Stab.scala 175:24]
  wire  last_merger_71_reset; // @[Stab.scala 175:24]
  wire  last_merger_71_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_71_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_71_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_71_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_71_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_71_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_71_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_71_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_71_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_71_clock; // @[Decoupled.scala 361:21]
  wire  last_q_71_reset; // @[Decoupled.scala 361:21]
  wire  last_q_71_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_71_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_71_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_71_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_71_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_71_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_72_clock; // @[Stab.scala 175:24]
  wire  last_merger_72_reset; // @[Stab.scala 175:24]
  wire  last_merger_72_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_72_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_72_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_72_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_72_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_72_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_72_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_72_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_72_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_72_clock; // @[Decoupled.scala 361:21]
  wire  last_q_72_reset; // @[Decoupled.scala 361:21]
  wire  last_q_72_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_72_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_72_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_72_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_72_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_72_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_73_clock; // @[Stab.scala 175:24]
  wire  last_merger_73_reset; // @[Stab.scala 175:24]
  wire  last_merger_73_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_73_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_73_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_73_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_73_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_73_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_73_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_73_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_73_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_73_clock; // @[Decoupled.scala 361:21]
  wire  last_q_73_reset; // @[Decoupled.scala 361:21]
  wire  last_q_73_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_73_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_73_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_73_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_73_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_73_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_74_clock; // @[Stab.scala 175:24]
  wire  last_merger_74_reset; // @[Stab.scala 175:24]
  wire  last_merger_74_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_74_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_74_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_74_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_74_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_74_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_74_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_74_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_74_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_74_clock; // @[Decoupled.scala 361:21]
  wire  last_q_74_reset; // @[Decoupled.scala 361:21]
  wire  last_q_74_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_74_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_74_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_74_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_74_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_74_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_75_clock; // @[Stab.scala 175:24]
  wire  last_merger_75_reset; // @[Stab.scala 175:24]
  wire  last_merger_75_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_75_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_75_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_75_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_75_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_75_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_75_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_75_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_75_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_75_clock; // @[Decoupled.scala 361:21]
  wire  last_q_75_reset; // @[Decoupled.scala 361:21]
  wire  last_q_75_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_75_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_75_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_75_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_75_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_75_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_76_clock; // @[Stab.scala 175:24]
  wire  last_merger_76_reset; // @[Stab.scala 175:24]
  wire  last_merger_76_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_76_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_76_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_76_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_76_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_76_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_76_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_76_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_76_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_76_clock; // @[Decoupled.scala 361:21]
  wire  last_q_76_reset; // @[Decoupled.scala 361:21]
  wire  last_q_76_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_76_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_76_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_76_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_76_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_76_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_77_clock; // @[Stab.scala 175:24]
  wire  last_merger_77_reset; // @[Stab.scala 175:24]
  wire  last_merger_77_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_77_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_77_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_77_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_77_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_77_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_77_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_77_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_77_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_77_clock; // @[Decoupled.scala 361:21]
  wire  last_q_77_reset; // @[Decoupled.scala 361:21]
  wire  last_q_77_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_77_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_77_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_77_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_77_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_77_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_78_clock; // @[Stab.scala 175:24]
  wire  last_merger_78_reset; // @[Stab.scala 175:24]
  wire  last_merger_78_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_78_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_78_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_78_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_78_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_78_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_78_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_78_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_78_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_78_clock; // @[Decoupled.scala 361:21]
  wire  last_q_78_reset; // @[Decoupled.scala 361:21]
  wire  last_q_78_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_78_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_78_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_78_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_78_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_78_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_79_clock; // @[Stab.scala 175:24]
  wire  last_merger_79_reset; // @[Stab.scala 175:24]
  wire  last_merger_79_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_79_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_79_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_79_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_79_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_79_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_79_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_79_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_79_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_79_clock; // @[Decoupled.scala 361:21]
  wire  last_q_79_reset; // @[Decoupled.scala 361:21]
  wire  last_q_79_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_79_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_79_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_79_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_79_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_79_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_80_clock; // @[Stab.scala 175:24]
  wire  last_merger_80_reset; // @[Stab.scala 175:24]
  wire  last_merger_80_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_80_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_80_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_80_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_80_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_80_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_80_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_80_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_80_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_80_clock; // @[Decoupled.scala 361:21]
  wire  last_q_80_reset; // @[Decoupled.scala 361:21]
  wire  last_q_80_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_80_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_80_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_80_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_80_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_80_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_81_clock; // @[Stab.scala 175:24]
  wire  last_merger_81_reset; // @[Stab.scala 175:24]
  wire  last_merger_81_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_81_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_81_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_81_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_81_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_81_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_81_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_81_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_81_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_81_clock; // @[Decoupled.scala 361:21]
  wire  last_q_81_reset; // @[Decoupled.scala 361:21]
  wire  last_q_81_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_81_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_81_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_81_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_81_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_81_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_82_clock; // @[Stab.scala 175:24]
  wire  last_merger_82_reset; // @[Stab.scala 175:24]
  wire  last_merger_82_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_82_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_82_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_82_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_82_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_82_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_82_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_82_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_82_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_82_clock; // @[Decoupled.scala 361:21]
  wire  last_q_82_reset; // @[Decoupled.scala 361:21]
  wire  last_q_82_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_82_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_82_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_82_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_82_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_82_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_83_clock; // @[Stab.scala 175:24]
  wire  last_merger_83_reset; // @[Stab.scala 175:24]
  wire  last_merger_83_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_83_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_83_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_83_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_83_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_83_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_83_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_83_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_83_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_83_clock; // @[Decoupled.scala 361:21]
  wire  last_q_83_reset; // @[Decoupled.scala 361:21]
  wire  last_q_83_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_83_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_83_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_83_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_83_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_83_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_84_clock; // @[Stab.scala 175:24]
  wire  last_merger_84_reset; // @[Stab.scala 175:24]
  wire  last_merger_84_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_84_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_84_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_84_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_84_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_84_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_84_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_84_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_84_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_84_clock; // @[Decoupled.scala 361:21]
  wire  last_q_84_reset; // @[Decoupled.scala 361:21]
  wire  last_q_84_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_84_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_84_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_84_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_84_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_84_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_85_clock; // @[Stab.scala 175:24]
  wire  last_merger_85_reset; // @[Stab.scala 175:24]
  wire  last_merger_85_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_85_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_85_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_85_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_85_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_85_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_85_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_85_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_85_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_85_clock; // @[Decoupled.scala 361:21]
  wire  last_q_85_reset; // @[Decoupled.scala 361:21]
  wire  last_q_85_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_85_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_85_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_85_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_85_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_85_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_86_clock; // @[Stab.scala 175:24]
  wire  last_merger_86_reset; // @[Stab.scala 175:24]
  wire  last_merger_86_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_86_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_86_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_86_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_86_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_86_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_86_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_86_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_86_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_86_clock; // @[Decoupled.scala 361:21]
  wire  last_q_86_reset; // @[Decoupled.scala 361:21]
  wire  last_q_86_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_86_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_86_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_86_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_86_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_86_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_87_clock; // @[Stab.scala 175:24]
  wire  last_merger_87_reset; // @[Stab.scala 175:24]
  wire  last_merger_87_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_87_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_87_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_87_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_87_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_87_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_87_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_87_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_87_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_87_clock; // @[Decoupled.scala 361:21]
  wire  last_q_87_reset; // @[Decoupled.scala 361:21]
  wire  last_q_87_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_87_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_87_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_87_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_87_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_87_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_88_clock; // @[Stab.scala 175:24]
  wire  last_merger_88_reset; // @[Stab.scala 175:24]
  wire  last_merger_88_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_88_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_88_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_88_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_88_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_88_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_88_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_88_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_88_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_88_clock; // @[Decoupled.scala 361:21]
  wire  last_q_88_reset; // @[Decoupled.scala 361:21]
  wire  last_q_88_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_88_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_88_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_88_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_88_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_88_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_89_clock; // @[Stab.scala 175:24]
  wire  last_merger_89_reset; // @[Stab.scala 175:24]
  wire  last_merger_89_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_89_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_89_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_89_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_89_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_89_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_89_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_89_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_89_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_89_clock; // @[Decoupled.scala 361:21]
  wire  last_q_89_reset; // @[Decoupled.scala 361:21]
  wire  last_q_89_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_89_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_89_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_89_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_89_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_89_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_90_clock; // @[Stab.scala 175:24]
  wire  last_merger_90_reset; // @[Stab.scala 175:24]
  wire  last_merger_90_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_90_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_90_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_90_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_90_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_90_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_90_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_90_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_90_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_90_clock; // @[Decoupled.scala 361:21]
  wire  last_q_90_reset; // @[Decoupled.scala 361:21]
  wire  last_q_90_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_90_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_90_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_90_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_90_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_90_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_91_clock; // @[Stab.scala 175:24]
  wire  last_merger_91_reset; // @[Stab.scala 175:24]
  wire  last_merger_91_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_91_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_91_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_91_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_91_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_91_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_91_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_91_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_91_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_91_clock; // @[Decoupled.scala 361:21]
  wire  last_q_91_reset; // @[Decoupled.scala 361:21]
  wire  last_q_91_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_91_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_91_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_91_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_91_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_91_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_92_clock; // @[Stab.scala 175:24]
  wire  last_merger_92_reset; // @[Stab.scala 175:24]
  wire  last_merger_92_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_92_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_92_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_92_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_92_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_92_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_92_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_92_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_92_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_92_clock; // @[Decoupled.scala 361:21]
  wire  last_q_92_reset; // @[Decoupled.scala 361:21]
  wire  last_q_92_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_92_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_92_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_92_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_92_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_92_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_93_clock; // @[Stab.scala 175:24]
  wire  last_merger_93_reset; // @[Stab.scala 175:24]
  wire  last_merger_93_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_93_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_93_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_93_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_93_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_93_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_93_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_93_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_93_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_93_clock; // @[Decoupled.scala 361:21]
  wire  last_q_93_reset; // @[Decoupled.scala 361:21]
  wire  last_q_93_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_93_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_93_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_93_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_93_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_93_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_94_clock; // @[Stab.scala 175:24]
  wire  last_merger_94_reset; // @[Stab.scala 175:24]
  wire  last_merger_94_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_94_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_94_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_94_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_94_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_94_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_94_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_94_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_94_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_94_clock; // @[Decoupled.scala 361:21]
  wire  last_q_94_reset; // @[Decoupled.scala 361:21]
  wire  last_q_94_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_94_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_94_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_94_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_94_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_94_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_95_clock; // @[Stab.scala 175:24]
  wire  last_merger_95_reset; // @[Stab.scala 175:24]
  wire  last_merger_95_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_95_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_95_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_95_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_95_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_95_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_95_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_95_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_95_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_95_clock; // @[Decoupled.scala 361:21]
  wire  last_q_95_reset; // @[Decoupled.scala 361:21]
  wire  last_q_95_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_95_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_95_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_95_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_95_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_95_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_96_clock; // @[Stab.scala 175:24]
  wire  last_merger_96_reset; // @[Stab.scala 175:24]
  wire  last_merger_96_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_96_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_96_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_96_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_96_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_96_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_96_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_96_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_96_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_96_clock; // @[Decoupled.scala 361:21]
  wire  last_q_96_reset; // @[Decoupled.scala 361:21]
  wire  last_q_96_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_96_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_96_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_96_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_96_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_96_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_97_clock; // @[Stab.scala 175:24]
  wire  last_merger_97_reset; // @[Stab.scala 175:24]
  wire  last_merger_97_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_97_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_97_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_97_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_97_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_97_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_97_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_97_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_97_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_97_clock; // @[Decoupled.scala 361:21]
  wire  last_q_97_reset; // @[Decoupled.scala 361:21]
  wire  last_q_97_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_97_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_97_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_97_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_97_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_97_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_98_clock; // @[Stab.scala 175:24]
  wire  last_merger_98_reset; // @[Stab.scala 175:24]
  wire  last_merger_98_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_98_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_98_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_98_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_98_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_98_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_98_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_98_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_98_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_98_clock; // @[Decoupled.scala 361:21]
  wire  last_q_98_reset; // @[Decoupled.scala 361:21]
  wire  last_q_98_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_98_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_98_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_98_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_98_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_98_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_99_clock; // @[Stab.scala 175:24]
  wire  last_merger_99_reset; // @[Stab.scala 175:24]
  wire  last_merger_99_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_99_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_99_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_99_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_99_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_99_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_99_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_99_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_99_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_99_clock; // @[Decoupled.scala 361:21]
  wire  last_q_99_reset; // @[Decoupled.scala 361:21]
  wire  last_q_99_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_99_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_99_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_99_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_99_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_99_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_100_clock; // @[Stab.scala 175:24]
  wire  last_merger_100_reset; // @[Stab.scala 175:24]
  wire  last_merger_100_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_100_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_100_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_100_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_100_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_100_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_100_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_100_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_100_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_100_clock; // @[Decoupled.scala 361:21]
  wire  last_q_100_reset; // @[Decoupled.scala 361:21]
  wire  last_q_100_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_100_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_100_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_100_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_100_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_100_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_101_clock; // @[Stab.scala 175:24]
  wire  last_merger_101_reset; // @[Stab.scala 175:24]
  wire  last_merger_101_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_101_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_101_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_101_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_101_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_101_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_101_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_101_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_101_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_101_clock; // @[Decoupled.scala 361:21]
  wire  last_q_101_reset; // @[Decoupled.scala 361:21]
  wire  last_q_101_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_101_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_101_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_101_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_101_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_101_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_102_clock; // @[Stab.scala 175:24]
  wire  last_merger_102_reset; // @[Stab.scala 175:24]
  wire  last_merger_102_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_102_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_102_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_102_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_102_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_102_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_102_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_102_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_102_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_102_clock; // @[Decoupled.scala 361:21]
  wire  last_q_102_reset; // @[Decoupled.scala 361:21]
  wire  last_q_102_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_102_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_102_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_102_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_102_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_102_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_103_clock; // @[Stab.scala 175:24]
  wire  last_merger_103_reset; // @[Stab.scala 175:24]
  wire  last_merger_103_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_103_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_103_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_103_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_103_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_103_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_103_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_103_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_103_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_103_clock; // @[Decoupled.scala 361:21]
  wire  last_q_103_reset; // @[Decoupled.scala 361:21]
  wire  last_q_103_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_103_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_103_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_103_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_103_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_103_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_104_clock; // @[Stab.scala 175:24]
  wire  last_merger_104_reset; // @[Stab.scala 175:24]
  wire  last_merger_104_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_104_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_104_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_104_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_104_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_104_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_104_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_104_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_104_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_104_clock; // @[Decoupled.scala 361:21]
  wire  last_q_104_reset; // @[Decoupled.scala 361:21]
  wire  last_q_104_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_104_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_104_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_104_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_104_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_104_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_105_clock; // @[Stab.scala 175:24]
  wire  last_merger_105_reset; // @[Stab.scala 175:24]
  wire  last_merger_105_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_105_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_105_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_105_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_105_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_105_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_105_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_105_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_105_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_105_clock; // @[Decoupled.scala 361:21]
  wire  last_q_105_reset; // @[Decoupled.scala 361:21]
  wire  last_q_105_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_105_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_105_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_105_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_105_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_105_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_106_clock; // @[Stab.scala 175:24]
  wire  last_merger_106_reset; // @[Stab.scala 175:24]
  wire  last_merger_106_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_106_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_106_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_106_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_106_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_106_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_106_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_106_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_106_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_106_clock; // @[Decoupled.scala 361:21]
  wire  last_q_106_reset; // @[Decoupled.scala 361:21]
  wire  last_q_106_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_106_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_106_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_106_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_106_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_106_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_107_clock; // @[Stab.scala 175:24]
  wire  last_merger_107_reset; // @[Stab.scala 175:24]
  wire  last_merger_107_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_107_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_107_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_107_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_107_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_107_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_107_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_107_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_107_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_107_clock; // @[Decoupled.scala 361:21]
  wire  last_q_107_reset; // @[Decoupled.scala 361:21]
  wire  last_q_107_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_107_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_107_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_107_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_107_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_107_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_108_clock; // @[Stab.scala 175:24]
  wire  last_merger_108_reset; // @[Stab.scala 175:24]
  wire  last_merger_108_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_108_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_108_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_108_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_108_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_108_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_108_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_108_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_108_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_108_clock; // @[Decoupled.scala 361:21]
  wire  last_q_108_reset; // @[Decoupled.scala 361:21]
  wire  last_q_108_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_108_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_108_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_108_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_108_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_108_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_109_clock; // @[Stab.scala 175:24]
  wire  last_merger_109_reset; // @[Stab.scala 175:24]
  wire  last_merger_109_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_109_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_109_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_109_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_109_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_109_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_109_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_109_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_109_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_109_clock; // @[Decoupled.scala 361:21]
  wire  last_q_109_reset; // @[Decoupled.scala 361:21]
  wire  last_q_109_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_109_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_109_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_109_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_109_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_109_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_110_clock; // @[Stab.scala 175:24]
  wire  last_merger_110_reset; // @[Stab.scala 175:24]
  wire  last_merger_110_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_110_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_110_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_110_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_110_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_110_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_110_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_110_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_110_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_110_clock; // @[Decoupled.scala 361:21]
  wire  last_q_110_reset; // @[Decoupled.scala 361:21]
  wire  last_q_110_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_110_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_110_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_110_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_110_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_110_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_111_clock; // @[Stab.scala 175:24]
  wire  last_merger_111_reset; // @[Stab.scala 175:24]
  wire  last_merger_111_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_111_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_111_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_111_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_111_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_111_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_111_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_111_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_111_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_111_clock; // @[Decoupled.scala 361:21]
  wire  last_q_111_reset; // @[Decoupled.scala 361:21]
  wire  last_q_111_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_111_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_111_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_111_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_111_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_111_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_112_clock; // @[Stab.scala 175:24]
  wire  last_merger_112_reset; // @[Stab.scala 175:24]
  wire  last_merger_112_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_112_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_112_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_112_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_112_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_112_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_112_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_112_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_112_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_112_clock; // @[Decoupled.scala 361:21]
  wire  last_q_112_reset; // @[Decoupled.scala 361:21]
  wire  last_q_112_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_112_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_112_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_112_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_112_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_112_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_113_clock; // @[Stab.scala 175:24]
  wire  last_merger_113_reset; // @[Stab.scala 175:24]
  wire  last_merger_113_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_113_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_113_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_113_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_113_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_113_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_113_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_113_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_113_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_113_clock; // @[Decoupled.scala 361:21]
  wire  last_q_113_reset; // @[Decoupled.scala 361:21]
  wire  last_q_113_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_113_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_113_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_113_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_113_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_113_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_114_clock; // @[Stab.scala 175:24]
  wire  last_merger_114_reset; // @[Stab.scala 175:24]
  wire  last_merger_114_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_114_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_114_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_114_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_114_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_114_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_114_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_114_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_114_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_114_clock; // @[Decoupled.scala 361:21]
  wire  last_q_114_reset; // @[Decoupled.scala 361:21]
  wire  last_q_114_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_114_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_114_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_114_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_114_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_114_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_115_clock; // @[Stab.scala 175:24]
  wire  last_merger_115_reset; // @[Stab.scala 175:24]
  wire  last_merger_115_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_115_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_115_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_115_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_115_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_115_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_115_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_115_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_115_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_115_clock; // @[Decoupled.scala 361:21]
  wire  last_q_115_reset; // @[Decoupled.scala 361:21]
  wire  last_q_115_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_115_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_115_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_115_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_115_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_115_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_116_clock; // @[Stab.scala 175:24]
  wire  last_merger_116_reset; // @[Stab.scala 175:24]
  wire  last_merger_116_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_116_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_116_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_116_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_116_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_116_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_116_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_116_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_116_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_116_clock; // @[Decoupled.scala 361:21]
  wire  last_q_116_reset; // @[Decoupled.scala 361:21]
  wire  last_q_116_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_116_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_116_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_116_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_116_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_116_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_117_clock; // @[Stab.scala 175:24]
  wire  last_merger_117_reset; // @[Stab.scala 175:24]
  wire  last_merger_117_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_117_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_117_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_117_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_117_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_117_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_117_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_117_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_117_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_117_clock; // @[Decoupled.scala 361:21]
  wire  last_q_117_reset; // @[Decoupled.scala 361:21]
  wire  last_q_117_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_117_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_117_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_117_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_117_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_117_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_118_clock; // @[Stab.scala 175:24]
  wire  last_merger_118_reset; // @[Stab.scala 175:24]
  wire  last_merger_118_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_118_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_118_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_118_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_118_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_118_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_118_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_118_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_118_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_118_clock; // @[Decoupled.scala 361:21]
  wire  last_q_118_reset; // @[Decoupled.scala 361:21]
  wire  last_q_118_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_118_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_118_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_118_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_118_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_118_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_119_clock; // @[Stab.scala 175:24]
  wire  last_merger_119_reset; // @[Stab.scala 175:24]
  wire  last_merger_119_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_119_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_119_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_119_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_119_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_119_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_119_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_119_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_119_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_119_clock; // @[Decoupled.scala 361:21]
  wire  last_q_119_reset; // @[Decoupled.scala 361:21]
  wire  last_q_119_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_119_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_119_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_119_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_119_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_119_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_120_clock; // @[Stab.scala 175:24]
  wire  last_merger_120_reset; // @[Stab.scala 175:24]
  wire  last_merger_120_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_120_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_120_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_120_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_120_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_120_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_120_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_120_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_120_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_120_clock; // @[Decoupled.scala 361:21]
  wire  last_q_120_reset; // @[Decoupled.scala 361:21]
  wire  last_q_120_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_120_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_120_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_120_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_120_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_120_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_121_clock; // @[Stab.scala 175:24]
  wire  last_merger_121_reset; // @[Stab.scala 175:24]
  wire  last_merger_121_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_121_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_121_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_121_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_121_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_121_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_121_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_121_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_121_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_121_clock; // @[Decoupled.scala 361:21]
  wire  last_q_121_reset; // @[Decoupled.scala 361:21]
  wire  last_q_121_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_121_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_121_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_121_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_121_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_121_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_122_clock; // @[Stab.scala 175:24]
  wire  last_merger_122_reset; // @[Stab.scala 175:24]
  wire  last_merger_122_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_122_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_122_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_122_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_122_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_122_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_122_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_122_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_122_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_122_clock; // @[Decoupled.scala 361:21]
  wire  last_q_122_reset; // @[Decoupled.scala 361:21]
  wire  last_q_122_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_122_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_122_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_122_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_122_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_122_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_123_clock; // @[Stab.scala 175:24]
  wire  last_merger_123_reset; // @[Stab.scala 175:24]
  wire  last_merger_123_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_123_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_123_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_123_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_123_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_123_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_123_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_123_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_123_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_123_clock; // @[Decoupled.scala 361:21]
  wire  last_q_123_reset; // @[Decoupled.scala 361:21]
  wire  last_q_123_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_123_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_123_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_123_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_123_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_123_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_124_clock; // @[Stab.scala 175:24]
  wire  last_merger_124_reset; // @[Stab.scala 175:24]
  wire  last_merger_124_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_124_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_124_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_124_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_124_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_124_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_124_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_124_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_124_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_124_clock; // @[Decoupled.scala 361:21]
  wire  last_q_124_reset; // @[Decoupled.scala 361:21]
  wire  last_q_124_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_124_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_124_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_124_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_124_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_124_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_125_clock; // @[Stab.scala 175:24]
  wire  last_merger_125_reset; // @[Stab.scala 175:24]
  wire  last_merger_125_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_125_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_125_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_125_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_125_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_125_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_125_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_125_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_125_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_125_clock; // @[Decoupled.scala 361:21]
  wire  last_q_125_reset; // @[Decoupled.scala 361:21]
  wire  last_q_125_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_125_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_125_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_125_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_125_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_125_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_126_clock; // @[Stab.scala 175:24]
  wire  last_merger_126_reset; // @[Stab.scala 175:24]
  wire  last_merger_126_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_126_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_126_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_126_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_126_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_126_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_126_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_126_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_126_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_126_clock; // @[Decoupled.scala 361:21]
  wire  last_q_126_reset; // @[Decoupled.scala 361:21]
  wire  last_q_126_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_126_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_126_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_126_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_126_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_126_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_127_clock; // @[Stab.scala 175:24]
  wire  last_merger_127_reset; // @[Stab.scala 175:24]
  wire  last_merger_127_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_127_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_127_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_127_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_127_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_127_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_127_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_127_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_127_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_127_clock; // @[Decoupled.scala 361:21]
  wire  last_q_127_reset; // @[Decoupled.scala 361:21]
  wire  last_q_127_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_127_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_127_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_127_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_127_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_127_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_128_clock; // @[Stab.scala 175:24]
  wire  last_merger_128_reset; // @[Stab.scala 175:24]
  wire  last_merger_128_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_128_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_128_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_128_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_128_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_128_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_128_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_128_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_128_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_128_clock; // @[Decoupled.scala 361:21]
  wire  last_q_128_reset; // @[Decoupled.scala 361:21]
  wire  last_q_128_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_128_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_128_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_128_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_128_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_128_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_129_clock; // @[Stab.scala 175:24]
  wire  last_merger_129_reset; // @[Stab.scala 175:24]
  wire  last_merger_129_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_129_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_129_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_129_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_129_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_129_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_129_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_129_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_129_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_129_clock; // @[Decoupled.scala 361:21]
  wire  last_q_129_reset; // @[Decoupled.scala 361:21]
  wire  last_q_129_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_129_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_129_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_129_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_129_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_129_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_130_clock; // @[Stab.scala 175:24]
  wire  last_merger_130_reset; // @[Stab.scala 175:24]
  wire  last_merger_130_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_130_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_130_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_130_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_130_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_130_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_130_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_130_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_130_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_130_clock; // @[Decoupled.scala 361:21]
  wire  last_q_130_reset; // @[Decoupled.scala 361:21]
  wire  last_q_130_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_130_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_130_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_130_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_130_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_130_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_131_clock; // @[Stab.scala 175:24]
  wire  last_merger_131_reset; // @[Stab.scala 175:24]
  wire  last_merger_131_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_131_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_131_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_131_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_131_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_131_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_131_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_131_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_131_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_131_clock; // @[Decoupled.scala 361:21]
  wire  last_q_131_reset; // @[Decoupled.scala 361:21]
  wire  last_q_131_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_131_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_131_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_131_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_131_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_131_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_132_clock; // @[Stab.scala 175:24]
  wire  last_merger_132_reset; // @[Stab.scala 175:24]
  wire  last_merger_132_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_132_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_132_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_132_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_132_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_132_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_132_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_132_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_132_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_132_clock; // @[Decoupled.scala 361:21]
  wire  last_q_132_reset; // @[Decoupled.scala 361:21]
  wire  last_q_132_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_132_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_132_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_132_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_132_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_132_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_133_clock; // @[Stab.scala 175:24]
  wire  last_merger_133_reset; // @[Stab.scala 175:24]
  wire  last_merger_133_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_133_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_133_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_133_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_133_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_133_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_133_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_133_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_133_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_133_clock; // @[Decoupled.scala 361:21]
  wire  last_q_133_reset; // @[Decoupled.scala 361:21]
  wire  last_q_133_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_133_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_133_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_133_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_133_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_133_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_134_clock; // @[Stab.scala 175:24]
  wire  last_merger_134_reset; // @[Stab.scala 175:24]
  wire  last_merger_134_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_134_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_134_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_134_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_134_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_134_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_134_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_134_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_134_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_134_clock; // @[Decoupled.scala 361:21]
  wire  last_q_134_reset; // @[Decoupled.scala 361:21]
  wire  last_q_134_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_134_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_134_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_134_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_134_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_134_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_135_clock; // @[Stab.scala 175:24]
  wire  last_merger_135_reset; // @[Stab.scala 175:24]
  wire  last_merger_135_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_135_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_135_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_135_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_135_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_135_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_135_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_135_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_135_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_135_clock; // @[Decoupled.scala 361:21]
  wire  last_q_135_reset; // @[Decoupled.scala 361:21]
  wire  last_q_135_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_135_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_135_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_135_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_135_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_135_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_136_clock; // @[Stab.scala 175:24]
  wire  last_merger_136_reset; // @[Stab.scala 175:24]
  wire  last_merger_136_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_136_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_136_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_136_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_136_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_136_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_136_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_136_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_136_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_136_clock; // @[Decoupled.scala 361:21]
  wire  last_q_136_reset; // @[Decoupled.scala 361:21]
  wire  last_q_136_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_136_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_136_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_136_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_136_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_136_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_137_clock; // @[Stab.scala 175:24]
  wire  last_merger_137_reset; // @[Stab.scala 175:24]
  wire  last_merger_137_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_137_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_137_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_137_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_137_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_137_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_137_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_137_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_137_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_137_clock; // @[Decoupled.scala 361:21]
  wire  last_q_137_reset; // @[Decoupled.scala 361:21]
  wire  last_q_137_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_137_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_137_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_137_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_137_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_137_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_138_clock; // @[Stab.scala 175:24]
  wire  last_merger_138_reset; // @[Stab.scala 175:24]
  wire  last_merger_138_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_138_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_138_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_138_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_138_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_138_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_138_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_138_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_138_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_138_clock; // @[Decoupled.scala 361:21]
  wire  last_q_138_reset; // @[Decoupled.scala 361:21]
  wire  last_q_138_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_138_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_138_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_138_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_138_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_138_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_139_clock; // @[Stab.scala 175:24]
  wire  last_merger_139_reset; // @[Stab.scala 175:24]
  wire  last_merger_139_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_139_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_139_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_139_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_139_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_139_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_139_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_139_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_139_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_139_clock; // @[Decoupled.scala 361:21]
  wire  last_q_139_reset; // @[Decoupled.scala 361:21]
  wire  last_q_139_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_139_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_139_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_139_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_139_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_139_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_140_clock; // @[Stab.scala 175:24]
  wire  last_merger_140_reset; // @[Stab.scala 175:24]
  wire  last_merger_140_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_140_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_140_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_140_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_140_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_140_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_140_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_140_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_140_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_140_clock; // @[Decoupled.scala 361:21]
  wire  last_q_140_reset; // @[Decoupled.scala 361:21]
  wire  last_q_140_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_140_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_140_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_140_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_140_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_140_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_141_clock; // @[Stab.scala 175:24]
  wire  last_merger_141_reset; // @[Stab.scala 175:24]
  wire  last_merger_141_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_141_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_141_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_141_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_141_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_141_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_141_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_141_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_141_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_141_clock; // @[Decoupled.scala 361:21]
  wire  last_q_141_reset; // @[Decoupled.scala 361:21]
  wire  last_q_141_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_141_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_141_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_141_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_141_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_141_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_142_clock; // @[Stab.scala 175:24]
  wire  last_merger_142_reset; // @[Stab.scala 175:24]
  wire  last_merger_142_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_142_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_142_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_142_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_142_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_142_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_142_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_142_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_142_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_142_clock; // @[Decoupled.scala 361:21]
  wire  last_q_142_reset; // @[Decoupled.scala 361:21]
  wire  last_q_142_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_142_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_142_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_142_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_142_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_142_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_143_clock; // @[Stab.scala 175:24]
  wire  last_merger_143_reset; // @[Stab.scala 175:24]
  wire  last_merger_143_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_143_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_143_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_143_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_143_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_143_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_143_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_143_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_143_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_143_clock; // @[Decoupled.scala 361:21]
  wire  last_q_143_reset; // @[Decoupled.scala 361:21]
  wire  last_q_143_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_143_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_143_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_143_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_143_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_143_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_144_clock; // @[Stab.scala 175:24]
  wire  last_merger_144_reset; // @[Stab.scala 175:24]
  wire  last_merger_144_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_144_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_144_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_144_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_144_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_144_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_144_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_144_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_144_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_144_clock; // @[Decoupled.scala 361:21]
  wire  last_q_144_reset; // @[Decoupled.scala 361:21]
  wire  last_q_144_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_144_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_144_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_144_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_144_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_144_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_145_clock; // @[Stab.scala 175:24]
  wire  last_merger_145_reset; // @[Stab.scala 175:24]
  wire  last_merger_145_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_145_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_145_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_145_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_145_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_145_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_145_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_145_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_145_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_145_clock; // @[Decoupled.scala 361:21]
  wire  last_q_145_reset; // @[Decoupled.scala 361:21]
  wire  last_q_145_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_145_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_145_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_145_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_145_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_145_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_146_clock; // @[Stab.scala 175:24]
  wire  last_merger_146_reset; // @[Stab.scala 175:24]
  wire  last_merger_146_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_146_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_146_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_146_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_146_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_146_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_146_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_146_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_146_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_146_clock; // @[Decoupled.scala 361:21]
  wire  last_q_146_reset; // @[Decoupled.scala 361:21]
  wire  last_q_146_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_146_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_146_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_146_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_146_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_146_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_147_clock; // @[Stab.scala 175:24]
  wire  last_merger_147_reset; // @[Stab.scala 175:24]
  wire  last_merger_147_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_147_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_147_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_147_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_147_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_147_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_147_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_147_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_147_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_147_clock; // @[Decoupled.scala 361:21]
  wire  last_q_147_reset; // @[Decoupled.scala 361:21]
  wire  last_q_147_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_147_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_147_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_147_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_147_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_147_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_148_clock; // @[Stab.scala 175:24]
  wire  last_merger_148_reset; // @[Stab.scala 175:24]
  wire  last_merger_148_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_148_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_148_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_148_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_148_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_148_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_148_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_148_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_148_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_148_clock; // @[Decoupled.scala 361:21]
  wire  last_q_148_reset; // @[Decoupled.scala 361:21]
  wire  last_q_148_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_148_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_148_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_148_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_148_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_148_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_149_clock; // @[Stab.scala 175:24]
  wire  last_merger_149_reset; // @[Stab.scala 175:24]
  wire  last_merger_149_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_149_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_149_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_149_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_149_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_149_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_149_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_149_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_149_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_149_clock; // @[Decoupled.scala 361:21]
  wire  last_q_149_reset; // @[Decoupled.scala 361:21]
  wire  last_q_149_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_149_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_149_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_149_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_149_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_149_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_150_clock; // @[Stab.scala 175:24]
  wire  last_merger_150_reset; // @[Stab.scala 175:24]
  wire  last_merger_150_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_150_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_150_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_150_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_150_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_150_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_150_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_150_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_150_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_150_clock; // @[Decoupled.scala 361:21]
  wire  last_q_150_reset; // @[Decoupled.scala 361:21]
  wire  last_q_150_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_150_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_150_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_150_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_150_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_150_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_151_clock; // @[Stab.scala 175:24]
  wire  last_merger_151_reset; // @[Stab.scala 175:24]
  wire  last_merger_151_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_151_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_151_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_151_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_151_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_151_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_151_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_151_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_151_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_151_clock; // @[Decoupled.scala 361:21]
  wire  last_q_151_reset; // @[Decoupled.scala 361:21]
  wire  last_q_151_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_151_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_151_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_151_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_151_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_151_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_152_clock; // @[Stab.scala 175:24]
  wire  last_merger_152_reset; // @[Stab.scala 175:24]
  wire  last_merger_152_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_152_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_152_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_152_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_152_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_152_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_152_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_152_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_152_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_152_clock; // @[Decoupled.scala 361:21]
  wire  last_q_152_reset; // @[Decoupled.scala 361:21]
  wire  last_q_152_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_152_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_152_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_152_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_152_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_152_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_153_clock; // @[Stab.scala 175:24]
  wire  last_merger_153_reset; // @[Stab.scala 175:24]
  wire  last_merger_153_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_153_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_153_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_153_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_153_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_153_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_153_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_153_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_153_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_153_clock; // @[Decoupled.scala 361:21]
  wire  last_q_153_reset; // @[Decoupled.scala 361:21]
  wire  last_q_153_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_153_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_153_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_153_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_153_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_153_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_154_clock; // @[Stab.scala 175:24]
  wire  last_merger_154_reset; // @[Stab.scala 175:24]
  wire  last_merger_154_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_154_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_154_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_154_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_154_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_154_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_154_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_154_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_154_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_154_clock; // @[Decoupled.scala 361:21]
  wire  last_q_154_reset; // @[Decoupled.scala 361:21]
  wire  last_q_154_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_154_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_154_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_154_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_154_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_154_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_155_clock; // @[Stab.scala 175:24]
  wire  last_merger_155_reset; // @[Stab.scala 175:24]
  wire  last_merger_155_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_155_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_155_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_155_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_155_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_155_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_155_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_155_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_155_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_155_clock; // @[Decoupled.scala 361:21]
  wire  last_q_155_reset; // @[Decoupled.scala 361:21]
  wire  last_q_155_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_155_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_155_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_155_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_155_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_155_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_156_clock; // @[Stab.scala 175:24]
  wire  last_merger_156_reset; // @[Stab.scala 175:24]
  wire  last_merger_156_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_156_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_156_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_156_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_156_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_156_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_156_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_156_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_156_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_156_clock; // @[Decoupled.scala 361:21]
  wire  last_q_156_reset; // @[Decoupled.scala 361:21]
  wire  last_q_156_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_156_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_156_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_156_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_156_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_156_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_157_clock; // @[Stab.scala 175:24]
  wire  last_merger_157_reset; // @[Stab.scala 175:24]
  wire  last_merger_157_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_157_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_157_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_157_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_157_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_157_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_157_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_157_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_157_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_157_clock; // @[Decoupled.scala 361:21]
  wire  last_q_157_reset; // @[Decoupled.scala 361:21]
  wire  last_q_157_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_157_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_157_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_157_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_157_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_157_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_158_clock; // @[Stab.scala 175:24]
  wire  last_merger_158_reset; // @[Stab.scala 175:24]
  wire  last_merger_158_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_158_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_158_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_158_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_158_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_158_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_158_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_158_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_158_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_158_clock; // @[Decoupled.scala 361:21]
  wire  last_q_158_reset; // @[Decoupled.scala 361:21]
  wire  last_q_158_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_158_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_158_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_158_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_158_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_158_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_159_clock; // @[Stab.scala 175:24]
  wire  last_merger_159_reset; // @[Stab.scala 175:24]
  wire  last_merger_159_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_159_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_159_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_159_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_159_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_159_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_159_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_159_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_159_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_159_clock; // @[Decoupled.scala 361:21]
  wire  last_q_159_reset; // @[Decoupled.scala 361:21]
  wire  last_q_159_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_159_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_159_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_159_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_159_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_159_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_160_clock; // @[Stab.scala 175:24]
  wire  last_merger_160_reset; // @[Stab.scala 175:24]
  wire  last_merger_160_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_160_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_160_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_160_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_160_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_160_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_160_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_160_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_160_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_160_clock; // @[Decoupled.scala 361:21]
  wire  last_q_160_reset; // @[Decoupled.scala 361:21]
  wire  last_q_160_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_160_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_160_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_160_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_160_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_160_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_161_clock; // @[Stab.scala 175:24]
  wire  last_merger_161_reset; // @[Stab.scala 175:24]
  wire  last_merger_161_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_161_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_161_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_161_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_161_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_161_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_161_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_161_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_161_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_161_clock; // @[Decoupled.scala 361:21]
  wire  last_q_161_reset; // @[Decoupled.scala 361:21]
  wire  last_q_161_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_161_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_161_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_161_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_161_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_161_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_162_clock; // @[Stab.scala 175:24]
  wire  last_merger_162_reset; // @[Stab.scala 175:24]
  wire  last_merger_162_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_162_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_162_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_162_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_162_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_162_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_162_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_162_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_162_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_162_clock; // @[Decoupled.scala 361:21]
  wire  last_q_162_reset; // @[Decoupled.scala 361:21]
  wire  last_q_162_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_162_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_162_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_162_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_162_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_162_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_163_clock; // @[Stab.scala 175:24]
  wire  last_merger_163_reset; // @[Stab.scala 175:24]
  wire  last_merger_163_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_163_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_163_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_163_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_163_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_163_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_163_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_163_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_163_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_163_clock; // @[Decoupled.scala 361:21]
  wire  last_q_163_reset; // @[Decoupled.scala 361:21]
  wire  last_q_163_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_163_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_163_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_163_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_163_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_163_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_164_clock; // @[Stab.scala 175:24]
  wire  last_merger_164_reset; // @[Stab.scala 175:24]
  wire  last_merger_164_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_164_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_164_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_164_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_164_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_164_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_164_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_164_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_164_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_164_clock; // @[Decoupled.scala 361:21]
  wire  last_q_164_reset; // @[Decoupled.scala 361:21]
  wire  last_q_164_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_164_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_164_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_164_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_164_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_164_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_165_clock; // @[Stab.scala 175:24]
  wire  last_merger_165_reset; // @[Stab.scala 175:24]
  wire  last_merger_165_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_165_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_165_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_165_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_165_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_165_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_165_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_165_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_165_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_165_clock; // @[Decoupled.scala 361:21]
  wire  last_q_165_reset; // @[Decoupled.scala 361:21]
  wire  last_q_165_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_165_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_165_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_165_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_165_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_165_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_166_clock; // @[Stab.scala 175:24]
  wire  last_merger_166_reset; // @[Stab.scala 175:24]
  wire  last_merger_166_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_166_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_166_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_166_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_166_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_166_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_166_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_166_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_166_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_166_clock; // @[Decoupled.scala 361:21]
  wire  last_q_166_reset; // @[Decoupled.scala 361:21]
  wire  last_q_166_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_166_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_166_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_166_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_166_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_166_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_167_clock; // @[Stab.scala 175:24]
  wire  last_merger_167_reset; // @[Stab.scala 175:24]
  wire  last_merger_167_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_167_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_167_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_167_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_167_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_167_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_167_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_167_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_167_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_167_clock; // @[Decoupled.scala 361:21]
  wire  last_q_167_reset; // @[Decoupled.scala 361:21]
  wire  last_q_167_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_167_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_167_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_167_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_167_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_167_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_168_clock; // @[Stab.scala 175:24]
  wire  last_merger_168_reset; // @[Stab.scala 175:24]
  wire  last_merger_168_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_168_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_168_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_168_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_168_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_168_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_168_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_168_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_168_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_168_clock; // @[Decoupled.scala 361:21]
  wire  last_q_168_reset; // @[Decoupled.scala 361:21]
  wire  last_q_168_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_168_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_168_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_168_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_168_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_168_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_169_clock; // @[Stab.scala 175:24]
  wire  last_merger_169_reset; // @[Stab.scala 175:24]
  wire  last_merger_169_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_169_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_169_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_169_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_169_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_169_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_169_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_169_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_169_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_169_clock; // @[Decoupled.scala 361:21]
  wire  last_q_169_reset; // @[Decoupled.scala 361:21]
  wire  last_q_169_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_169_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_169_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_169_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_169_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_169_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_170_clock; // @[Stab.scala 175:24]
  wire  last_merger_170_reset; // @[Stab.scala 175:24]
  wire  last_merger_170_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_170_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_170_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_170_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_170_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_170_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_170_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_170_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_170_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_170_clock; // @[Decoupled.scala 361:21]
  wire  last_q_170_reset; // @[Decoupled.scala 361:21]
  wire  last_q_170_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_170_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_170_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_170_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_170_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_170_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_171_clock; // @[Stab.scala 175:24]
  wire  last_merger_171_reset; // @[Stab.scala 175:24]
  wire  last_merger_171_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_171_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_171_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_171_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_171_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_171_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_171_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_171_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_171_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_171_clock; // @[Decoupled.scala 361:21]
  wire  last_q_171_reset; // @[Decoupled.scala 361:21]
  wire  last_q_171_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_171_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_171_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_171_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_171_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_171_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_172_clock; // @[Stab.scala 175:24]
  wire  last_merger_172_reset; // @[Stab.scala 175:24]
  wire  last_merger_172_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_172_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_172_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_172_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_172_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_172_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_172_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_172_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_172_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_172_clock; // @[Decoupled.scala 361:21]
  wire  last_q_172_reset; // @[Decoupled.scala 361:21]
  wire  last_q_172_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_172_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_172_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_172_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_172_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_172_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_173_clock; // @[Stab.scala 175:24]
  wire  last_merger_173_reset; // @[Stab.scala 175:24]
  wire  last_merger_173_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_173_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_173_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_173_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_173_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_173_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_173_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_173_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_173_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_173_clock; // @[Decoupled.scala 361:21]
  wire  last_q_173_reset; // @[Decoupled.scala 361:21]
  wire  last_q_173_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_173_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_173_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_173_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_173_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_173_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_174_clock; // @[Stab.scala 175:24]
  wire  last_merger_174_reset; // @[Stab.scala 175:24]
  wire  last_merger_174_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_174_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_174_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_174_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_174_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_174_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_174_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_174_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_174_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_174_clock; // @[Decoupled.scala 361:21]
  wire  last_q_174_reset; // @[Decoupled.scala 361:21]
  wire  last_q_174_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_174_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_174_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_174_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_174_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_174_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_175_clock; // @[Stab.scala 175:24]
  wire  last_merger_175_reset; // @[Stab.scala 175:24]
  wire  last_merger_175_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_175_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_175_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_175_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_175_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_175_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_175_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_175_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_175_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_175_clock; // @[Decoupled.scala 361:21]
  wire  last_q_175_reset; // @[Decoupled.scala 361:21]
  wire  last_q_175_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_175_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_175_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_175_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_175_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_175_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_176_clock; // @[Stab.scala 175:24]
  wire  last_merger_176_reset; // @[Stab.scala 175:24]
  wire  last_merger_176_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_176_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_176_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_176_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_176_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_176_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_176_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_176_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_176_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_176_clock; // @[Decoupled.scala 361:21]
  wire  last_q_176_reset; // @[Decoupled.scala 361:21]
  wire  last_q_176_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_176_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_176_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_176_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_176_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_176_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_177_clock; // @[Stab.scala 175:24]
  wire  last_merger_177_reset; // @[Stab.scala 175:24]
  wire  last_merger_177_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_177_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_177_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_177_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_177_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_177_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_177_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_177_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_177_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_177_clock; // @[Decoupled.scala 361:21]
  wire  last_q_177_reset; // @[Decoupled.scala 361:21]
  wire  last_q_177_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_177_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_177_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_177_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_177_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_177_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_178_clock; // @[Stab.scala 175:24]
  wire  last_merger_178_reset; // @[Stab.scala 175:24]
  wire  last_merger_178_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_178_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_178_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_178_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_178_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_178_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_178_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_178_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_178_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_178_clock; // @[Decoupled.scala 361:21]
  wire  last_q_178_reset; // @[Decoupled.scala 361:21]
  wire  last_q_178_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_178_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_178_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_178_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_178_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_178_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_179_clock; // @[Stab.scala 175:24]
  wire  last_merger_179_reset; // @[Stab.scala 175:24]
  wire  last_merger_179_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_179_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_179_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_179_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_179_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_179_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_179_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_179_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_179_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_179_clock; // @[Decoupled.scala 361:21]
  wire  last_q_179_reset; // @[Decoupled.scala 361:21]
  wire  last_q_179_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_179_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_179_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_179_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_179_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_179_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_180_clock; // @[Stab.scala 175:24]
  wire  last_merger_180_reset; // @[Stab.scala 175:24]
  wire  last_merger_180_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_180_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_180_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_180_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_180_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_180_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_180_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_180_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_180_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_180_clock; // @[Decoupled.scala 361:21]
  wire  last_q_180_reset; // @[Decoupled.scala 361:21]
  wire  last_q_180_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_180_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_180_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_180_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_180_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_180_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_181_clock; // @[Stab.scala 175:24]
  wire  last_merger_181_reset; // @[Stab.scala 175:24]
  wire  last_merger_181_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_181_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_181_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_181_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_181_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_181_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_181_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_181_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_181_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_181_clock; // @[Decoupled.scala 361:21]
  wire  last_q_181_reset; // @[Decoupled.scala 361:21]
  wire  last_q_181_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_181_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_181_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_181_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_181_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_181_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_182_clock; // @[Stab.scala 175:24]
  wire  last_merger_182_reset; // @[Stab.scala 175:24]
  wire  last_merger_182_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_182_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_182_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_182_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_182_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_182_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_182_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_182_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_182_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_182_clock; // @[Decoupled.scala 361:21]
  wire  last_q_182_reset; // @[Decoupled.scala 361:21]
  wire  last_q_182_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_182_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_182_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_182_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_182_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_182_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_183_clock; // @[Stab.scala 175:24]
  wire  last_merger_183_reset; // @[Stab.scala 175:24]
  wire  last_merger_183_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_183_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_183_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_183_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_183_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_183_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_183_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_183_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_183_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_183_clock; // @[Decoupled.scala 361:21]
  wire  last_q_183_reset; // @[Decoupled.scala 361:21]
  wire  last_q_183_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_183_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_183_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_183_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_183_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_183_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_184_clock; // @[Stab.scala 175:24]
  wire  last_merger_184_reset; // @[Stab.scala 175:24]
  wire  last_merger_184_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_184_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_184_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_184_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_184_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_184_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_184_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_184_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_184_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_184_clock; // @[Decoupled.scala 361:21]
  wire  last_q_184_reset; // @[Decoupled.scala 361:21]
  wire  last_q_184_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_184_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_184_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_184_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_184_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_184_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_185_clock; // @[Stab.scala 175:24]
  wire  last_merger_185_reset; // @[Stab.scala 175:24]
  wire  last_merger_185_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_185_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_185_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_185_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_185_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_185_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_185_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_185_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_185_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_185_clock; // @[Decoupled.scala 361:21]
  wire  last_q_185_reset; // @[Decoupled.scala 361:21]
  wire  last_q_185_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_185_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_185_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_185_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_185_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_185_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_186_clock; // @[Stab.scala 175:24]
  wire  last_merger_186_reset; // @[Stab.scala 175:24]
  wire  last_merger_186_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_186_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_186_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_186_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_186_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_186_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_186_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_186_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_186_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_186_clock; // @[Decoupled.scala 361:21]
  wire  last_q_186_reset; // @[Decoupled.scala 361:21]
  wire  last_q_186_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_186_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_186_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_186_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_186_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_186_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_187_clock; // @[Stab.scala 175:24]
  wire  last_merger_187_reset; // @[Stab.scala 175:24]
  wire  last_merger_187_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_187_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_187_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_187_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_187_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_187_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_187_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_187_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_187_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_187_clock; // @[Decoupled.scala 361:21]
  wire  last_q_187_reset; // @[Decoupled.scala 361:21]
  wire  last_q_187_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_187_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_187_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_187_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_187_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_187_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_188_clock; // @[Stab.scala 175:24]
  wire  last_merger_188_reset; // @[Stab.scala 175:24]
  wire  last_merger_188_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_188_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_188_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_188_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_188_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_188_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_188_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_188_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_188_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_188_clock; // @[Decoupled.scala 361:21]
  wire  last_q_188_reset; // @[Decoupled.scala 361:21]
  wire  last_q_188_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_188_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_188_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_188_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_188_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_188_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_189_clock; // @[Stab.scala 175:24]
  wire  last_merger_189_reset; // @[Stab.scala 175:24]
  wire  last_merger_189_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_189_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_189_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_189_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_189_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_189_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_189_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_189_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_189_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_189_clock; // @[Decoupled.scala 361:21]
  wire  last_q_189_reset; // @[Decoupled.scala 361:21]
  wire  last_q_189_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_189_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_189_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_189_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_189_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_189_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_190_clock; // @[Stab.scala 175:24]
  wire  last_merger_190_reset; // @[Stab.scala 175:24]
  wire  last_merger_190_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_190_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_190_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_190_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_190_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_190_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_190_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_190_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_190_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_190_clock; // @[Decoupled.scala 361:21]
  wire  last_q_190_reset; // @[Decoupled.scala 361:21]
  wire  last_q_190_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_190_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_190_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_190_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_190_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_190_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_191_clock; // @[Stab.scala 175:24]
  wire  last_merger_191_reset; // @[Stab.scala 175:24]
  wire  last_merger_191_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_191_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_191_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_191_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_191_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_191_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_191_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_191_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_191_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_191_clock; // @[Decoupled.scala 361:21]
  wire  last_q_191_reset; // @[Decoupled.scala 361:21]
  wire  last_q_191_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_191_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_191_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_191_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_191_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_191_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_192_clock; // @[Stab.scala 175:24]
  wire  last_merger_192_reset; // @[Stab.scala 175:24]
  wire  last_merger_192_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_192_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_192_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_192_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_192_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_192_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_192_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_192_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_192_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_192_clock; // @[Decoupled.scala 361:21]
  wire  last_q_192_reset; // @[Decoupled.scala 361:21]
  wire  last_q_192_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_192_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_192_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_192_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_192_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_192_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_193_clock; // @[Stab.scala 175:24]
  wire  last_merger_193_reset; // @[Stab.scala 175:24]
  wire  last_merger_193_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_193_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_193_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_193_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_193_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_193_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_193_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_193_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_193_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_193_clock; // @[Decoupled.scala 361:21]
  wire  last_q_193_reset; // @[Decoupled.scala 361:21]
  wire  last_q_193_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_193_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_193_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_193_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_193_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_193_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_194_clock; // @[Stab.scala 175:24]
  wire  last_merger_194_reset; // @[Stab.scala 175:24]
  wire  last_merger_194_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_194_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_194_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_194_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_194_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_194_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_194_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_194_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_194_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_194_clock; // @[Decoupled.scala 361:21]
  wire  last_q_194_reset; // @[Decoupled.scala 361:21]
  wire  last_q_194_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_194_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_194_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_194_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_194_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_194_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_195_clock; // @[Stab.scala 175:24]
  wire  last_merger_195_reset; // @[Stab.scala 175:24]
  wire  last_merger_195_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_195_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_195_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_195_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_195_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_195_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_195_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_195_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_195_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_195_clock; // @[Decoupled.scala 361:21]
  wire  last_q_195_reset; // @[Decoupled.scala 361:21]
  wire  last_q_195_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_195_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_195_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_195_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_195_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_195_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_196_clock; // @[Stab.scala 175:24]
  wire  last_merger_196_reset; // @[Stab.scala 175:24]
  wire  last_merger_196_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_196_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_196_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_196_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_196_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_196_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_196_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_196_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_196_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_196_clock; // @[Decoupled.scala 361:21]
  wire  last_q_196_reset; // @[Decoupled.scala 361:21]
  wire  last_q_196_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_196_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_196_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_196_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_196_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_196_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_197_clock; // @[Stab.scala 175:24]
  wire  last_merger_197_reset; // @[Stab.scala 175:24]
  wire  last_merger_197_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_197_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_197_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_197_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_197_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_197_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_197_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_197_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_197_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_197_clock; // @[Decoupled.scala 361:21]
  wire  last_q_197_reset; // @[Decoupled.scala 361:21]
  wire  last_q_197_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_197_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_197_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_197_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_197_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_197_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_198_clock; // @[Stab.scala 175:24]
  wire  last_merger_198_reset; // @[Stab.scala 175:24]
  wire  last_merger_198_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_198_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_198_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_198_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_198_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_198_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_198_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_198_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_198_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_198_clock; // @[Decoupled.scala 361:21]
  wire  last_q_198_reset; // @[Decoupled.scala 361:21]
  wire  last_q_198_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_198_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_198_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_198_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_198_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_198_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_199_clock; // @[Stab.scala 175:24]
  wire  last_merger_199_reset; // @[Stab.scala 175:24]
  wire  last_merger_199_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_199_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_199_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_199_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_199_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_199_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_199_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_199_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_199_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_199_clock; // @[Decoupled.scala 361:21]
  wire  last_q_199_reset; // @[Decoupled.scala 361:21]
  wire  last_q_199_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_199_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_199_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_199_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_199_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_199_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_200_clock; // @[Stab.scala 175:24]
  wire  last_merger_200_reset; // @[Stab.scala 175:24]
  wire  last_merger_200_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_200_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_200_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_200_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_200_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_200_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_200_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_200_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_200_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_200_clock; // @[Decoupled.scala 361:21]
  wire  last_q_200_reset; // @[Decoupled.scala 361:21]
  wire  last_q_200_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_200_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_200_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_200_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_200_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_200_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_201_clock; // @[Stab.scala 175:24]
  wire  last_merger_201_reset; // @[Stab.scala 175:24]
  wire  last_merger_201_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_201_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_201_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_201_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_201_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_201_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_201_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_201_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_201_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_201_clock; // @[Decoupled.scala 361:21]
  wire  last_q_201_reset; // @[Decoupled.scala 361:21]
  wire  last_q_201_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_201_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_201_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_201_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_201_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_201_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_202_clock; // @[Stab.scala 175:24]
  wire  last_merger_202_reset; // @[Stab.scala 175:24]
  wire  last_merger_202_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_202_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_202_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_202_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_202_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_202_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_202_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_202_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_202_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_202_clock; // @[Decoupled.scala 361:21]
  wire  last_q_202_reset; // @[Decoupled.scala 361:21]
  wire  last_q_202_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_202_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_202_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_202_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_202_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_202_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_203_clock; // @[Stab.scala 175:24]
  wire  last_merger_203_reset; // @[Stab.scala 175:24]
  wire  last_merger_203_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_203_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_203_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_203_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_203_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_203_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_203_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_203_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_203_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_203_clock; // @[Decoupled.scala 361:21]
  wire  last_q_203_reset; // @[Decoupled.scala 361:21]
  wire  last_q_203_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_203_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_203_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_203_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_203_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_203_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_204_clock; // @[Stab.scala 175:24]
  wire  last_merger_204_reset; // @[Stab.scala 175:24]
  wire  last_merger_204_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_204_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_204_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_204_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_204_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_204_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_204_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_204_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_204_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_204_clock; // @[Decoupled.scala 361:21]
  wire  last_q_204_reset; // @[Decoupled.scala 361:21]
  wire  last_q_204_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_204_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_204_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_204_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_204_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_204_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_205_clock; // @[Stab.scala 175:24]
  wire  last_merger_205_reset; // @[Stab.scala 175:24]
  wire  last_merger_205_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_205_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_205_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_205_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_205_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_205_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_205_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_205_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_205_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_205_clock; // @[Decoupled.scala 361:21]
  wire  last_q_205_reset; // @[Decoupled.scala 361:21]
  wire  last_q_205_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_205_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_205_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_205_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_205_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_205_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_206_clock; // @[Stab.scala 175:24]
  wire  last_merger_206_reset; // @[Stab.scala 175:24]
  wire  last_merger_206_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_206_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_206_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_206_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_206_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_206_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_206_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_206_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_206_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_206_clock; // @[Decoupled.scala 361:21]
  wire  last_q_206_reset; // @[Decoupled.scala 361:21]
  wire  last_q_206_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_206_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_206_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_206_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_206_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_206_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_207_clock; // @[Stab.scala 175:24]
  wire  last_merger_207_reset; // @[Stab.scala 175:24]
  wire  last_merger_207_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_207_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_207_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_207_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_207_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_207_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_207_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_207_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_207_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_207_clock; // @[Decoupled.scala 361:21]
  wire  last_q_207_reset; // @[Decoupled.scala 361:21]
  wire  last_q_207_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_207_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_207_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_207_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_207_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_207_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_208_clock; // @[Stab.scala 175:24]
  wire  last_merger_208_reset; // @[Stab.scala 175:24]
  wire  last_merger_208_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_208_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_208_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_208_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_208_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_208_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_208_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_208_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_208_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_208_clock; // @[Decoupled.scala 361:21]
  wire  last_q_208_reset; // @[Decoupled.scala 361:21]
  wire  last_q_208_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_208_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_208_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_208_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_208_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_208_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_209_clock; // @[Stab.scala 175:24]
  wire  last_merger_209_reset; // @[Stab.scala 175:24]
  wire  last_merger_209_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_209_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_209_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_209_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_209_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_209_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_209_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_209_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_209_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_209_clock; // @[Decoupled.scala 361:21]
  wire  last_q_209_reset; // @[Decoupled.scala 361:21]
  wire  last_q_209_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_209_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_209_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_209_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_209_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_209_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_210_clock; // @[Stab.scala 175:24]
  wire  last_merger_210_reset; // @[Stab.scala 175:24]
  wire  last_merger_210_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_210_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_210_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_210_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_210_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_210_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_210_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_210_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_210_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_210_clock; // @[Decoupled.scala 361:21]
  wire  last_q_210_reset; // @[Decoupled.scala 361:21]
  wire  last_q_210_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_210_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_210_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_210_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_210_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_210_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_211_clock; // @[Stab.scala 175:24]
  wire  last_merger_211_reset; // @[Stab.scala 175:24]
  wire  last_merger_211_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_211_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_211_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_211_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_211_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_211_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_211_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_211_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_211_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_211_clock; // @[Decoupled.scala 361:21]
  wire  last_q_211_reset; // @[Decoupled.scala 361:21]
  wire  last_q_211_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_211_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_211_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_211_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_211_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_211_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_212_clock; // @[Stab.scala 175:24]
  wire  last_merger_212_reset; // @[Stab.scala 175:24]
  wire  last_merger_212_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_212_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_212_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_212_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_212_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_212_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_212_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_212_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_212_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_212_clock; // @[Decoupled.scala 361:21]
  wire  last_q_212_reset; // @[Decoupled.scala 361:21]
  wire  last_q_212_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_212_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_212_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_212_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_212_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_212_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_213_clock; // @[Stab.scala 175:24]
  wire  last_merger_213_reset; // @[Stab.scala 175:24]
  wire  last_merger_213_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_213_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_213_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_213_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_213_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_213_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_213_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_213_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_213_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_213_clock; // @[Decoupled.scala 361:21]
  wire  last_q_213_reset; // @[Decoupled.scala 361:21]
  wire  last_q_213_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_213_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_213_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_213_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_213_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_213_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_214_clock; // @[Stab.scala 175:24]
  wire  last_merger_214_reset; // @[Stab.scala 175:24]
  wire  last_merger_214_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_214_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_214_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_214_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_214_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_214_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_214_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_214_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_214_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_214_clock; // @[Decoupled.scala 361:21]
  wire  last_q_214_reset; // @[Decoupled.scala 361:21]
  wire  last_q_214_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_214_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_214_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_214_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_214_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_214_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_215_clock; // @[Stab.scala 175:24]
  wire  last_merger_215_reset; // @[Stab.scala 175:24]
  wire  last_merger_215_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_215_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_215_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_215_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_215_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_215_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_215_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_215_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_215_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_215_clock; // @[Decoupled.scala 361:21]
  wire  last_q_215_reset; // @[Decoupled.scala 361:21]
  wire  last_q_215_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_215_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_215_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_215_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_215_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_215_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_216_clock; // @[Stab.scala 175:24]
  wire  last_merger_216_reset; // @[Stab.scala 175:24]
  wire  last_merger_216_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_216_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_216_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_216_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_216_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_216_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_216_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_216_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_216_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_216_clock; // @[Decoupled.scala 361:21]
  wire  last_q_216_reset; // @[Decoupled.scala 361:21]
  wire  last_q_216_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_216_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_216_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_216_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_216_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_216_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_217_clock; // @[Stab.scala 175:24]
  wire  last_merger_217_reset; // @[Stab.scala 175:24]
  wire  last_merger_217_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_217_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_217_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_217_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_217_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_217_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_217_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_217_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_217_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_217_clock; // @[Decoupled.scala 361:21]
  wire  last_q_217_reset; // @[Decoupled.scala 361:21]
  wire  last_q_217_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_217_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_217_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_217_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_217_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_217_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_218_clock; // @[Stab.scala 175:24]
  wire  last_merger_218_reset; // @[Stab.scala 175:24]
  wire  last_merger_218_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_218_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_218_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_218_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_218_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_218_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_218_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_218_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_218_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_218_clock; // @[Decoupled.scala 361:21]
  wire  last_q_218_reset; // @[Decoupled.scala 361:21]
  wire  last_q_218_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_218_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_218_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_218_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_218_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_218_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_219_clock; // @[Stab.scala 175:24]
  wire  last_merger_219_reset; // @[Stab.scala 175:24]
  wire  last_merger_219_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_219_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_219_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_219_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_219_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_219_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_219_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_219_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_219_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_219_clock; // @[Decoupled.scala 361:21]
  wire  last_q_219_reset; // @[Decoupled.scala 361:21]
  wire  last_q_219_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_219_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_219_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_219_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_219_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_219_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_220_clock; // @[Stab.scala 175:24]
  wire  last_merger_220_reset; // @[Stab.scala 175:24]
  wire  last_merger_220_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_220_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_220_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_220_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_220_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_220_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_220_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_220_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_220_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_220_clock; // @[Decoupled.scala 361:21]
  wire  last_q_220_reset; // @[Decoupled.scala 361:21]
  wire  last_q_220_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_220_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_220_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_220_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_220_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_220_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_221_clock; // @[Stab.scala 175:24]
  wire  last_merger_221_reset; // @[Stab.scala 175:24]
  wire  last_merger_221_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_221_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_221_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_221_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_221_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_221_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_221_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_221_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_221_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_221_clock; // @[Decoupled.scala 361:21]
  wire  last_q_221_reset; // @[Decoupled.scala 361:21]
  wire  last_q_221_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_221_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_221_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_221_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_221_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_221_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_222_clock; // @[Stab.scala 175:24]
  wire  last_merger_222_reset; // @[Stab.scala 175:24]
  wire  last_merger_222_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_222_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_222_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_222_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_222_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_222_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_222_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_222_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_222_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_222_clock; // @[Decoupled.scala 361:21]
  wire  last_q_222_reset; // @[Decoupled.scala 361:21]
  wire  last_q_222_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_222_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_222_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_222_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_222_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_222_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_223_clock; // @[Stab.scala 175:24]
  wire  last_merger_223_reset; // @[Stab.scala 175:24]
  wire  last_merger_223_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_223_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_223_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_223_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_223_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_223_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_223_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_223_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_223_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_223_clock; // @[Decoupled.scala 361:21]
  wire  last_q_223_reset; // @[Decoupled.scala 361:21]
  wire  last_q_223_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_223_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_223_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_223_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_223_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_223_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_224_clock; // @[Stab.scala 175:24]
  wire  last_merger_224_reset; // @[Stab.scala 175:24]
  wire  last_merger_224_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_224_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_224_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_224_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_224_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_224_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_224_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_224_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_224_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_224_clock; // @[Decoupled.scala 361:21]
  wire  last_q_224_reset; // @[Decoupled.scala 361:21]
  wire  last_q_224_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_224_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_224_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_224_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_224_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_224_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_225_clock; // @[Stab.scala 175:24]
  wire  last_merger_225_reset; // @[Stab.scala 175:24]
  wire  last_merger_225_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_225_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_225_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_225_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_225_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_225_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_225_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_225_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_225_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_225_clock; // @[Decoupled.scala 361:21]
  wire  last_q_225_reset; // @[Decoupled.scala 361:21]
  wire  last_q_225_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_225_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_225_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_225_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_225_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_225_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_226_clock; // @[Stab.scala 175:24]
  wire  last_merger_226_reset; // @[Stab.scala 175:24]
  wire  last_merger_226_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_226_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_226_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_226_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_226_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_226_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_226_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_226_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_226_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_226_clock; // @[Decoupled.scala 361:21]
  wire  last_q_226_reset; // @[Decoupled.scala 361:21]
  wire  last_q_226_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_226_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_226_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_226_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_226_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_226_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_227_clock; // @[Stab.scala 175:24]
  wire  last_merger_227_reset; // @[Stab.scala 175:24]
  wire  last_merger_227_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_227_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_227_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_227_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_227_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_227_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_227_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_227_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_227_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_227_clock; // @[Decoupled.scala 361:21]
  wire  last_q_227_reset; // @[Decoupled.scala 361:21]
  wire  last_q_227_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_227_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_227_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_227_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_227_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_227_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_228_clock; // @[Stab.scala 175:24]
  wire  last_merger_228_reset; // @[Stab.scala 175:24]
  wire  last_merger_228_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_228_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_228_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_228_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_228_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_228_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_228_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_228_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_228_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_228_clock; // @[Decoupled.scala 361:21]
  wire  last_q_228_reset; // @[Decoupled.scala 361:21]
  wire  last_q_228_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_228_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_228_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_228_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_228_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_228_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_229_clock; // @[Stab.scala 175:24]
  wire  last_merger_229_reset; // @[Stab.scala 175:24]
  wire  last_merger_229_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_229_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_229_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_229_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_229_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_229_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_229_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_229_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_229_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_229_clock; // @[Decoupled.scala 361:21]
  wire  last_q_229_reset; // @[Decoupled.scala 361:21]
  wire  last_q_229_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_229_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_229_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_229_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_229_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_229_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_230_clock; // @[Stab.scala 175:24]
  wire  last_merger_230_reset; // @[Stab.scala 175:24]
  wire  last_merger_230_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_230_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_230_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_230_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_230_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_230_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_230_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_230_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_230_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_230_clock; // @[Decoupled.scala 361:21]
  wire  last_q_230_reset; // @[Decoupled.scala 361:21]
  wire  last_q_230_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_230_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_230_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_230_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_230_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_230_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_231_clock; // @[Stab.scala 175:24]
  wire  last_merger_231_reset; // @[Stab.scala 175:24]
  wire  last_merger_231_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_231_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_231_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_231_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_231_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_231_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_231_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_231_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_231_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_231_clock; // @[Decoupled.scala 361:21]
  wire  last_q_231_reset; // @[Decoupled.scala 361:21]
  wire  last_q_231_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_231_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_231_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_231_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_231_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_231_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_232_clock; // @[Stab.scala 175:24]
  wire  last_merger_232_reset; // @[Stab.scala 175:24]
  wire  last_merger_232_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_232_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_232_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_232_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_232_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_232_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_232_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_232_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_232_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_232_clock; // @[Decoupled.scala 361:21]
  wire  last_q_232_reset; // @[Decoupled.scala 361:21]
  wire  last_q_232_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_232_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_232_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_232_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_232_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_232_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_233_clock; // @[Stab.scala 175:24]
  wire  last_merger_233_reset; // @[Stab.scala 175:24]
  wire  last_merger_233_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_233_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_233_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_233_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_233_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_233_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_233_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_233_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_233_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_233_clock; // @[Decoupled.scala 361:21]
  wire  last_q_233_reset; // @[Decoupled.scala 361:21]
  wire  last_q_233_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_233_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_233_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_233_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_233_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_233_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_234_clock; // @[Stab.scala 175:24]
  wire  last_merger_234_reset; // @[Stab.scala 175:24]
  wire  last_merger_234_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_234_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_234_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_234_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_234_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_234_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_234_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_234_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_234_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_234_clock; // @[Decoupled.scala 361:21]
  wire  last_q_234_reset; // @[Decoupled.scala 361:21]
  wire  last_q_234_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_234_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_234_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_234_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_234_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_234_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_235_clock; // @[Stab.scala 175:24]
  wire  last_merger_235_reset; // @[Stab.scala 175:24]
  wire  last_merger_235_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_235_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_235_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_235_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_235_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_235_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_235_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_235_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_235_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_235_clock; // @[Decoupled.scala 361:21]
  wire  last_q_235_reset; // @[Decoupled.scala 361:21]
  wire  last_q_235_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_235_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_235_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_235_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_235_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_235_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_236_clock; // @[Stab.scala 175:24]
  wire  last_merger_236_reset; // @[Stab.scala 175:24]
  wire  last_merger_236_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_236_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_236_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_236_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_236_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_236_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_236_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_236_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_236_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_236_clock; // @[Decoupled.scala 361:21]
  wire  last_q_236_reset; // @[Decoupled.scala 361:21]
  wire  last_q_236_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_236_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_236_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_236_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_236_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_236_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_237_clock; // @[Stab.scala 175:24]
  wire  last_merger_237_reset; // @[Stab.scala 175:24]
  wire  last_merger_237_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_237_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_237_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_237_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_237_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_237_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_237_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_237_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_237_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_237_clock; // @[Decoupled.scala 361:21]
  wire  last_q_237_reset; // @[Decoupled.scala 361:21]
  wire  last_q_237_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_237_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_237_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_237_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_237_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_237_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_238_clock; // @[Stab.scala 175:24]
  wire  last_merger_238_reset; // @[Stab.scala 175:24]
  wire  last_merger_238_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_238_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_238_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_238_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_238_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_238_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_238_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_238_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_238_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_238_clock; // @[Decoupled.scala 361:21]
  wire  last_q_238_reset; // @[Decoupled.scala 361:21]
  wire  last_q_238_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_238_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_238_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_238_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_238_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_238_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_239_clock; // @[Stab.scala 175:24]
  wire  last_merger_239_reset; // @[Stab.scala 175:24]
  wire  last_merger_239_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_239_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_239_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_239_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_239_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_239_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_239_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_239_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_239_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_239_clock; // @[Decoupled.scala 361:21]
  wire  last_q_239_reset; // @[Decoupled.scala 361:21]
  wire  last_q_239_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_239_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_239_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_239_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_239_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_239_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_240_clock; // @[Stab.scala 175:24]
  wire  last_merger_240_reset; // @[Stab.scala 175:24]
  wire  last_merger_240_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_240_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_240_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_240_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_240_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_240_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_240_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_240_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_240_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_240_clock; // @[Decoupled.scala 361:21]
  wire  last_q_240_reset; // @[Decoupled.scala 361:21]
  wire  last_q_240_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_240_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_240_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_240_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_240_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_240_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_241_clock; // @[Stab.scala 175:24]
  wire  last_merger_241_reset; // @[Stab.scala 175:24]
  wire  last_merger_241_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_241_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_241_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_241_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_241_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_241_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_241_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_241_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_241_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_241_clock; // @[Decoupled.scala 361:21]
  wire  last_q_241_reset; // @[Decoupled.scala 361:21]
  wire  last_q_241_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_241_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_241_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_241_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_241_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_241_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_242_clock; // @[Stab.scala 175:24]
  wire  last_merger_242_reset; // @[Stab.scala 175:24]
  wire  last_merger_242_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_242_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_242_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_242_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_242_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_242_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_242_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_242_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_242_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_242_clock; // @[Decoupled.scala 361:21]
  wire  last_q_242_reset; // @[Decoupled.scala 361:21]
  wire  last_q_242_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_242_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_242_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_242_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_242_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_242_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_243_clock; // @[Stab.scala 175:24]
  wire  last_merger_243_reset; // @[Stab.scala 175:24]
  wire  last_merger_243_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_243_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_243_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_243_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_243_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_243_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_243_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_243_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_243_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_243_clock; // @[Decoupled.scala 361:21]
  wire  last_q_243_reset; // @[Decoupled.scala 361:21]
  wire  last_q_243_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_243_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_243_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_243_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_243_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_243_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_244_clock; // @[Stab.scala 175:24]
  wire  last_merger_244_reset; // @[Stab.scala 175:24]
  wire  last_merger_244_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_244_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_244_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_244_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_244_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_244_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_244_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_244_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_244_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_244_clock; // @[Decoupled.scala 361:21]
  wire  last_q_244_reset; // @[Decoupled.scala 361:21]
  wire  last_q_244_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_244_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_244_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_244_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_244_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_244_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_245_clock; // @[Stab.scala 175:24]
  wire  last_merger_245_reset; // @[Stab.scala 175:24]
  wire  last_merger_245_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_245_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_245_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_245_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_245_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_245_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_245_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_245_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_245_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_245_clock; // @[Decoupled.scala 361:21]
  wire  last_q_245_reset; // @[Decoupled.scala 361:21]
  wire  last_q_245_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_245_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_245_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_245_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_245_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_245_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_246_clock; // @[Stab.scala 175:24]
  wire  last_merger_246_reset; // @[Stab.scala 175:24]
  wire  last_merger_246_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_246_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_246_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_246_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_246_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_246_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_246_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_246_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_246_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_246_clock; // @[Decoupled.scala 361:21]
  wire  last_q_246_reset; // @[Decoupled.scala 361:21]
  wire  last_q_246_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_246_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_246_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_246_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_246_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_246_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_247_clock; // @[Stab.scala 175:24]
  wire  last_merger_247_reset; // @[Stab.scala 175:24]
  wire  last_merger_247_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_247_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_247_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_247_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_247_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_247_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_247_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_247_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_247_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_247_clock; // @[Decoupled.scala 361:21]
  wire  last_q_247_reset; // @[Decoupled.scala 361:21]
  wire  last_q_247_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_247_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_247_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_247_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_247_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_247_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_248_clock; // @[Stab.scala 175:24]
  wire  last_merger_248_reset; // @[Stab.scala 175:24]
  wire  last_merger_248_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_248_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_248_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_248_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_248_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_248_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_248_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_248_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_248_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_248_clock; // @[Decoupled.scala 361:21]
  wire  last_q_248_reset; // @[Decoupled.scala 361:21]
  wire  last_q_248_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_248_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_248_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_248_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_248_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_248_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_249_clock; // @[Stab.scala 175:24]
  wire  last_merger_249_reset; // @[Stab.scala 175:24]
  wire  last_merger_249_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_249_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_249_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_249_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_249_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_249_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_249_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_249_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_249_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_249_clock; // @[Decoupled.scala 361:21]
  wire  last_q_249_reset; // @[Decoupled.scala 361:21]
  wire  last_q_249_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_249_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_249_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_249_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_249_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_249_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_250_clock; // @[Stab.scala 175:24]
  wire  last_merger_250_reset; // @[Stab.scala 175:24]
  wire  last_merger_250_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_250_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_250_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_250_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_250_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_250_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_250_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_250_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_250_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_250_clock; // @[Decoupled.scala 361:21]
  wire  last_q_250_reset; // @[Decoupled.scala 361:21]
  wire  last_q_250_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_250_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_250_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_250_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_250_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_250_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_251_clock; // @[Stab.scala 175:24]
  wire  last_merger_251_reset; // @[Stab.scala 175:24]
  wire  last_merger_251_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_251_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_251_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_251_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_251_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_251_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_251_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_251_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_251_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_251_clock; // @[Decoupled.scala 361:21]
  wire  last_q_251_reset; // @[Decoupled.scala 361:21]
  wire  last_q_251_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_251_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_251_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_251_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_251_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_251_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_252_clock; // @[Stab.scala 175:24]
  wire  last_merger_252_reset; // @[Stab.scala 175:24]
  wire  last_merger_252_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_252_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_252_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_252_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_252_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_252_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_252_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_252_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_252_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_252_clock; // @[Decoupled.scala 361:21]
  wire  last_q_252_reset; // @[Decoupled.scala 361:21]
  wire  last_q_252_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_252_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_252_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_252_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_252_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_252_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_253_clock; // @[Stab.scala 175:24]
  wire  last_merger_253_reset; // @[Stab.scala 175:24]
  wire  last_merger_253_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_253_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_253_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_253_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_253_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_253_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_253_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_253_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_253_io_result_bits; // @[Stab.scala 175:24]
  wire  last_q_253_clock; // @[Decoupled.scala 361:21]
  wire  last_q_253_reset; // @[Decoupled.scala 361:21]
  wire  last_q_253_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_253_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_253_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_q_253_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_q_253_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_q_253_io_deq_bits; // @[Decoupled.scala 361:21]
  wire  last_merger_254_clock; // @[Stab.scala 175:24]
  wire  last_merger_254_reset; // @[Stab.scala 175:24]
  wire  last_merger_254_io_stream1_ready; // @[Stab.scala 175:24]
  wire  last_merger_254_io_stream1_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_254_io_stream1_bits; // @[Stab.scala 175:24]
  wire  last_merger_254_io_stream2_ready; // @[Stab.scala 175:24]
  wire  last_merger_254_io_stream2_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_254_io_stream2_bits; // @[Stab.scala 175:24]
  wire  last_merger_254_io_result_ready; // @[Stab.scala 175:24]
  wire  last_merger_254_io_result_valid; // @[Stab.scala 175:24]
  wire [31:0] last_merger_254_io_result_bits; // @[Stab.scala 175:24]
  wire  last_clock; // @[Decoupled.scala 361:21]
  wire  last_reset; // @[Decoupled.scala 361:21]
  wire  last_io_enq_ready; // @[Decoupled.scala 361:21]
  wire  last_io_enq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_io_enq_bits; // @[Decoupled.scala 361:21]
  wire  last_io_deq_ready; // @[Decoupled.scala 361:21]
  wire  last_io_deq_valid; // @[Decoupled.scala 361:21]
  wire [31:0] last_io_deq_bits; // @[Decoupled.scala 361:21]
  StreamMerger last_merger ( // @[Stab.scala 175:24]
    .clock(last_merger_clock),
    .reset(last_merger_reset),
    .io_stream1_ready(last_merger_io_stream1_ready),
    .io_stream1_valid(last_merger_io_stream1_valid),
    .io_stream1_bits(last_merger_io_stream1_bits),
    .io_stream2_ready(last_merger_io_stream2_ready),
    .io_stream2_valid(last_merger_io_stream2_valid),
    .io_stream2_bits(last_merger_io_stream2_bits),
    .io_result_ready(last_merger_io_result_ready),
    .io_result_valid(last_merger_io_result_valid),
    .io_result_bits(last_merger_io_result_bits)
  );
  Queue last_q ( // @[Decoupled.scala 361:21]
    .clock(last_q_clock),
    .reset(last_q_reset),
    .io_enq_ready(last_q_io_enq_ready),
    .io_enq_valid(last_q_io_enq_valid),
    .io_enq_bits(last_q_io_enq_bits),
    .io_deq_ready(last_q_io_deq_ready),
    .io_deq_valid(last_q_io_deq_valid),
    .io_deq_bits(last_q_io_deq_bits)
  );
  StreamMerger_1 last_merger_1 ( // @[Stab.scala 175:24]
    .clock(last_merger_1_clock),
    .reset(last_merger_1_reset),
    .io_stream1_ready(last_merger_1_io_stream1_ready),
    .io_stream1_valid(last_merger_1_io_stream1_valid),
    .io_stream1_bits(last_merger_1_io_stream1_bits),
    .io_stream2_ready(last_merger_1_io_stream2_ready),
    .io_stream2_valid(last_merger_1_io_stream2_valid),
    .io_stream2_bits(last_merger_1_io_stream2_bits),
    .io_result_ready(last_merger_1_io_result_ready),
    .io_result_valid(last_merger_1_io_result_valid),
    .io_result_bits(last_merger_1_io_result_bits)
  );
  Queue last_q_1 ( // @[Decoupled.scala 361:21]
    .clock(last_q_1_clock),
    .reset(last_q_1_reset),
    .io_enq_ready(last_q_1_io_enq_ready),
    .io_enq_valid(last_q_1_io_enq_valid),
    .io_enq_bits(last_q_1_io_enq_bits),
    .io_deq_ready(last_q_1_io_deq_ready),
    .io_deq_valid(last_q_1_io_deq_valid),
    .io_deq_bits(last_q_1_io_deq_bits)
  );
  StreamMerger_2 last_merger_2 ( // @[Stab.scala 175:24]
    .clock(last_merger_2_clock),
    .reset(last_merger_2_reset),
    .io_stream1_ready(last_merger_2_io_stream1_ready),
    .io_stream1_valid(last_merger_2_io_stream1_valid),
    .io_stream1_bits(last_merger_2_io_stream1_bits),
    .io_stream2_ready(last_merger_2_io_stream2_ready),
    .io_stream2_valid(last_merger_2_io_stream2_valid),
    .io_stream2_bits(last_merger_2_io_stream2_bits),
    .io_result_ready(last_merger_2_io_result_ready),
    .io_result_valid(last_merger_2_io_result_valid),
    .io_result_bits(last_merger_2_io_result_bits)
  );
  Queue last_q_2 ( // @[Decoupled.scala 361:21]
    .clock(last_q_2_clock),
    .reset(last_q_2_reset),
    .io_enq_ready(last_q_2_io_enq_ready),
    .io_enq_valid(last_q_2_io_enq_valid),
    .io_enq_bits(last_q_2_io_enq_bits),
    .io_deq_ready(last_q_2_io_deq_ready),
    .io_deq_valid(last_q_2_io_deq_valid),
    .io_deq_bits(last_q_2_io_deq_bits)
  );
  StreamMerger_3 last_merger_3 ( // @[Stab.scala 175:24]
    .clock(last_merger_3_clock),
    .reset(last_merger_3_reset),
    .io_stream1_ready(last_merger_3_io_stream1_ready),
    .io_stream1_valid(last_merger_3_io_stream1_valid),
    .io_stream1_bits(last_merger_3_io_stream1_bits),
    .io_stream2_ready(last_merger_3_io_stream2_ready),
    .io_stream2_valid(last_merger_3_io_stream2_valid),
    .io_stream2_bits(last_merger_3_io_stream2_bits),
    .io_result_ready(last_merger_3_io_result_ready),
    .io_result_valid(last_merger_3_io_result_valid),
    .io_result_bits(last_merger_3_io_result_bits)
  );
  Queue last_q_3 ( // @[Decoupled.scala 361:21]
    .clock(last_q_3_clock),
    .reset(last_q_3_reset),
    .io_enq_ready(last_q_3_io_enq_ready),
    .io_enq_valid(last_q_3_io_enq_valid),
    .io_enq_bits(last_q_3_io_enq_bits),
    .io_deq_ready(last_q_3_io_deq_ready),
    .io_deq_valid(last_q_3_io_deq_valid),
    .io_deq_bits(last_q_3_io_deq_bits)
  );
  StreamMerger_4 last_merger_4 ( // @[Stab.scala 175:24]
    .clock(last_merger_4_clock),
    .reset(last_merger_4_reset),
    .io_stream1_ready(last_merger_4_io_stream1_ready),
    .io_stream1_valid(last_merger_4_io_stream1_valid),
    .io_stream1_bits(last_merger_4_io_stream1_bits),
    .io_stream2_ready(last_merger_4_io_stream2_ready),
    .io_stream2_valid(last_merger_4_io_stream2_valid),
    .io_stream2_bits(last_merger_4_io_stream2_bits),
    .io_result_ready(last_merger_4_io_result_ready),
    .io_result_valid(last_merger_4_io_result_valid),
    .io_result_bits(last_merger_4_io_result_bits)
  );
  Queue last_q_4 ( // @[Decoupled.scala 361:21]
    .clock(last_q_4_clock),
    .reset(last_q_4_reset),
    .io_enq_ready(last_q_4_io_enq_ready),
    .io_enq_valid(last_q_4_io_enq_valid),
    .io_enq_bits(last_q_4_io_enq_bits),
    .io_deq_ready(last_q_4_io_deq_ready),
    .io_deq_valid(last_q_4_io_deq_valid),
    .io_deq_bits(last_q_4_io_deq_bits)
  );
  StreamMerger_5 last_merger_5 ( // @[Stab.scala 175:24]
    .clock(last_merger_5_clock),
    .reset(last_merger_5_reset),
    .io_stream1_ready(last_merger_5_io_stream1_ready),
    .io_stream1_valid(last_merger_5_io_stream1_valid),
    .io_stream1_bits(last_merger_5_io_stream1_bits),
    .io_stream2_ready(last_merger_5_io_stream2_ready),
    .io_stream2_valid(last_merger_5_io_stream2_valid),
    .io_stream2_bits(last_merger_5_io_stream2_bits),
    .io_result_ready(last_merger_5_io_result_ready),
    .io_result_valid(last_merger_5_io_result_valid),
    .io_result_bits(last_merger_5_io_result_bits)
  );
  Queue last_q_5 ( // @[Decoupled.scala 361:21]
    .clock(last_q_5_clock),
    .reset(last_q_5_reset),
    .io_enq_ready(last_q_5_io_enq_ready),
    .io_enq_valid(last_q_5_io_enq_valid),
    .io_enq_bits(last_q_5_io_enq_bits),
    .io_deq_ready(last_q_5_io_deq_ready),
    .io_deq_valid(last_q_5_io_deq_valid),
    .io_deq_bits(last_q_5_io_deq_bits)
  );
  StreamMerger_6 last_merger_6 ( // @[Stab.scala 175:24]
    .clock(last_merger_6_clock),
    .reset(last_merger_6_reset),
    .io_stream1_ready(last_merger_6_io_stream1_ready),
    .io_stream1_valid(last_merger_6_io_stream1_valid),
    .io_stream1_bits(last_merger_6_io_stream1_bits),
    .io_stream2_ready(last_merger_6_io_stream2_ready),
    .io_stream2_valid(last_merger_6_io_stream2_valid),
    .io_stream2_bits(last_merger_6_io_stream2_bits),
    .io_result_ready(last_merger_6_io_result_ready),
    .io_result_valid(last_merger_6_io_result_valid),
    .io_result_bits(last_merger_6_io_result_bits)
  );
  Queue last_q_6 ( // @[Decoupled.scala 361:21]
    .clock(last_q_6_clock),
    .reset(last_q_6_reset),
    .io_enq_ready(last_q_6_io_enq_ready),
    .io_enq_valid(last_q_6_io_enq_valid),
    .io_enq_bits(last_q_6_io_enq_bits),
    .io_deq_ready(last_q_6_io_deq_ready),
    .io_deq_valid(last_q_6_io_deq_valid),
    .io_deq_bits(last_q_6_io_deq_bits)
  );
  StreamMerger_7 last_merger_7 ( // @[Stab.scala 175:24]
    .clock(last_merger_7_clock),
    .reset(last_merger_7_reset),
    .io_stream1_ready(last_merger_7_io_stream1_ready),
    .io_stream1_valid(last_merger_7_io_stream1_valid),
    .io_stream1_bits(last_merger_7_io_stream1_bits),
    .io_stream2_ready(last_merger_7_io_stream2_ready),
    .io_stream2_valid(last_merger_7_io_stream2_valid),
    .io_stream2_bits(last_merger_7_io_stream2_bits),
    .io_result_ready(last_merger_7_io_result_ready),
    .io_result_valid(last_merger_7_io_result_valid),
    .io_result_bits(last_merger_7_io_result_bits)
  );
  Queue last_q_7 ( // @[Decoupled.scala 361:21]
    .clock(last_q_7_clock),
    .reset(last_q_7_reset),
    .io_enq_ready(last_q_7_io_enq_ready),
    .io_enq_valid(last_q_7_io_enq_valid),
    .io_enq_bits(last_q_7_io_enq_bits),
    .io_deq_ready(last_q_7_io_deq_ready),
    .io_deq_valid(last_q_7_io_deq_valid),
    .io_deq_bits(last_q_7_io_deq_bits)
  );
  StreamMerger_8 last_merger_8 ( // @[Stab.scala 175:24]
    .clock(last_merger_8_clock),
    .reset(last_merger_8_reset),
    .io_stream1_ready(last_merger_8_io_stream1_ready),
    .io_stream1_valid(last_merger_8_io_stream1_valid),
    .io_stream1_bits(last_merger_8_io_stream1_bits),
    .io_stream2_ready(last_merger_8_io_stream2_ready),
    .io_stream2_valid(last_merger_8_io_stream2_valid),
    .io_stream2_bits(last_merger_8_io_stream2_bits),
    .io_result_ready(last_merger_8_io_result_ready),
    .io_result_valid(last_merger_8_io_result_valid),
    .io_result_bits(last_merger_8_io_result_bits)
  );
  Queue last_q_8 ( // @[Decoupled.scala 361:21]
    .clock(last_q_8_clock),
    .reset(last_q_8_reset),
    .io_enq_ready(last_q_8_io_enq_ready),
    .io_enq_valid(last_q_8_io_enq_valid),
    .io_enq_bits(last_q_8_io_enq_bits),
    .io_deq_ready(last_q_8_io_deq_ready),
    .io_deq_valid(last_q_8_io_deq_valid),
    .io_deq_bits(last_q_8_io_deq_bits)
  );
  StreamMerger_9 last_merger_9 ( // @[Stab.scala 175:24]
    .clock(last_merger_9_clock),
    .reset(last_merger_9_reset),
    .io_stream1_ready(last_merger_9_io_stream1_ready),
    .io_stream1_valid(last_merger_9_io_stream1_valid),
    .io_stream1_bits(last_merger_9_io_stream1_bits),
    .io_stream2_ready(last_merger_9_io_stream2_ready),
    .io_stream2_valid(last_merger_9_io_stream2_valid),
    .io_stream2_bits(last_merger_9_io_stream2_bits),
    .io_result_ready(last_merger_9_io_result_ready),
    .io_result_valid(last_merger_9_io_result_valid),
    .io_result_bits(last_merger_9_io_result_bits)
  );
  Queue last_q_9 ( // @[Decoupled.scala 361:21]
    .clock(last_q_9_clock),
    .reset(last_q_9_reset),
    .io_enq_ready(last_q_9_io_enq_ready),
    .io_enq_valid(last_q_9_io_enq_valid),
    .io_enq_bits(last_q_9_io_enq_bits),
    .io_deq_ready(last_q_9_io_deq_ready),
    .io_deq_valid(last_q_9_io_deq_valid),
    .io_deq_bits(last_q_9_io_deq_bits)
  );
  StreamMerger_10 last_merger_10 ( // @[Stab.scala 175:24]
    .clock(last_merger_10_clock),
    .reset(last_merger_10_reset),
    .io_stream1_ready(last_merger_10_io_stream1_ready),
    .io_stream1_valid(last_merger_10_io_stream1_valid),
    .io_stream1_bits(last_merger_10_io_stream1_bits),
    .io_stream2_ready(last_merger_10_io_stream2_ready),
    .io_stream2_valid(last_merger_10_io_stream2_valid),
    .io_stream2_bits(last_merger_10_io_stream2_bits),
    .io_result_ready(last_merger_10_io_result_ready),
    .io_result_valid(last_merger_10_io_result_valid),
    .io_result_bits(last_merger_10_io_result_bits)
  );
  Queue last_q_10 ( // @[Decoupled.scala 361:21]
    .clock(last_q_10_clock),
    .reset(last_q_10_reset),
    .io_enq_ready(last_q_10_io_enq_ready),
    .io_enq_valid(last_q_10_io_enq_valid),
    .io_enq_bits(last_q_10_io_enq_bits),
    .io_deq_ready(last_q_10_io_deq_ready),
    .io_deq_valid(last_q_10_io_deq_valid),
    .io_deq_bits(last_q_10_io_deq_bits)
  );
  StreamMerger_11 last_merger_11 ( // @[Stab.scala 175:24]
    .clock(last_merger_11_clock),
    .reset(last_merger_11_reset),
    .io_stream1_ready(last_merger_11_io_stream1_ready),
    .io_stream1_valid(last_merger_11_io_stream1_valid),
    .io_stream1_bits(last_merger_11_io_stream1_bits),
    .io_stream2_ready(last_merger_11_io_stream2_ready),
    .io_stream2_valid(last_merger_11_io_stream2_valid),
    .io_stream2_bits(last_merger_11_io_stream2_bits),
    .io_result_ready(last_merger_11_io_result_ready),
    .io_result_valid(last_merger_11_io_result_valid),
    .io_result_bits(last_merger_11_io_result_bits)
  );
  Queue last_q_11 ( // @[Decoupled.scala 361:21]
    .clock(last_q_11_clock),
    .reset(last_q_11_reset),
    .io_enq_ready(last_q_11_io_enq_ready),
    .io_enq_valid(last_q_11_io_enq_valid),
    .io_enq_bits(last_q_11_io_enq_bits),
    .io_deq_ready(last_q_11_io_deq_ready),
    .io_deq_valid(last_q_11_io_deq_valid),
    .io_deq_bits(last_q_11_io_deq_bits)
  );
  StreamMerger_12 last_merger_12 ( // @[Stab.scala 175:24]
    .clock(last_merger_12_clock),
    .reset(last_merger_12_reset),
    .io_stream1_ready(last_merger_12_io_stream1_ready),
    .io_stream1_valid(last_merger_12_io_stream1_valid),
    .io_stream1_bits(last_merger_12_io_stream1_bits),
    .io_stream2_ready(last_merger_12_io_stream2_ready),
    .io_stream2_valid(last_merger_12_io_stream2_valid),
    .io_stream2_bits(last_merger_12_io_stream2_bits),
    .io_result_ready(last_merger_12_io_result_ready),
    .io_result_valid(last_merger_12_io_result_valid),
    .io_result_bits(last_merger_12_io_result_bits)
  );
  Queue last_q_12 ( // @[Decoupled.scala 361:21]
    .clock(last_q_12_clock),
    .reset(last_q_12_reset),
    .io_enq_ready(last_q_12_io_enq_ready),
    .io_enq_valid(last_q_12_io_enq_valid),
    .io_enq_bits(last_q_12_io_enq_bits),
    .io_deq_ready(last_q_12_io_deq_ready),
    .io_deq_valid(last_q_12_io_deq_valid),
    .io_deq_bits(last_q_12_io_deq_bits)
  );
  StreamMerger_13 last_merger_13 ( // @[Stab.scala 175:24]
    .clock(last_merger_13_clock),
    .reset(last_merger_13_reset),
    .io_stream1_ready(last_merger_13_io_stream1_ready),
    .io_stream1_valid(last_merger_13_io_stream1_valid),
    .io_stream1_bits(last_merger_13_io_stream1_bits),
    .io_stream2_ready(last_merger_13_io_stream2_ready),
    .io_stream2_valid(last_merger_13_io_stream2_valid),
    .io_stream2_bits(last_merger_13_io_stream2_bits),
    .io_result_ready(last_merger_13_io_result_ready),
    .io_result_valid(last_merger_13_io_result_valid),
    .io_result_bits(last_merger_13_io_result_bits)
  );
  Queue last_q_13 ( // @[Decoupled.scala 361:21]
    .clock(last_q_13_clock),
    .reset(last_q_13_reset),
    .io_enq_ready(last_q_13_io_enq_ready),
    .io_enq_valid(last_q_13_io_enq_valid),
    .io_enq_bits(last_q_13_io_enq_bits),
    .io_deq_ready(last_q_13_io_deq_ready),
    .io_deq_valid(last_q_13_io_deq_valid),
    .io_deq_bits(last_q_13_io_deq_bits)
  );
  StreamMerger_14 last_merger_14 ( // @[Stab.scala 175:24]
    .clock(last_merger_14_clock),
    .reset(last_merger_14_reset),
    .io_stream1_ready(last_merger_14_io_stream1_ready),
    .io_stream1_valid(last_merger_14_io_stream1_valid),
    .io_stream1_bits(last_merger_14_io_stream1_bits),
    .io_stream2_ready(last_merger_14_io_stream2_ready),
    .io_stream2_valid(last_merger_14_io_stream2_valid),
    .io_stream2_bits(last_merger_14_io_stream2_bits),
    .io_result_ready(last_merger_14_io_result_ready),
    .io_result_valid(last_merger_14_io_result_valid),
    .io_result_bits(last_merger_14_io_result_bits)
  );
  Queue last_q_14 ( // @[Decoupled.scala 361:21]
    .clock(last_q_14_clock),
    .reset(last_q_14_reset),
    .io_enq_ready(last_q_14_io_enq_ready),
    .io_enq_valid(last_q_14_io_enq_valid),
    .io_enq_bits(last_q_14_io_enq_bits),
    .io_deq_ready(last_q_14_io_deq_ready),
    .io_deq_valid(last_q_14_io_deq_valid),
    .io_deq_bits(last_q_14_io_deq_bits)
  );
  StreamMerger_15 last_merger_15 ( // @[Stab.scala 175:24]
    .clock(last_merger_15_clock),
    .reset(last_merger_15_reset),
    .io_stream1_ready(last_merger_15_io_stream1_ready),
    .io_stream1_valid(last_merger_15_io_stream1_valid),
    .io_stream1_bits(last_merger_15_io_stream1_bits),
    .io_stream2_ready(last_merger_15_io_stream2_ready),
    .io_stream2_valid(last_merger_15_io_stream2_valid),
    .io_stream2_bits(last_merger_15_io_stream2_bits),
    .io_result_ready(last_merger_15_io_result_ready),
    .io_result_valid(last_merger_15_io_result_valid),
    .io_result_bits(last_merger_15_io_result_bits)
  );
  Queue last_q_15 ( // @[Decoupled.scala 361:21]
    .clock(last_q_15_clock),
    .reset(last_q_15_reset),
    .io_enq_ready(last_q_15_io_enq_ready),
    .io_enq_valid(last_q_15_io_enq_valid),
    .io_enq_bits(last_q_15_io_enq_bits),
    .io_deq_ready(last_q_15_io_deq_ready),
    .io_deq_valid(last_q_15_io_deq_valid),
    .io_deq_bits(last_q_15_io_deq_bits)
  );
  StreamMerger_16 last_merger_16 ( // @[Stab.scala 175:24]
    .clock(last_merger_16_clock),
    .reset(last_merger_16_reset),
    .io_stream1_ready(last_merger_16_io_stream1_ready),
    .io_stream1_valid(last_merger_16_io_stream1_valid),
    .io_stream1_bits(last_merger_16_io_stream1_bits),
    .io_stream2_ready(last_merger_16_io_stream2_ready),
    .io_stream2_valid(last_merger_16_io_stream2_valid),
    .io_stream2_bits(last_merger_16_io_stream2_bits),
    .io_result_ready(last_merger_16_io_result_ready),
    .io_result_valid(last_merger_16_io_result_valid),
    .io_result_bits(last_merger_16_io_result_bits)
  );
  Queue last_q_16 ( // @[Decoupled.scala 361:21]
    .clock(last_q_16_clock),
    .reset(last_q_16_reset),
    .io_enq_ready(last_q_16_io_enq_ready),
    .io_enq_valid(last_q_16_io_enq_valid),
    .io_enq_bits(last_q_16_io_enq_bits),
    .io_deq_ready(last_q_16_io_deq_ready),
    .io_deq_valid(last_q_16_io_deq_valid),
    .io_deq_bits(last_q_16_io_deq_bits)
  );
  StreamMerger_17 last_merger_17 ( // @[Stab.scala 175:24]
    .clock(last_merger_17_clock),
    .reset(last_merger_17_reset),
    .io_stream1_ready(last_merger_17_io_stream1_ready),
    .io_stream1_valid(last_merger_17_io_stream1_valid),
    .io_stream1_bits(last_merger_17_io_stream1_bits),
    .io_stream2_ready(last_merger_17_io_stream2_ready),
    .io_stream2_valid(last_merger_17_io_stream2_valid),
    .io_stream2_bits(last_merger_17_io_stream2_bits),
    .io_result_ready(last_merger_17_io_result_ready),
    .io_result_valid(last_merger_17_io_result_valid),
    .io_result_bits(last_merger_17_io_result_bits)
  );
  Queue last_q_17 ( // @[Decoupled.scala 361:21]
    .clock(last_q_17_clock),
    .reset(last_q_17_reset),
    .io_enq_ready(last_q_17_io_enq_ready),
    .io_enq_valid(last_q_17_io_enq_valid),
    .io_enq_bits(last_q_17_io_enq_bits),
    .io_deq_ready(last_q_17_io_deq_ready),
    .io_deq_valid(last_q_17_io_deq_valid),
    .io_deq_bits(last_q_17_io_deq_bits)
  );
  StreamMerger_18 last_merger_18 ( // @[Stab.scala 175:24]
    .clock(last_merger_18_clock),
    .reset(last_merger_18_reset),
    .io_stream1_ready(last_merger_18_io_stream1_ready),
    .io_stream1_valid(last_merger_18_io_stream1_valid),
    .io_stream1_bits(last_merger_18_io_stream1_bits),
    .io_stream2_ready(last_merger_18_io_stream2_ready),
    .io_stream2_valid(last_merger_18_io_stream2_valid),
    .io_stream2_bits(last_merger_18_io_stream2_bits),
    .io_result_ready(last_merger_18_io_result_ready),
    .io_result_valid(last_merger_18_io_result_valid),
    .io_result_bits(last_merger_18_io_result_bits)
  );
  Queue last_q_18 ( // @[Decoupled.scala 361:21]
    .clock(last_q_18_clock),
    .reset(last_q_18_reset),
    .io_enq_ready(last_q_18_io_enq_ready),
    .io_enq_valid(last_q_18_io_enq_valid),
    .io_enq_bits(last_q_18_io_enq_bits),
    .io_deq_ready(last_q_18_io_deq_ready),
    .io_deq_valid(last_q_18_io_deq_valid),
    .io_deq_bits(last_q_18_io_deq_bits)
  );
  StreamMerger_19 last_merger_19 ( // @[Stab.scala 175:24]
    .clock(last_merger_19_clock),
    .reset(last_merger_19_reset),
    .io_stream1_ready(last_merger_19_io_stream1_ready),
    .io_stream1_valid(last_merger_19_io_stream1_valid),
    .io_stream1_bits(last_merger_19_io_stream1_bits),
    .io_stream2_ready(last_merger_19_io_stream2_ready),
    .io_stream2_valid(last_merger_19_io_stream2_valid),
    .io_stream2_bits(last_merger_19_io_stream2_bits),
    .io_result_ready(last_merger_19_io_result_ready),
    .io_result_valid(last_merger_19_io_result_valid),
    .io_result_bits(last_merger_19_io_result_bits)
  );
  Queue last_q_19 ( // @[Decoupled.scala 361:21]
    .clock(last_q_19_clock),
    .reset(last_q_19_reset),
    .io_enq_ready(last_q_19_io_enq_ready),
    .io_enq_valid(last_q_19_io_enq_valid),
    .io_enq_bits(last_q_19_io_enq_bits),
    .io_deq_ready(last_q_19_io_deq_ready),
    .io_deq_valid(last_q_19_io_deq_valid),
    .io_deq_bits(last_q_19_io_deq_bits)
  );
  StreamMerger_20 last_merger_20 ( // @[Stab.scala 175:24]
    .clock(last_merger_20_clock),
    .reset(last_merger_20_reset),
    .io_stream1_ready(last_merger_20_io_stream1_ready),
    .io_stream1_valid(last_merger_20_io_stream1_valid),
    .io_stream1_bits(last_merger_20_io_stream1_bits),
    .io_stream2_ready(last_merger_20_io_stream2_ready),
    .io_stream2_valid(last_merger_20_io_stream2_valid),
    .io_stream2_bits(last_merger_20_io_stream2_bits),
    .io_result_ready(last_merger_20_io_result_ready),
    .io_result_valid(last_merger_20_io_result_valid),
    .io_result_bits(last_merger_20_io_result_bits)
  );
  Queue last_q_20 ( // @[Decoupled.scala 361:21]
    .clock(last_q_20_clock),
    .reset(last_q_20_reset),
    .io_enq_ready(last_q_20_io_enq_ready),
    .io_enq_valid(last_q_20_io_enq_valid),
    .io_enq_bits(last_q_20_io_enq_bits),
    .io_deq_ready(last_q_20_io_deq_ready),
    .io_deq_valid(last_q_20_io_deq_valid),
    .io_deq_bits(last_q_20_io_deq_bits)
  );
  StreamMerger_21 last_merger_21 ( // @[Stab.scala 175:24]
    .clock(last_merger_21_clock),
    .reset(last_merger_21_reset),
    .io_stream1_ready(last_merger_21_io_stream1_ready),
    .io_stream1_valid(last_merger_21_io_stream1_valid),
    .io_stream1_bits(last_merger_21_io_stream1_bits),
    .io_stream2_ready(last_merger_21_io_stream2_ready),
    .io_stream2_valid(last_merger_21_io_stream2_valid),
    .io_stream2_bits(last_merger_21_io_stream2_bits),
    .io_result_ready(last_merger_21_io_result_ready),
    .io_result_valid(last_merger_21_io_result_valid),
    .io_result_bits(last_merger_21_io_result_bits)
  );
  Queue last_q_21 ( // @[Decoupled.scala 361:21]
    .clock(last_q_21_clock),
    .reset(last_q_21_reset),
    .io_enq_ready(last_q_21_io_enq_ready),
    .io_enq_valid(last_q_21_io_enq_valid),
    .io_enq_bits(last_q_21_io_enq_bits),
    .io_deq_ready(last_q_21_io_deq_ready),
    .io_deq_valid(last_q_21_io_deq_valid),
    .io_deq_bits(last_q_21_io_deq_bits)
  );
  StreamMerger_22 last_merger_22 ( // @[Stab.scala 175:24]
    .clock(last_merger_22_clock),
    .reset(last_merger_22_reset),
    .io_stream1_ready(last_merger_22_io_stream1_ready),
    .io_stream1_valid(last_merger_22_io_stream1_valid),
    .io_stream1_bits(last_merger_22_io_stream1_bits),
    .io_stream2_ready(last_merger_22_io_stream2_ready),
    .io_stream2_valid(last_merger_22_io_stream2_valid),
    .io_stream2_bits(last_merger_22_io_stream2_bits),
    .io_result_ready(last_merger_22_io_result_ready),
    .io_result_valid(last_merger_22_io_result_valid),
    .io_result_bits(last_merger_22_io_result_bits)
  );
  Queue last_q_22 ( // @[Decoupled.scala 361:21]
    .clock(last_q_22_clock),
    .reset(last_q_22_reset),
    .io_enq_ready(last_q_22_io_enq_ready),
    .io_enq_valid(last_q_22_io_enq_valid),
    .io_enq_bits(last_q_22_io_enq_bits),
    .io_deq_ready(last_q_22_io_deq_ready),
    .io_deq_valid(last_q_22_io_deq_valid),
    .io_deq_bits(last_q_22_io_deq_bits)
  );
  StreamMerger_23 last_merger_23 ( // @[Stab.scala 175:24]
    .clock(last_merger_23_clock),
    .reset(last_merger_23_reset),
    .io_stream1_ready(last_merger_23_io_stream1_ready),
    .io_stream1_valid(last_merger_23_io_stream1_valid),
    .io_stream1_bits(last_merger_23_io_stream1_bits),
    .io_stream2_ready(last_merger_23_io_stream2_ready),
    .io_stream2_valid(last_merger_23_io_stream2_valid),
    .io_stream2_bits(last_merger_23_io_stream2_bits),
    .io_result_ready(last_merger_23_io_result_ready),
    .io_result_valid(last_merger_23_io_result_valid),
    .io_result_bits(last_merger_23_io_result_bits)
  );
  Queue last_q_23 ( // @[Decoupled.scala 361:21]
    .clock(last_q_23_clock),
    .reset(last_q_23_reset),
    .io_enq_ready(last_q_23_io_enq_ready),
    .io_enq_valid(last_q_23_io_enq_valid),
    .io_enq_bits(last_q_23_io_enq_bits),
    .io_deq_ready(last_q_23_io_deq_ready),
    .io_deq_valid(last_q_23_io_deq_valid),
    .io_deq_bits(last_q_23_io_deq_bits)
  );
  StreamMerger_24 last_merger_24 ( // @[Stab.scala 175:24]
    .clock(last_merger_24_clock),
    .reset(last_merger_24_reset),
    .io_stream1_ready(last_merger_24_io_stream1_ready),
    .io_stream1_valid(last_merger_24_io_stream1_valid),
    .io_stream1_bits(last_merger_24_io_stream1_bits),
    .io_stream2_ready(last_merger_24_io_stream2_ready),
    .io_stream2_valid(last_merger_24_io_stream2_valid),
    .io_stream2_bits(last_merger_24_io_stream2_bits),
    .io_result_ready(last_merger_24_io_result_ready),
    .io_result_valid(last_merger_24_io_result_valid),
    .io_result_bits(last_merger_24_io_result_bits)
  );
  Queue last_q_24 ( // @[Decoupled.scala 361:21]
    .clock(last_q_24_clock),
    .reset(last_q_24_reset),
    .io_enq_ready(last_q_24_io_enq_ready),
    .io_enq_valid(last_q_24_io_enq_valid),
    .io_enq_bits(last_q_24_io_enq_bits),
    .io_deq_ready(last_q_24_io_deq_ready),
    .io_deq_valid(last_q_24_io_deq_valid),
    .io_deq_bits(last_q_24_io_deq_bits)
  );
  StreamMerger_25 last_merger_25 ( // @[Stab.scala 175:24]
    .clock(last_merger_25_clock),
    .reset(last_merger_25_reset),
    .io_stream1_ready(last_merger_25_io_stream1_ready),
    .io_stream1_valid(last_merger_25_io_stream1_valid),
    .io_stream1_bits(last_merger_25_io_stream1_bits),
    .io_stream2_ready(last_merger_25_io_stream2_ready),
    .io_stream2_valid(last_merger_25_io_stream2_valid),
    .io_stream2_bits(last_merger_25_io_stream2_bits),
    .io_result_ready(last_merger_25_io_result_ready),
    .io_result_valid(last_merger_25_io_result_valid),
    .io_result_bits(last_merger_25_io_result_bits)
  );
  Queue last_q_25 ( // @[Decoupled.scala 361:21]
    .clock(last_q_25_clock),
    .reset(last_q_25_reset),
    .io_enq_ready(last_q_25_io_enq_ready),
    .io_enq_valid(last_q_25_io_enq_valid),
    .io_enq_bits(last_q_25_io_enq_bits),
    .io_deq_ready(last_q_25_io_deq_ready),
    .io_deq_valid(last_q_25_io_deq_valid),
    .io_deq_bits(last_q_25_io_deq_bits)
  );
  StreamMerger_26 last_merger_26 ( // @[Stab.scala 175:24]
    .clock(last_merger_26_clock),
    .reset(last_merger_26_reset),
    .io_stream1_ready(last_merger_26_io_stream1_ready),
    .io_stream1_valid(last_merger_26_io_stream1_valid),
    .io_stream1_bits(last_merger_26_io_stream1_bits),
    .io_stream2_ready(last_merger_26_io_stream2_ready),
    .io_stream2_valid(last_merger_26_io_stream2_valid),
    .io_stream2_bits(last_merger_26_io_stream2_bits),
    .io_result_ready(last_merger_26_io_result_ready),
    .io_result_valid(last_merger_26_io_result_valid),
    .io_result_bits(last_merger_26_io_result_bits)
  );
  Queue last_q_26 ( // @[Decoupled.scala 361:21]
    .clock(last_q_26_clock),
    .reset(last_q_26_reset),
    .io_enq_ready(last_q_26_io_enq_ready),
    .io_enq_valid(last_q_26_io_enq_valid),
    .io_enq_bits(last_q_26_io_enq_bits),
    .io_deq_ready(last_q_26_io_deq_ready),
    .io_deq_valid(last_q_26_io_deq_valid),
    .io_deq_bits(last_q_26_io_deq_bits)
  );
  StreamMerger_27 last_merger_27 ( // @[Stab.scala 175:24]
    .clock(last_merger_27_clock),
    .reset(last_merger_27_reset),
    .io_stream1_ready(last_merger_27_io_stream1_ready),
    .io_stream1_valid(last_merger_27_io_stream1_valid),
    .io_stream1_bits(last_merger_27_io_stream1_bits),
    .io_stream2_ready(last_merger_27_io_stream2_ready),
    .io_stream2_valid(last_merger_27_io_stream2_valid),
    .io_stream2_bits(last_merger_27_io_stream2_bits),
    .io_result_ready(last_merger_27_io_result_ready),
    .io_result_valid(last_merger_27_io_result_valid),
    .io_result_bits(last_merger_27_io_result_bits)
  );
  Queue last_q_27 ( // @[Decoupled.scala 361:21]
    .clock(last_q_27_clock),
    .reset(last_q_27_reset),
    .io_enq_ready(last_q_27_io_enq_ready),
    .io_enq_valid(last_q_27_io_enq_valid),
    .io_enq_bits(last_q_27_io_enq_bits),
    .io_deq_ready(last_q_27_io_deq_ready),
    .io_deq_valid(last_q_27_io_deq_valid),
    .io_deq_bits(last_q_27_io_deq_bits)
  );
  StreamMerger_28 last_merger_28 ( // @[Stab.scala 175:24]
    .clock(last_merger_28_clock),
    .reset(last_merger_28_reset),
    .io_stream1_ready(last_merger_28_io_stream1_ready),
    .io_stream1_valid(last_merger_28_io_stream1_valid),
    .io_stream1_bits(last_merger_28_io_stream1_bits),
    .io_stream2_ready(last_merger_28_io_stream2_ready),
    .io_stream2_valid(last_merger_28_io_stream2_valid),
    .io_stream2_bits(last_merger_28_io_stream2_bits),
    .io_result_ready(last_merger_28_io_result_ready),
    .io_result_valid(last_merger_28_io_result_valid),
    .io_result_bits(last_merger_28_io_result_bits)
  );
  Queue last_q_28 ( // @[Decoupled.scala 361:21]
    .clock(last_q_28_clock),
    .reset(last_q_28_reset),
    .io_enq_ready(last_q_28_io_enq_ready),
    .io_enq_valid(last_q_28_io_enq_valid),
    .io_enq_bits(last_q_28_io_enq_bits),
    .io_deq_ready(last_q_28_io_deq_ready),
    .io_deq_valid(last_q_28_io_deq_valid),
    .io_deq_bits(last_q_28_io_deq_bits)
  );
  StreamMerger_29 last_merger_29 ( // @[Stab.scala 175:24]
    .clock(last_merger_29_clock),
    .reset(last_merger_29_reset),
    .io_stream1_ready(last_merger_29_io_stream1_ready),
    .io_stream1_valid(last_merger_29_io_stream1_valid),
    .io_stream1_bits(last_merger_29_io_stream1_bits),
    .io_stream2_ready(last_merger_29_io_stream2_ready),
    .io_stream2_valid(last_merger_29_io_stream2_valid),
    .io_stream2_bits(last_merger_29_io_stream2_bits),
    .io_result_ready(last_merger_29_io_result_ready),
    .io_result_valid(last_merger_29_io_result_valid),
    .io_result_bits(last_merger_29_io_result_bits)
  );
  Queue last_q_29 ( // @[Decoupled.scala 361:21]
    .clock(last_q_29_clock),
    .reset(last_q_29_reset),
    .io_enq_ready(last_q_29_io_enq_ready),
    .io_enq_valid(last_q_29_io_enq_valid),
    .io_enq_bits(last_q_29_io_enq_bits),
    .io_deq_ready(last_q_29_io_deq_ready),
    .io_deq_valid(last_q_29_io_deq_valid),
    .io_deq_bits(last_q_29_io_deq_bits)
  );
  StreamMerger_30 last_merger_30 ( // @[Stab.scala 175:24]
    .clock(last_merger_30_clock),
    .reset(last_merger_30_reset),
    .io_stream1_ready(last_merger_30_io_stream1_ready),
    .io_stream1_valid(last_merger_30_io_stream1_valid),
    .io_stream1_bits(last_merger_30_io_stream1_bits),
    .io_stream2_ready(last_merger_30_io_stream2_ready),
    .io_stream2_valid(last_merger_30_io_stream2_valid),
    .io_stream2_bits(last_merger_30_io_stream2_bits),
    .io_result_ready(last_merger_30_io_result_ready),
    .io_result_valid(last_merger_30_io_result_valid),
    .io_result_bits(last_merger_30_io_result_bits)
  );
  Queue last_q_30 ( // @[Decoupled.scala 361:21]
    .clock(last_q_30_clock),
    .reset(last_q_30_reset),
    .io_enq_ready(last_q_30_io_enq_ready),
    .io_enq_valid(last_q_30_io_enq_valid),
    .io_enq_bits(last_q_30_io_enq_bits),
    .io_deq_ready(last_q_30_io_deq_ready),
    .io_deq_valid(last_q_30_io_deq_valid),
    .io_deq_bits(last_q_30_io_deq_bits)
  );
  StreamMerger_31 last_merger_31 ( // @[Stab.scala 175:24]
    .clock(last_merger_31_clock),
    .reset(last_merger_31_reset),
    .io_stream1_ready(last_merger_31_io_stream1_ready),
    .io_stream1_valid(last_merger_31_io_stream1_valid),
    .io_stream1_bits(last_merger_31_io_stream1_bits),
    .io_stream2_ready(last_merger_31_io_stream2_ready),
    .io_stream2_valid(last_merger_31_io_stream2_valid),
    .io_stream2_bits(last_merger_31_io_stream2_bits),
    .io_result_ready(last_merger_31_io_result_ready),
    .io_result_valid(last_merger_31_io_result_valid),
    .io_result_bits(last_merger_31_io_result_bits)
  );
  Queue last_q_31 ( // @[Decoupled.scala 361:21]
    .clock(last_q_31_clock),
    .reset(last_q_31_reset),
    .io_enq_ready(last_q_31_io_enq_ready),
    .io_enq_valid(last_q_31_io_enq_valid),
    .io_enq_bits(last_q_31_io_enq_bits),
    .io_deq_ready(last_q_31_io_deq_ready),
    .io_deq_valid(last_q_31_io_deq_valid),
    .io_deq_bits(last_q_31_io_deq_bits)
  );
  StreamMerger_32 last_merger_32 ( // @[Stab.scala 175:24]
    .clock(last_merger_32_clock),
    .reset(last_merger_32_reset),
    .io_stream1_ready(last_merger_32_io_stream1_ready),
    .io_stream1_valid(last_merger_32_io_stream1_valid),
    .io_stream1_bits(last_merger_32_io_stream1_bits),
    .io_stream2_ready(last_merger_32_io_stream2_ready),
    .io_stream2_valid(last_merger_32_io_stream2_valid),
    .io_stream2_bits(last_merger_32_io_stream2_bits),
    .io_result_ready(last_merger_32_io_result_ready),
    .io_result_valid(last_merger_32_io_result_valid),
    .io_result_bits(last_merger_32_io_result_bits)
  );
  Queue last_q_32 ( // @[Decoupled.scala 361:21]
    .clock(last_q_32_clock),
    .reset(last_q_32_reset),
    .io_enq_ready(last_q_32_io_enq_ready),
    .io_enq_valid(last_q_32_io_enq_valid),
    .io_enq_bits(last_q_32_io_enq_bits),
    .io_deq_ready(last_q_32_io_deq_ready),
    .io_deq_valid(last_q_32_io_deq_valid),
    .io_deq_bits(last_q_32_io_deq_bits)
  );
  StreamMerger_33 last_merger_33 ( // @[Stab.scala 175:24]
    .clock(last_merger_33_clock),
    .reset(last_merger_33_reset),
    .io_stream1_ready(last_merger_33_io_stream1_ready),
    .io_stream1_valid(last_merger_33_io_stream1_valid),
    .io_stream1_bits(last_merger_33_io_stream1_bits),
    .io_stream2_ready(last_merger_33_io_stream2_ready),
    .io_stream2_valid(last_merger_33_io_stream2_valid),
    .io_stream2_bits(last_merger_33_io_stream2_bits),
    .io_result_ready(last_merger_33_io_result_ready),
    .io_result_valid(last_merger_33_io_result_valid),
    .io_result_bits(last_merger_33_io_result_bits)
  );
  Queue last_q_33 ( // @[Decoupled.scala 361:21]
    .clock(last_q_33_clock),
    .reset(last_q_33_reset),
    .io_enq_ready(last_q_33_io_enq_ready),
    .io_enq_valid(last_q_33_io_enq_valid),
    .io_enq_bits(last_q_33_io_enq_bits),
    .io_deq_ready(last_q_33_io_deq_ready),
    .io_deq_valid(last_q_33_io_deq_valid),
    .io_deq_bits(last_q_33_io_deq_bits)
  );
  StreamMerger_34 last_merger_34 ( // @[Stab.scala 175:24]
    .clock(last_merger_34_clock),
    .reset(last_merger_34_reset),
    .io_stream1_ready(last_merger_34_io_stream1_ready),
    .io_stream1_valid(last_merger_34_io_stream1_valid),
    .io_stream1_bits(last_merger_34_io_stream1_bits),
    .io_stream2_ready(last_merger_34_io_stream2_ready),
    .io_stream2_valid(last_merger_34_io_stream2_valid),
    .io_stream2_bits(last_merger_34_io_stream2_bits),
    .io_result_ready(last_merger_34_io_result_ready),
    .io_result_valid(last_merger_34_io_result_valid),
    .io_result_bits(last_merger_34_io_result_bits)
  );
  Queue last_q_34 ( // @[Decoupled.scala 361:21]
    .clock(last_q_34_clock),
    .reset(last_q_34_reset),
    .io_enq_ready(last_q_34_io_enq_ready),
    .io_enq_valid(last_q_34_io_enq_valid),
    .io_enq_bits(last_q_34_io_enq_bits),
    .io_deq_ready(last_q_34_io_deq_ready),
    .io_deq_valid(last_q_34_io_deq_valid),
    .io_deq_bits(last_q_34_io_deq_bits)
  );
  StreamMerger_35 last_merger_35 ( // @[Stab.scala 175:24]
    .clock(last_merger_35_clock),
    .reset(last_merger_35_reset),
    .io_stream1_ready(last_merger_35_io_stream1_ready),
    .io_stream1_valid(last_merger_35_io_stream1_valid),
    .io_stream1_bits(last_merger_35_io_stream1_bits),
    .io_stream2_ready(last_merger_35_io_stream2_ready),
    .io_stream2_valid(last_merger_35_io_stream2_valid),
    .io_stream2_bits(last_merger_35_io_stream2_bits),
    .io_result_ready(last_merger_35_io_result_ready),
    .io_result_valid(last_merger_35_io_result_valid),
    .io_result_bits(last_merger_35_io_result_bits)
  );
  Queue last_q_35 ( // @[Decoupled.scala 361:21]
    .clock(last_q_35_clock),
    .reset(last_q_35_reset),
    .io_enq_ready(last_q_35_io_enq_ready),
    .io_enq_valid(last_q_35_io_enq_valid),
    .io_enq_bits(last_q_35_io_enq_bits),
    .io_deq_ready(last_q_35_io_deq_ready),
    .io_deq_valid(last_q_35_io_deq_valid),
    .io_deq_bits(last_q_35_io_deq_bits)
  );
  StreamMerger_36 last_merger_36 ( // @[Stab.scala 175:24]
    .clock(last_merger_36_clock),
    .reset(last_merger_36_reset),
    .io_stream1_ready(last_merger_36_io_stream1_ready),
    .io_stream1_valid(last_merger_36_io_stream1_valid),
    .io_stream1_bits(last_merger_36_io_stream1_bits),
    .io_stream2_ready(last_merger_36_io_stream2_ready),
    .io_stream2_valid(last_merger_36_io_stream2_valid),
    .io_stream2_bits(last_merger_36_io_stream2_bits),
    .io_result_ready(last_merger_36_io_result_ready),
    .io_result_valid(last_merger_36_io_result_valid),
    .io_result_bits(last_merger_36_io_result_bits)
  );
  Queue last_q_36 ( // @[Decoupled.scala 361:21]
    .clock(last_q_36_clock),
    .reset(last_q_36_reset),
    .io_enq_ready(last_q_36_io_enq_ready),
    .io_enq_valid(last_q_36_io_enq_valid),
    .io_enq_bits(last_q_36_io_enq_bits),
    .io_deq_ready(last_q_36_io_deq_ready),
    .io_deq_valid(last_q_36_io_deq_valid),
    .io_deq_bits(last_q_36_io_deq_bits)
  );
  StreamMerger_37 last_merger_37 ( // @[Stab.scala 175:24]
    .clock(last_merger_37_clock),
    .reset(last_merger_37_reset),
    .io_stream1_ready(last_merger_37_io_stream1_ready),
    .io_stream1_valid(last_merger_37_io_stream1_valid),
    .io_stream1_bits(last_merger_37_io_stream1_bits),
    .io_stream2_ready(last_merger_37_io_stream2_ready),
    .io_stream2_valid(last_merger_37_io_stream2_valid),
    .io_stream2_bits(last_merger_37_io_stream2_bits),
    .io_result_ready(last_merger_37_io_result_ready),
    .io_result_valid(last_merger_37_io_result_valid),
    .io_result_bits(last_merger_37_io_result_bits)
  );
  Queue last_q_37 ( // @[Decoupled.scala 361:21]
    .clock(last_q_37_clock),
    .reset(last_q_37_reset),
    .io_enq_ready(last_q_37_io_enq_ready),
    .io_enq_valid(last_q_37_io_enq_valid),
    .io_enq_bits(last_q_37_io_enq_bits),
    .io_deq_ready(last_q_37_io_deq_ready),
    .io_deq_valid(last_q_37_io_deq_valid),
    .io_deq_bits(last_q_37_io_deq_bits)
  );
  StreamMerger_38 last_merger_38 ( // @[Stab.scala 175:24]
    .clock(last_merger_38_clock),
    .reset(last_merger_38_reset),
    .io_stream1_ready(last_merger_38_io_stream1_ready),
    .io_stream1_valid(last_merger_38_io_stream1_valid),
    .io_stream1_bits(last_merger_38_io_stream1_bits),
    .io_stream2_ready(last_merger_38_io_stream2_ready),
    .io_stream2_valid(last_merger_38_io_stream2_valid),
    .io_stream2_bits(last_merger_38_io_stream2_bits),
    .io_result_ready(last_merger_38_io_result_ready),
    .io_result_valid(last_merger_38_io_result_valid),
    .io_result_bits(last_merger_38_io_result_bits)
  );
  Queue last_q_38 ( // @[Decoupled.scala 361:21]
    .clock(last_q_38_clock),
    .reset(last_q_38_reset),
    .io_enq_ready(last_q_38_io_enq_ready),
    .io_enq_valid(last_q_38_io_enq_valid),
    .io_enq_bits(last_q_38_io_enq_bits),
    .io_deq_ready(last_q_38_io_deq_ready),
    .io_deq_valid(last_q_38_io_deq_valid),
    .io_deq_bits(last_q_38_io_deq_bits)
  );
  StreamMerger_39 last_merger_39 ( // @[Stab.scala 175:24]
    .clock(last_merger_39_clock),
    .reset(last_merger_39_reset),
    .io_stream1_ready(last_merger_39_io_stream1_ready),
    .io_stream1_valid(last_merger_39_io_stream1_valid),
    .io_stream1_bits(last_merger_39_io_stream1_bits),
    .io_stream2_ready(last_merger_39_io_stream2_ready),
    .io_stream2_valid(last_merger_39_io_stream2_valid),
    .io_stream2_bits(last_merger_39_io_stream2_bits),
    .io_result_ready(last_merger_39_io_result_ready),
    .io_result_valid(last_merger_39_io_result_valid),
    .io_result_bits(last_merger_39_io_result_bits)
  );
  Queue last_q_39 ( // @[Decoupled.scala 361:21]
    .clock(last_q_39_clock),
    .reset(last_q_39_reset),
    .io_enq_ready(last_q_39_io_enq_ready),
    .io_enq_valid(last_q_39_io_enq_valid),
    .io_enq_bits(last_q_39_io_enq_bits),
    .io_deq_ready(last_q_39_io_deq_ready),
    .io_deq_valid(last_q_39_io_deq_valid),
    .io_deq_bits(last_q_39_io_deq_bits)
  );
  StreamMerger_40 last_merger_40 ( // @[Stab.scala 175:24]
    .clock(last_merger_40_clock),
    .reset(last_merger_40_reset),
    .io_stream1_ready(last_merger_40_io_stream1_ready),
    .io_stream1_valid(last_merger_40_io_stream1_valid),
    .io_stream1_bits(last_merger_40_io_stream1_bits),
    .io_stream2_ready(last_merger_40_io_stream2_ready),
    .io_stream2_valid(last_merger_40_io_stream2_valid),
    .io_stream2_bits(last_merger_40_io_stream2_bits),
    .io_result_ready(last_merger_40_io_result_ready),
    .io_result_valid(last_merger_40_io_result_valid),
    .io_result_bits(last_merger_40_io_result_bits)
  );
  Queue last_q_40 ( // @[Decoupled.scala 361:21]
    .clock(last_q_40_clock),
    .reset(last_q_40_reset),
    .io_enq_ready(last_q_40_io_enq_ready),
    .io_enq_valid(last_q_40_io_enq_valid),
    .io_enq_bits(last_q_40_io_enq_bits),
    .io_deq_ready(last_q_40_io_deq_ready),
    .io_deq_valid(last_q_40_io_deq_valid),
    .io_deq_bits(last_q_40_io_deq_bits)
  );
  StreamMerger_41 last_merger_41 ( // @[Stab.scala 175:24]
    .clock(last_merger_41_clock),
    .reset(last_merger_41_reset),
    .io_stream1_ready(last_merger_41_io_stream1_ready),
    .io_stream1_valid(last_merger_41_io_stream1_valid),
    .io_stream1_bits(last_merger_41_io_stream1_bits),
    .io_stream2_ready(last_merger_41_io_stream2_ready),
    .io_stream2_valid(last_merger_41_io_stream2_valid),
    .io_stream2_bits(last_merger_41_io_stream2_bits),
    .io_result_ready(last_merger_41_io_result_ready),
    .io_result_valid(last_merger_41_io_result_valid),
    .io_result_bits(last_merger_41_io_result_bits)
  );
  Queue last_q_41 ( // @[Decoupled.scala 361:21]
    .clock(last_q_41_clock),
    .reset(last_q_41_reset),
    .io_enq_ready(last_q_41_io_enq_ready),
    .io_enq_valid(last_q_41_io_enq_valid),
    .io_enq_bits(last_q_41_io_enq_bits),
    .io_deq_ready(last_q_41_io_deq_ready),
    .io_deq_valid(last_q_41_io_deq_valid),
    .io_deq_bits(last_q_41_io_deq_bits)
  );
  StreamMerger_42 last_merger_42 ( // @[Stab.scala 175:24]
    .clock(last_merger_42_clock),
    .reset(last_merger_42_reset),
    .io_stream1_ready(last_merger_42_io_stream1_ready),
    .io_stream1_valid(last_merger_42_io_stream1_valid),
    .io_stream1_bits(last_merger_42_io_stream1_bits),
    .io_stream2_ready(last_merger_42_io_stream2_ready),
    .io_stream2_valid(last_merger_42_io_stream2_valid),
    .io_stream2_bits(last_merger_42_io_stream2_bits),
    .io_result_ready(last_merger_42_io_result_ready),
    .io_result_valid(last_merger_42_io_result_valid),
    .io_result_bits(last_merger_42_io_result_bits)
  );
  Queue last_q_42 ( // @[Decoupled.scala 361:21]
    .clock(last_q_42_clock),
    .reset(last_q_42_reset),
    .io_enq_ready(last_q_42_io_enq_ready),
    .io_enq_valid(last_q_42_io_enq_valid),
    .io_enq_bits(last_q_42_io_enq_bits),
    .io_deq_ready(last_q_42_io_deq_ready),
    .io_deq_valid(last_q_42_io_deq_valid),
    .io_deq_bits(last_q_42_io_deq_bits)
  );
  StreamMerger_43 last_merger_43 ( // @[Stab.scala 175:24]
    .clock(last_merger_43_clock),
    .reset(last_merger_43_reset),
    .io_stream1_ready(last_merger_43_io_stream1_ready),
    .io_stream1_valid(last_merger_43_io_stream1_valid),
    .io_stream1_bits(last_merger_43_io_stream1_bits),
    .io_stream2_ready(last_merger_43_io_stream2_ready),
    .io_stream2_valid(last_merger_43_io_stream2_valid),
    .io_stream2_bits(last_merger_43_io_stream2_bits),
    .io_result_ready(last_merger_43_io_result_ready),
    .io_result_valid(last_merger_43_io_result_valid),
    .io_result_bits(last_merger_43_io_result_bits)
  );
  Queue last_q_43 ( // @[Decoupled.scala 361:21]
    .clock(last_q_43_clock),
    .reset(last_q_43_reset),
    .io_enq_ready(last_q_43_io_enq_ready),
    .io_enq_valid(last_q_43_io_enq_valid),
    .io_enq_bits(last_q_43_io_enq_bits),
    .io_deq_ready(last_q_43_io_deq_ready),
    .io_deq_valid(last_q_43_io_deq_valid),
    .io_deq_bits(last_q_43_io_deq_bits)
  );
  StreamMerger_44 last_merger_44 ( // @[Stab.scala 175:24]
    .clock(last_merger_44_clock),
    .reset(last_merger_44_reset),
    .io_stream1_ready(last_merger_44_io_stream1_ready),
    .io_stream1_valid(last_merger_44_io_stream1_valid),
    .io_stream1_bits(last_merger_44_io_stream1_bits),
    .io_stream2_ready(last_merger_44_io_stream2_ready),
    .io_stream2_valid(last_merger_44_io_stream2_valid),
    .io_stream2_bits(last_merger_44_io_stream2_bits),
    .io_result_ready(last_merger_44_io_result_ready),
    .io_result_valid(last_merger_44_io_result_valid),
    .io_result_bits(last_merger_44_io_result_bits)
  );
  Queue last_q_44 ( // @[Decoupled.scala 361:21]
    .clock(last_q_44_clock),
    .reset(last_q_44_reset),
    .io_enq_ready(last_q_44_io_enq_ready),
    .io_enq_valid(last_q_44_io_enq_valid),
    .io_enq_bits(last_q_44_io_enq_bits),
    .io_deq_ready(last_q_44_io_deq_ready),
    .io_deq_valid(last_q_44_io_deq_valid),
    .io_deq_bits(last_q_44_io_deq_bits)
  );
  StreamMerger_45 last_merger_45 ( // @[Stab.scala 175:24]
    .clock(last_merger_45_clock),
    .reset(last_merger_45_reset),
    .io_stream1_ready(last_merger_45_io_stream1_ready),
    .io_stream1_valid(last_merger_45_io_stream1_valid),
    .io_stream1_bits(last_merger_45_io_stream1_bits),
    .io_stream2_ready(last_merger_45_io_stream2_ready),
    .io_stream2_valid(last_merger_45_io_stream2_valid),
    .io_stream2_bits(last_merger_45_io_stream2_bits),
    .io_result_ready(last_merger_45_io_result_ready),
    .io_result_valid(last_merger_45_io_result_valid),
    .io_result_bits(last_merger_45_io_result_bits)
  );
  Queue last_q_45 ( // @[Decoupled.scala 361:21]
    .clock(last_q_45_clock),
    .reset(last_q_45_reset),
    .io_enq_ready(last_q_45_io_enq_ready),
    .io_enq_valid(last_q_45_io_enq_valid),
    .io_enq_bits(last_q_45_io_enq_bits),
    .io_deq_ready(last_q_45_io_deq_ready),
    .io_deq_valid(last_q_45_io_deq_valid),
    .io_deq_bits(last_q_45_io_deq_bits)
  );
  StreamMerger_46 last_merger_46 ( // @[Stab.scala 175:24]
    .clock(last_merger_46_clock),
    .reset(last_merger_46_reset),
    .io_stream1_ready(last_merger_46_io_stream1_ready),
    .io_stream1_valid(last_merger_46_io_stream1_valid),
    .io_stream1_bits(last_merger_46_io_stream1_bits),
    .io_stream2_ready(last_merger_46_io_stream2_ready),
    .io_stream2_valid(last_merger_46_io_stream2_valid),
    .io_stream2_bits(last_merger_46_io_stream2_bits),
    .io_result_ready(last_merger_46_io_result_ready),
    .io_result_valid(last_merger_46_io_result_valid),
    .io_result_bits(last_merger_46_io_result_bits)
  );
  Queue last_q_46 ( // @[Decoupled.scala 361:21]
    .clock(last_q_46_clock),
    .reset(last_q_46_reset),
    .io_enq_ready(last_q_46_io_enq_ready),
    .io_enq_valid(last_q_46_io_enq_valid),
    .io_enq_bits(last_q_46_io_enq_bits),
    .io_deq_ready(last_q_46_io_deq_ready),
    .io_deq_valid(last_q_46_io_deq_valid),
    .io_deq_bits(last_q_46_io_deq_bits)
  );
  StreamMerger_47 last_merger_47 ( // @[Stab.scala 175:24]
    .clock(last_merger_47_clock),
    .reset(last_merger_47_reset),
    .io_stream1_ready(last_merger_47_io_stream1_ready),
    .io_stream1_valid(last_merger_47_io_stream1_valid),
    .io_stream1_bits(last_merger_47_io_stream1_bits),
    .io_stream2_ready(last_merger_47_io_stream2_ready),
    .io_stream2_valid(last_merger_47_io_stream2_valid),
    .io_stream2_bits(last_merger_47_io_stream2_bits),
    .io_result_ready(last_merger_47_io_result_ready),
    .io_result_valid(last_merger_47_io_result_valid),
    .io_result_bits(last_merger_47_io_result_bits)
  );
  Queue last_q_47 ( // @[Decoupled.scala 361:21]
    .clock(last_q_47_clock),
    .reset(last_q_47_reset),
    .io_enq_ready(last_q_47_io_enq_ready),
    .io_enq_valid(last_q_47_io_enq_valid),
    .io_enq_bits(last_q_47_io_enq_bits),
    .io_deq_ready(last_q_47_io_deq_ready),
    .io_deq_valid(last_q_47_io_deq_valid),
    .io_deq_bits(last_q_47_io_deq_bits)
  );
  StreamMerger_48 last_merger_48 ( // @[Stab.scala 175:24]
    .clock(last_merger_48_clock),
    .reset(last_merger_48_reset),
    .io_stream1_ready(last_merger_48_io_stream1_ready),
    .io_stream1_valid(last_merger_48_io_stream1_valid),
    .io_stream1_bits(last_merger_48_io_stream1_bits),
    .io_stream2_ready(last_merger_48_io_stream2_ready),
    .io_stream2_valid(last_merger_48_io_stream2_valid),
    .io_stream2_bits(last_merger_48_io_stream2_bits),
    .io_result_ready(last_merger_48_io_result_ready),
    .io_result_valid(last_merger_48_io_result_valid),
    .io_result_bits(last_merger_48_io_result_bits)
  );
  Queue last_q_48 ( // @[Decoupled.scala 361:21]
    .clock(last_q_48_clock),
    .reset(last_q_48_reset),
    .io_enq_ready(last_q_48_io_enq_ready),
    .io_enq_valid(last_q_48_io_enq_valid),
    .io_enq_bits(last_q_48_io_enq_bits),
    .io_deq_ready(last_q_48_io_deq_ready),
    .io_deq_valid(last_q_48_io_deq_valid),
    .io_deq_bits(last_q_48_io_deq_bits)
  );
  StreamMerger_49 last_merger_49 ( // @[Stab.scala 175:24]
    .clock(last_merger_49_clock),
    .reset(last_merger_49_reset),
    .io_stream1_ready(last_merger_49_io_stream1_ready),
    .io_stream1_valid(last_merger_49_io_stream1_valid),
    .io_stream1_bits(last_merger_49_io_stream1_bits),
    .io_stream2_ready(last_merger_49_io_stream2_ready),
    .io_stream2_valid(last_merger_49_io_stream2_valid),
    .io_stream2_bits(last_merger_49_io_stream2_bits),
    .io_result_ready(last_merger_49_io_result_ready),
    .io_result_valid(last_merger_49_io_result_valid),
    .io_result_bits(last_merger_49_io_result_bits)
  );
  Queue last_q_49 ( // @[Decoupled.scala 361:21]
    .clock(last_q_49_clock),
    .reset(last_q_49_reset),
    .io_enq_ready(last_q_49_io_enq_ready),
    .io_enq_valid(last_q_49_io_enq_valid),
    .io_enq_bits(last_q_49_io_enq_bits),
    .io_deq_ready(last_q_49_io_deq_ready),
    .io_deq_valid(last_q_49_io_deq_valid),
    .io_deq_bits(last_q_49_io_deq_bits)
  );
  StreamMerger_50 last_merger_50 ( // @[Stab.scala 175:24]
    .clock(last_merger_50_clock),
    .reset(last_merger_50_reset),
    .io_stream1_ready(last_merger_50_io_stream1_ready),
    .io_stream1_valid(last_merger_50_io_stream1_valid),
    .io_stream1_bits(last_merger_50_io_stream1_bits),
    .io_stream2_ready(last_merger_50_io_stream2_ready),
    .io_stream2_valid(last_merger_50_io_stream2_valid),
    .io_stream2_bits(last_merger_50_io_stream2_bits),
    .io_result_ready(last_merger_50_io_result_ready),
    .io_result_valid(last_merger_50_io_result_valid),
    .io_result_bits(last_merger_50_io_result_bits)
  );
  Queue last_q_50 ( // @[Decoupled.scala 361:21]
    .clock(last_q_50_clock),
    .reset(last_q_50_reset),
    .io_enq_ready(last_q_50_io_enq_ready),
    .io_enq_valid(last_q_50_io_enq_valid),
    .io_enq_bits(last_q_50_io_enq_bits),
    .io_deq_ready(last_q_50_io_deq_ready),
    .io_deq_valid(last_q_50_io_deq_valid),
    .io_deq_bits(last_q_50_io_deq_bits)
  );
  StreamMerger_51 last_merger_51 ( // @[Stab.scala 175:24]
    .clock(last_merger_51_clock),
    .reset(last_merger_51_reset),
    .io_stream1_ready(last_merger_51_io_stream1_ready),
    .io_stream1_valid(last_merger_51_io_stream1_valid),
    .io_stream1_bits(last_merger_51_io_stream1_bits),
    .io_stream2_ready(last_merger_51_io_stream2_ready),
    .io_stream2_valid(last_merger_51_io_stream2_valid),
    .io_stream2_bits(last_merger_51_io_stream2_bits),
    .io_result_ready(last_merger_51_io_result_ready),
    .io_result_valid(last_merger_51_io_result_valid),
    .io_result_bits(last_merger_51_io_result_bits)
  );
  Queue last_q_51 ( // @[Decoupled.scala 361:21]
    .clock(last_q_51_clock),
    .reset(last_q_51_reset),
    .io_enq_ready(last_q_51_io_enq_ready),
    .io_enq_valid(last_q_51_io_enq_valid),
    .io_enq_bits(last_q_51_io_enq_bits),
    .io_deq_ready(last_q_51_io_deq_ready),
    .io_deq_valid(last_q_51_io_deq_valid),
    .io_deq_bits(last_q_51_io_deq_bits)
  );
  StreamMerger_52 last_merger_52 ( // @[Stab.scala 175:24]
    .clock(last_merger_52_clock),
    .reset(last_merger_52_reset),
    .io_stream1_ready(last_merger_52_io_stream1_ready),
    .io_stream1_valid(last_merger_52_io_stream1_valid),
    .io_stream1_bits(last_merger_52_io_stream1_bits),
    .io_stream2_ready(last_merger_52_io_stream2_ready),
    .io_stream2_valid(last_merger_52_io_stream2_valid),
    .io_stream2_bits(last_merger_52_io_stream2_bits),
    .io_result_ready(last_merger_52_io_result_ready),
    .io_result_valid(last_merger_52_io_result_valid),
    .io_result_bits(last_merger_52_io_result_bits)
  );
  Queue last_q_52 ( // @[Decoupled.scala 361:21]
    .clock(last_q_52_clock),
    .reset(last_q_52_reset),
    .io_enq_ready(last_q_52_io_enq_ready),
    .io_enq_valid(last_q_52_io_enq_valid),
    .io_enq_bits(last_q_52_io_enq_bits),
    .io_deq_ready(last_q_52_io_deq_ready),
    .io_deq_valid(last_q_52_io_deq_valid),
    .io_deq_bits(last_q_52_io_deq_bits)
  );
  StreamMerger_53 last_merger_53 ( // @[Stab.scala 175:24]
    .clock(last_merger_53_clock),
    .reset(last_merger_53_reset),
    .io_stream1_ready(last_merger_53_io_stream1_ready),
    .io_stream1_valid(last_merger_53_io_stream1_valid),
    .io_stream1_bits(last_merger_53_io_stream1_bits),
    .io_stream2_ready(last_merger_53_io_stream2_ready),
    .io_stream2_valid(last_merger_53_io_stream2_valid),
    .io_stream2_bits(last_merger_53_io_stream2_bits),
    .io_result_ready(last_merger_53_io_result_ready),
    .io_result_valid(last_merger_53_io_result_valid),
    .io_result_bits(last_merger_53_io_result_bits)
  );
  Queue last_q_53 ( // @[Decoupled.scala 361:21]
    .clock(last_q_53_clock),
    .reset(last_q_53_reset),
    .io_enq_ready(last_q_53_io_enq_ready),
    .io_enq_valid(last_q_53_io_enq_valid),
    .io_enq_bits(last_q_53_io_enq_bits),
    .io_deq_ready(last_q_53_io_deq_ready),
    .io_deq_valid(last_q_53_io_deq_valid),
    .io_deq_bits(last_q_53_io_deq_bits)
  );
  StreamMerger_54 last_merger_54 ( // @[Stab.scala 175:24]
    .clock(last_merger_54_clock),
    .reset(last_merger_54_reset),
    .io_stream1_ready(last_merger_54_io_stream1_ready),
    .io_stream1_valid(last_merger_54_io_stream1_valid),
    .io_stream1_bits(last_merger_54_io_stream1_bits),
    .io_stream2_ready(last_merger_54_io_stream2_ready),
    .io_stream2_valid(last_merger_54_io_stream2_valid),
    .io_stream2_bits(last_merger_54_io_stream2_bits),
    .io_result_ready(last_merger_54_io_result_ready),
    .io_result_valid(last_merger_54_io_result_valid),
    .io_result_bits(last_merger_54_io_result_bits)
  );
  Queue last_q_54 ( // @[Decoupled.scala 361:21]
    .clock(last_q_54_clock),
    .reset(last_q_54_reset),
    .io_enq_ready(last_q_54_io_enq_ready),
    .io_enq_valid(last_q_54_io_enq_valid),
    .io_enq_bits(last_q_54_io_enq_bits),
    .io_deq_ready(last_q_54_io_deq_ready),
    .io_deq_valid(last_q_54_io_deq_valid),
    .io_deq_bits(last_q_54_io_deq_bits)
  );
  StreamMerger_55 last_merger_55 ( // @[Stab.scala 175:24]
    .clock(last_merger_55_clock),
    .reset(last_merger_55_reset),
    .io_stream1_ready(last_merger_55_io_stream1_ready),
    .io_stream1_valid(last_merger_55_io_stream1_valid),
    .io_stream1_bits(last_merger_55_io_stream1_bits),
    .io_stream2_ready(last_merger_55_io_stream2_ready),
    .io_stream2_valid(last_merger_55_io_stream2_valid),
    .io_stream2_bits(last_merger_55_io_stream2_bits),
    .io_result_ready(last_merger_55_io_result_ready),
    .io_result_valid(last_merger_55_io_result_valid),
    .io_result_bits(last_merger_55_io_result_bits)
  );
  Queue last_q_55 ( // @[Decoupled.scala 361:21]
    .clock(last_q_55_clock),
    .reset(last_q_55_reset),
    .io_enq_ready(last_q_55_io_enq_ready),
    .io_enq_valid(last_q_55_io_enq_valid),
    .io_enq_bits(last_q_55_io_enq_bits),
    .io_deq_ready(last_q_55_io_deq_ready),
    .io_deq_valid(last_q_55_io_deq_valid),
    .io_deq_bits(last_q_55_io_deq_bits)
  );
  StreamMerger_56 last_merger_56 ( // @[Stab.scala 175:24]
    .clock(last_merger_56_clock),
    .reset(last_merger_56_reset),
    .io_stream1_ready(last_merger_56_io_stream1_ready),
    .io_stream1_valid(last_merger_56_io_stream1_valid),
    .io_stream1_bits(last_merger_56_io_stream1_bits),
    .io_stream2_ready(last_merger_56_io_stream2_ready),
    .io_stream2_valid(last_merger_56_io_stream2_valid),
    .io_stream2_bits(last_merger_56_io_stream2_bits),
    .io_result_ready(last_merger_56_io_result_ready),
    .io_result_valid(last_merger_56_io_result_valid),
    .io_result_bits(last_merger_56_io_result_bits)
  );
  Queue last_q_56 ( // @[Decoupled.scala 361:21]
    .clock(last_q_56_clock),
    .reset(last_q_56_reset),
    .io_enq_ready(last_q_56_io_enq_ready),
    .io_enq_valid(last_q_56_io_enq_valid),
    .io_enq_bits(last_q_56_io_enq_bits),
    .io_deq_ready(last_q_56_io_deq_ready),
    .io_deq_valid(last_q_56_io_deq_valid),
    .io_deq_bits(last_q_56_io_deq_bits)
  );
  StreamMerger_57 last_merger_57 ( // @[Stab.scala 175:24]
    .clock(last_merger_57_clock),
    .reset(last_merger_57_reset),
    .io_stream1_ready(last_merger_57_io_stream1_ready),
    .io_stream1_valid(last_merger_57_io_stream1_valid),
    .io_stream1_bits(last_merger_57_io_stream1_bits),
    .io_stream2_ready(last_merger_57_io_stream2_ready),
    .io_stream2_valid(last_merger_57_io_stream2_valid),
    .io_stream2_bits(last_merger_57_io_stream2_bits),
    .io_result_ready(last_merger_57_io_result_ready),
    .io_result_valid(last_merger_57_io_result_valid),
    .io_result_bits(last_merger_57_io_result_bits)
  );
  Queue last_q_57 ( // @[Decoupled.scala 361:21]
    .clock(last_q_57_clock),
    .reset(last_q_57_reset),
    .io_enq_ready(last_q_57_io_enq_ready),
    .io_enq_valid(last_q_57_io_enq_valid),
    .io_enq_bits(last_q_57_io_enq_bits),
    .io_deq_ready(last_q_57_io_deq_ready),
    .io_deq_valid(last_q_57_io_deq_valid),
    .io_deq_bits(last_q_57_io_deq_bits)
  );
  StreamMerger_58 last_merger_58 ( // @[Stab.scala 175:24]
    .clock(last_merger_58_clock),
    .reset(last_merger_58_reset),
    .io_stream1_ready(last_merger_58_io_stream1_ready),
    .io_stream1_valid(last_merger_58_io_stream1_valid),
    .io_stream1_bits(last_merger_58_io_stream1_bits),
    .io_stream2_ready(last_merger_58_io_stream2_ready),
    .io_stream2_valid(last_merger_58_io_stream2_valid),
    .io_stream2_bits(last_merger_58_io_stream2_bits),
    .io_result_ready(last_merger_58_io_result_ready),
    .io_result_valid(last_merger_58_io_result_valid),
    .io_result_bits(last_merger_58_io_result_bits)
  );
  Queue last_q_58 ( // @[Decoupled.scala 361:21]
    .clock(last_q_58_clock),
    .reset(last_q_58_reset),
    .io_enq_ready(last_q_58_io_enq_ready),
    .io_enq_valid(last_q_58_io_enq_valid),
    .io_enq_bits(last_q_58_io_enq_bits),
    .io_deq_ready(last_q_58_io_deq_ready),
    .io_deq_valid(last_q_58_io_deq_valid),
    .io_deq_bits(last_q_58_io_deq_bits)
  );
  StreamMerger_59 last_merger_59 ( // @[Stab.scala 175:24]
    .clock(last_merger_59_clock),
    .reset(last_merger_59_reset),
    .io_stream1_ready(last_merger_59_io_stream1_ready),
    .io_stream1_valid(last_merger_59_io_stream1_valid),
    .io_stream1_bits(last_merger_59_io_stream1_bits),
    .io_stream2_ready(last_merger_59_io_stream2_ready),
    .io_stream2_valid(last_merger_59_io_stream2_valid),
    .io_stream2_bits(last_merger_59_io_stream2_bits),
    .io_result_ready(last_merger_59_io_result_ready),
    .io_result_valid(last_merger_59_io_result_valid),
    .io_result_bits(last_merger_59_io_result_bits)
  );
  Queue last_q_59 ( // @[Decoupled.scala 361:21]
    .clock(last_q_59_clock),
    .reset(last_q_59_reset),
    .io_enq_ready(last_q_59_io_enq_ready),
    .io_enq_valid(last_q_59_io_enq_valid),
    .io_enq_bits(last_q_59_io_enq_bits),
    .io_deq_ready(last_q_59_io_deq_ready),
    .io_deq_valid(last_q_59_io_deq_valid),
    .io_deq_bits(last_q_59_io_deq_bits)
  );
  StreamMerger_60 last_merger_60 ( // @[Stab.scala 175:24]
    .clock(last_merger_60_clock),
    .reset(last_merger_60_reset),
    .io_stream1_ready(last_merger_60_io_stream1_ready),
    .io_stream1_valid(last_merger_60_io_stream1_valid),
    .io_stream1_bits(last_merger_60_io_stream1_bits),
    .io_stream2_ready(last_merger_60_io_stream2_ready),
    .io_stream2_valid(last_merger_60_io_stream2_valid),
    .io_stream2_bits(last_merger_60_io_stream2_bits),
    .io_result_ready(last_merger_60_io_result_ready),
    .io_result_valid(last_merger_60_io_result_valid),
    .io_result_bits(last_merger_60_io_result_bits)
  );
  Queue last_q_60 ( // @[Decoupled.scala 361:21]
    .clock(last_q_60_clock),
    .reset(last_q_60_reset),
    .io_enq_ready(last_q_60_io_enq_ready),
    .io_enq_valid(last_q_60_io_enq_valid),
    .io_enq_bits(last_q_60_io_enq_bits),
    .io_deq_ready(last_q_60_io_deq_ready),
    .io_deq_valid(last_q_60_io_deq_valid),
    .io_deq_bits(last_q_60_io_deq_bits)
  );
  StreamMerger_61 last_merger_61 ( // @[Stab.scala 175:24]
    .clock(last_merger_61_clock),
    .reset(last_merger_61_reset),
    .io_stream1_ready(last_merger_61_io_stream1_ready),
    .io_stream1_valid(last_merger_61_io_stream1_valid),
    .io_stream1_bits(last_merger_61_io_stream1_bits),
    .io_stream2_ready(last_merger_61_io_stream2_ready),
    .io_stream2_valid(last_merger_61_io_stream2_valid),
    .io_stream2_bits(last_merger_61_io_stream2_bits),
    .io_result_ready(last_merger_61_io_result_ready),
    .io_result_valid(last_merger_61_io_result_valid),
    .io_result_bits(last_merger_61_io_result_bits)
  );
  Queue last_q_61 ( // @[Decoupled.scala 361:21]
    .clock(last_q_61_clock),
    .reset(last_q_61_reset),
    .io_enq_ready(last_q_61_io_enq_ready),
    .io_enq_valid(last_q_61_io_enq_valid),
    .io_enq_bits(last_q_61_io_enq_bits),
    .io_deq_ready(last_q_61_io_deq_ready),
    .io_deq_valid(last_q_61_io_deq_valid),
    .io_deq_bits(last_q_61_io_deq_bits)
  );
  StreamMerger_62 last_merger_62 ( // @[Stab.scala 175:24]
    .clock(last_merger_62_clock),
    .reset(last_merger_62_reset),
    .io_stream1_ready(last_merger_62_io_stream1_ready),
    .io_stream1_valid(last_merger_62_io_stream1_valid),
    .io_stream1_bits(last_merger_62_io_stream1_bits),
    .io_stream2_ready(last_merger_62_io_stream2_ready),
    .io_stream2_valid(last_merger_62_io_stream2_valid),
    .io_stream2_bits(last_merger_62_io_stream2_bits),
    .io_result_ready(last_merger_62_io_result_ready),
    .io_result_valid(last_merger_62_io_result_valid),
    .io_result_bits(last_merger_62_io_result_bits)
  );
  Queue last_q_62 ( // @[Decoupled.scala 361:21]
    .clock(last_q_62_clock),
    .reset(last_q_62_reset),
    .io_enq_ready(last_q_62_io_enq_ready),
    .io_enq_valid(last_q_62_io_enq_valid),
    .io_enq_bits(last_q_62_io_enq_bits),
    .io_deq_ready(last_q_62_io_deq_ready),
    .io_deq_valid(last_q_62_io_deq_valid),
    .io_deq_bits(last_q_62_io_deq_bits)
  );
  StreamMerger_63 last_merger_63 ( // @[Stab.scala 175:24]
    .clock(last_merger_63_clock),
    .reset(last_merger_63_reset),
    .io_stream1_ready(last_merger_63_io_stream1_ready),
    .io_stream1_valid(last_merger_63_io_stream1_valid),
    .io_stream1_bits(last_merger_63_io_stream1_bits),
    .io_stream2_ready(last_merger_63_io_stream2_ready),
    .io_stream2_valid(last_merger_63_io_stream2_valid),
    .io_stream2_bits(last_merger_63_io_stream2_bits),
    .io_result_ready(last_merger_63_io_result_ready),
    .io_result_valid(last_merger_63_io_result_valid),
    .io_result_bits(last_merger_63_io_result_bits)
  );
  Queue last_q_63 ( // @[Decoupled.scala 361:21]
    .clock(last_q_63_clock),
    .reset(last_q_63_reset),
    .io_enq_ready(last_q_63_io_enq_ready),
    .io_enq_valid(last_q_63_io_enq_valid),
    .io_enq_bits(last_q_63_io_enq_bits),
    .io_deq_ready(last_q_63_io_deq_ready),
    .io_deq_valid(last_q_63_io_deq_valid),
    .io_deq_bits(last_q_63_io_deq_bits)
  );
  StreamMerger_64 last_merger_64 ( // @[Stab.scala 175:24]
    .clock(last_merger_64_clock),
    .reset(last_merger_64_reset),
    .io_stream1_ready(last_merger_64_io_stream1_ready),
    .io_stream1_valid(last_merger_64_io_stream1_valid),
    .io_stream1_bits(last_merger_64_io_stream1_bits),
    .io_stream2_ready(last_merger_64_io_stream2_ready),
    .io_stream2_valid(last_merger_64_io_stream2_valid),
    .io_stream2_bits(last_merger_64_io_stream2_bits),
    .io_result_ready(last_merger_64_io_result_ready),
    .io_result_valid(last_merger_64_io_result_valid),
    .io_result_bits(last_merger_64_io_result_bits)
  );
  Queue last_q_64 ( // @[Decoupled.scala 361:21]
    .clock(last_q_64_clock),
    .reset(last_q_64_reset),
    .io_enq_ready(last_q_64_io_enq_ready),
    .io_enq_valid(last_q_64_io_enq_valid),
    .io_enq_bits(last_q_64_io_enq_bits),
    .io_deq_ready(last_q_64_io_deq_ready),
    .io_deq_valid(last_q_64_io_deq_valid),
    .io_deq_bits(last_q_64_io_deq_bits)
  );
  StreamMerger_65 last_merger_65 ( // @[Stab.scala 175:24]
    .clock(last_merger_65_clock),
    .reset(last_merger_65_reset),
    .io_stream1_ready(last_merger_65_io_stream1_ready),
    .io_stream1_valid(last_merger_65_io_stream1_valid),
    .io_stream1_bits(last_merger_65_io_stream1_bits),
    .io_stream2_ready(last_merger_65_io_stream2_ready),
    .io_stream2_valid(last_merger_65_io_stream2_valid),
    .io_stream2_bits(last_merger_65_io_stream2_bits),
    .io_result_ready(last_merger_65_io_result_ready),
    .io_result_valid(last_merger_65_io_result_valid),
    .io_result_bits(last_merger_65_io_result_bits)
  );
  Queue last_q_65 ( // @[Decoupled.scala 361:21]
    .clock(last_q_65_clock),
    .reset(last_q_65_reset),
    .io_enq_ready(last_q_65_io_enq_ready),
    .io_enq_valid(last_q_65_io_enq_valid),
    .io_enq_bits(last_q_65_io_enq_bits),
    .io_deq_ready(last_q_65_io_deq_ready),
    .io_deq_valid(last_q_65_io_deq_valid),
    .io_deq_bits(last_q_65_io_deq_bits)
  );
  StreamMerger_66 last_merger_66 ( // @[Stab.scala 175:24]
    .clock(last_merger_66_clock),
    .reset(last_merger_66_reset),
    .io_stream1_ready(last_merger_66_io_stream1_ready),
    .io_stream1_valid(last_merger_66_io_stream1_valid),
    .io_stream1_bits(last_merger_66_io_stream1_bits),
    .io_stream2_ready(last_merger_66_io_stream2_ready),
    .io_stream2_valid(last_merger_66_io_stream2_valid),
    .io_stream2_bits(last_merger_66_io_stream2_bits),
    .io_result_ready(last_merger_66_io_result_ready),
    .io_result_valid(last_merger_66_io_result_valid),
    .io_result_bits(last_merger_66_io_result_bits)
  );
  Queue last_q_66 ( // @[Decoupled.scala 361:21]
    .clock(last_q_66_clock),
    .reset(last_q_66_reset),
    .io_enq_ready(last_q_66_io_enq_ready),
    .io_enq_valid(last_q_66_io_enq_valid),
    .io_enq_bits(last_q_66_io_enq_bits),
    .io_deq_ready(last_q_66_io_deq_ready),
    .io_deq_valid(last_q_66_io_deq_valid),
    .io_deq_bits(last_q_66_io_deq_bits)
  );
  StreamMerger_67 last_merger_67 ( // @[Stab.scala 175:24]
    .clock(last_merger_67_clock),
    .reset(last_merger_67_reset),
    .io_stream1_ready(last_merger_67_io_stream1_ready),
    .io_stream1_valid(last_merger_67_io_stream1_valid),
    .io_stream1_bits(last_merger_67_io_stream1_bits),
    .io_stream2_ready(last_merger_67_io_stream2_ready),
    .io_stream2_valid(last_merger_67_io_stream2_valid),
    .io_stream2_bits(last_merger_67_io_stream2_bits),
    .io_result_ready(last_merger_67_io_result_ready),
    .io_result_valid(last_merger_67_io_result_valid),
    .io_result_bits(last_merger_67_io_result_bits)
  );
  Queue last_q_67 ( // @[Decoupled.scala 361:21]
    .clock(last_q_67_clock),
    .reset(last_q_67_reset),
    .io_enq_ready(last_q_67_io_enq_ready),
    .io_enq_valid(last_q_67_io_enq_valid),
    .io_enq_bits(last_q_67_io_enq_bits),
    .io_deq_ready(last_q_67_io_deq_ready),
    .io_deq_valid(last_q_67_io_deq_valid),
    .io_deq_bits(last_q_67_io_deq_bits)
  );
  StreamMerger_68 last_merger_68 ( // @[Stab.scala 175:24]
    .clock(last_merger_68_clock),
    .reset(last_merger_68_reset),
    .io_stream1_ready(last_merger_68_io_stream1_ready),
    .io_stream1_valid(last_merger_68_io_stream1_valid),
    .io_stream1_bits(last_merger_68_io_stream1_bits),
    .io_stream2_ready(last_merger_68_io_stream2_ready),
    .io_stream2_valid(last_merger_68_io_stream2_valid),
    .io_stream2_bits(last_merger_68_io_stream2_bits),
    .io_result_ready(last_merger_68_io_result_ready),
    .io_result_valid(last_merger_68_io_result_valid),
    .io_result_bits(last_merger_68_io_result_bits)
  );
  Queue last_q_68 ( // @[Decoupled.scala 361:21]
    .clock(last_q_68_clock),
    .reset(last_q_68_reset),
    .io_enq_ready(last_q_68_io_enq_ready),
    .io_enq_valid(last_q_68_io_enq_valid),
    .io_enq_bits(last_q_68_io_enq_bits),
    .io_deq_ready(last_q_68_io_deq_ready),
    .io_deq_valid(last_q_68_io_deq_valid),
    .io_deq_bits(last_q_68_io_deq_bits)
  );
  StreamMerger_69 last_merger_69 ( // @[Stab.scala 175:24]
    .clock(last_merger_69_clock),
    .reset(last_merger_69_reset),
    .io_stream1_ready(last_merger_69_io_stream1_ready),
    .io_stream1_valid(last_merger_69_io_stream1_valid),
    .io_stream1_bits(last_merger_69_io_stream1_bits),
    .io_stream2_ready(last_merger_69_io_stream2_ready),
    .io_stream2_valid(last_merger_69_io_stream2_valid),
    .io_stream2_bits(last_merger_69_io_stream2_bits),
    .io_result_ready(last_merger_69_io_result_ready),
    .io_result_valid(last_merger_69_io_result_valid),
    .io_result_bits(last_merger_69_io_result_bits)
  );
  Queue last_q_69 ( // @[Decoupled.scala 361:21]
    .clock(last_q_69_clock),
    .reset(last_q_69_reset),
    .io_enq_ready(last_q_69_io_enq_ready),
    .io_enq_valid(last_q_69_io_enq_valid),
    .io_enq_bits(last_q_69_io_enq_bits),
    .io_deq_ready(last_q_69_io_deq_ready),
    .io_deq_valid(last_q_69_io_deq_valid),
    .io_deq_bits(last_q_69_io_deq_bits)
  );
  StreamMerger_70 last_merger_70 ( // @[Stab.scala 175:24]
    .clock(last_merger_70_clock),
    .reset(last_merger_70_reset),
    .io_stream1_ready(last_merger_70_io_stream1_ready),
    .io_stream1_valid(last_merger_70_io_stream1_valid),
    .io_stream1_bits(last_merger_70_io_stream1_bits),
    .io_stream2_ready(last_merger_70_io_stream2_ready),
    .io_stream2_valid(last_merger_70_io_stream2_valid),
    .io_stream2_bits(last_merger_70_io_stream2_bits),
    .io_result_ready(last_merger_70_io_result_ready),
    .io_result_valid(last_merger_70_io_result_valid),
    .io_result_bits(last_merger_70_io_result_bits)
  );
  Queue last_q_70 ( // @[Decoupled.scala 361:21]
    .clock(last_q_70_clock),
    .reset(last_q_70_reset),
    .io_enq_ready(last_q_70_io_enq_ready),
    .io_enq_valid(last_q_70_io_enq_valid),
    .io_enq_bits(last_q_70_io_enq_bits),
    .io_deq_ready(last_q_70_io_deq_ready),
    .io_deq_valid(last_q_70_io_deq_valid),
    .io_deq_bits(last_q_70_io_deq_bits)
  );
  StreamMerger_71 last_merger_71 ( // @[Stab.scala 175:24]
    .clock(last_merger_71_clock),
    .reset(last_merger_71_reset),
    .io_stream1_ready(last_merger_71_io_stream1_ready),
    .io_stream1_valid(last_merger_71_io_stream1_valid),
    .io_stream1_bits(last_merger_71_io_stream1_bits),
    .io_stream2_ready(last_merger_71_io_stream2_ready),
    .io_stream2_valid(last_merger_71_io_stream2_valid),
    .io_stream2_bits(last_merger_71_io_stream2_bits),
    .io_result_ready(last_merger_71_io_result_ready),
    .io_result_valid(last_merger_71_io_result_valid),
    .io_result_bits(last_merger_71_io_result_bits)
  );
  Queue last_q_71 ( // @[Decoupled.scala 361:21]
    .clock(last_q_71_clock),
    .reset(last_q_71_reset),
    .io_enq_ready(last_q_71_io_enq_ready),
    .io_enq_valid(last_q_71_io_enq_valid),
    .io_enq_bits(last_q_71_io_enq_bits),
    .io_deq_ready(last_q_71_io_deq_ready),
    .io_deq_valid(last_q_71_io_deq_valid),
    .io_deq_bits(last_q_71_io_deq_bits)
  );
  StreamMerger_72 last_merger_72 ( // @[Stab.scala 175:24]
    .clock(last_merger_72_clock),
    .reset(last_merger_72_reset),
    .io_stream1_ready(last_merger_72_io_stream1_ready),
    .io_stream1_valid(last_merger_72_io_stream1_valid),
    .io_stream1_bits(last_merger_72_io_stream1_bits),
    .io_stream2_ready(last_merger_72_io_stream2_ready),
    .io_stream2_valid(last_merger_72_io_stream2_valid),
    .io_stream2_bits(last_merger_72_io_stream2_bits),
    .io_result_ready(last_merger_72_io_result_ready),
    .io_result_valid(last_merger_72_io_result_valid),
    .io_result_bits(last_merger_72_io_result_bits)
  );
  Queue last_q_72 ( // @[Decoupled.scala 361:21]
    .clock(last_q_72_clock),
    .reset(last_q_72_reset),
    .io_enq_ready(last_q_72_io_enq_ready),
    .io_enq_valid(last_q_72_io_enq_valid),
    .io_enq_bits(last_q_72_io_enq_bits),
    .io_deq_ready(last_q_72_io_deq_ready),
    .io_deq_valid(last_q_72_io_deq_valid),
    .io_deq_bits(last_q_72_io_deq_bits)
  );
  StreamMerger_73 last_merger_73 ( // @[Stab.scala 175:24]
    .clock(last_merger_73_clock),
    .reset(last_merger_73_reset),
    .io_stream1_ready(last_merger_73_io_stream1_ready),
    .io_stream1_valid(last_merger_73_io_stream1_valid),
    .io_stream1_bits(last_merger_73_io_stream1_bits),
    .io_stream2_ready(last_merger_73_io_stream2_ready),
    .io_stream2_valid(last_merger_73_io_stream2_valid),
    .io_stream2_bits(last_merger_73_io_stream2_bits),
    .io_result_ready(last_merger_73_io_result_ready),
    .io_result_valid(last_merger_73_io_result_valid),
    .io_result_bits(last_merger_73_io_result_bits)
  );
  Queue last_q_73 ( // @[Decoupled.scala 361:21]
    .clock(last_q_73_clock),
    .reset(last_q_73_reset),
    .io_enq_ready(last_q_73_io_enq_ready),
    .io_enq_valid(last_q_73_io_enq_valid),
    .io_enq_bits(last_q_73_io_enq_bits),
    .io_deq_ready(last_q_73_io_deq_ready),
    .io_deq_valid(last_q_73_io_deq_valid),
    .io_deq_bits(last_q_73_io_deq_bits)
  );
  StreamMerger_74 last_merger_74 ( // @[Stab.scala 175:24]
    .clock(last_merger_74_clock),
    .reset(last_merger_74_reset),
    .io_stream1_ready(last_merger_74_io_stream1_ready),
    .io_stream1_valid(last_merger_74_io_stream1_valid),
    .io_stream1_bits(last_merger_74_io_stream1_bits),
    .io_stream2_ready(last_merger_74_io_stream2_ready),
    .io_stream2_valid(last_merger_74_io_stream2_valid),
    .io_stream2_bits(last_merger_74_io_stream2_bits),
    .io_result_ready(last_merger_74_io_result_ready),
    .io_result_valid(last_merger_74_io_result_valid),
    .io_result_bits(last_merger_74_io_result_bits)
  );
  Queue last_q_74 ( // @[Decoupled.scala 361:21]
    .clock(last_q_74_clock),
    .reset(last_q_74_reset),
    .io_enq_ready(last_q_74_io_enq_ready),
    .io_enq_valid(last_q_74_io_enq_valid),
    .io_enq_bits(last_q_74_io_enq_bits),
    .io_deq_ready(last_q_74_io_deq_ready),
    .io_deq_valid(last_q_74_io_deq_valid),
    .io_deq_bits(last_q_74_io_deq_bits)
  );
  StreamMerger_75 last_merger_75 ( // @[Stab.scala 175:24]
    .clock(last_merger_75_clock),
    .reset(last_merger_75_reset),
    .io_stream1_ready(last_merger_75_io_stream1_ready),
    .io_stream1_valid(last_merger_75_io_stream1_valid),
    .io_stream1_bits(last_merger_75_io_stream1_bits),
    .io_stream2_ready(last_merger_75_io_stream2_ready),
    .io_stream2_valid(last_merger_75_io_stream2_valid),
    .io_stream2_bits(last_merger_75_io_stream2_bits),
    .io_result_ready(last_merger_75_io_result_ready),
    .io_result_valid(last_merger_75_io_result_valid),
    .io_result_bits(last_merger_75_io_result_bits)
  );
  Queue last_q_75 ( // @[Decoupled.scala 361:21]
    .clock(last_q_75_clock),
    .reset(last_q_75_reset),
    .io_enq_ready(last_q_75_io_enq_ready),
    .io_enq_valid(last_q_75_io_enq_valid),
    .io_enq_bits(last_q_75_io_enq_bits),
    .io_deq_ready(last_q_75_io_deq_ready),
    .io_deq_valid(last_q_75_io_deq_valid),
    .io_deq_bits(last_q_75_io_deq_bits)
  );
  StreamMerger_76 last_merger_76 ( // @[Stab.scala 175:24]
    .clock(last_merger_76_clock),
    .reset(last_merger_76_reset),
    .io_stream1_ready(last_merger_76_io_stream1_ready),
    .io_stream1_valid(last_merger_76_io_stream1_valid),
    .io_stream1_bits(last_merger_76_io_stream1_bits),
    .io_stream2_ready(last_merger_76_io_stream2_ready),
    .io_stream2_valid(last_merger_76_io_stream2_valid),
    .io_stream2_bits(last_merger_76_io_stream2_bits),
    .io_result_ready(last_merger_76_io_result_ready),
    .io_result_valid(last_merger_76_io_result_valid),
    .io_result_bits(last_merger_76_io_result_bits)
  );
  Queue last_q_76 ( // @[Decoupled.scala 361:21]
    .clock(last_q_76_clock),
    .reset(last_q_76_reset),
    .io_enq_ready(last_q_76_io_enq_ready),
    .io_enq_valid(last_q_76_io_enq_valid),
    .io_enq_bits(last_q_76_io_enq_bits),
    .io_deq_ready(last_q_76_io_deq_ready),
    .io_deq_valid(last_q_76_io_deq_valid),
    .io_deq_bits(last_q_76_io_deq_bits)
  );
  StreamMerger_77 last_merger_77 ( // @[Stab.scala 175:24]
    .clock(last_merger_77_clock),
    .reset(last_merger_77_reset),
    .io_stream1_ready(last_merger_77_io_stream1_ready),
    .io_stream1_valid(last_merger_77_io_stream1_valid),
    .io_stream1_bits(last_merger_77_io_stream1_bits),
    .io_stream2_ready(last_merger_77_io_stream2_ready),
    .io_stream2_valid(last_merger_77_io_stream2_valid),
    .io_stream2_bits(last_merger_77_io_stream2_bits),
    .io_result_ready(last_merger_77_io_result_ready),
    .io_result_valid(last_merger_77_io_result_valid),
    .io_result_bits(last_merger_77_io_result_bits)
  );
  Queue last_q_77 ( // @[Decoupled.scala 361:21]
    .clock(last_q_77_clock),
    .reset(last_q_77_reset),
    .io_enq_ready(last_q_77_io_enq_ready),
    .io_enq_valid(last_q_77_io_enq_valid),
    .io_enq_bits(last_q_77_io_enq_bits),
    .io_deq_ready(last_q_77_io_deq_ready),
    .io_deq_valid(last_q_77_io_deq_valid),
    .io_deq_bits(last_q_77_io_deq_bits)
  );
  StreamMerger_78 last_merger_78 ( // @[Stab.scala 175:24]
    .clock(last_merger_78_clock),
    .reset(last_merger_78_reset),
    .io_stream1_ready(last_merger_78_io_stream1_ready),
    .io_stream1_valid(last_merger_78_io_stream1_valid),
    .io_stream1_bits(last_merger_78_io_stream1_bits),
    .io_stream2_ready(last_merger_78_io_stream2_ready),
    .io_stream2_valid(last_merger_78_io_stream2_valid),
    .io_stream2_bits(last_merger_78_io_stream2_bits),
    .io_result_ready(last_merger_78_io_result_ready),
    .io_result_valid(last_merger_78_io_result_valid),
    .io_result_bits(last_merger_78_io_result_bits)
  );
  Queue last_q_78 ( // @[Decoupled.scala 361:21]
    .clock(last_q_78_clock),
    .reset(last_q_78_reset),
    .io_enq_ready(last_q_78_io_enq_ready),
    .io_enq_valid(last_q_78_io_enq_valid),
    .io_enq_bits(last_q_78_io_enq_bits),
    .io_deq_ready(last_q_78_io_deq_ready),
    .io_deq_valid(last_q_78_io_deq_valid),
    .io_deq_bits(last_q_78_io_deq_bits)
  );
  StreamMerger_79 last_merger_79 ( // @[Stab.scala 175:24]
    .clock(last_merger_79_clock),
    .reset(last_merger_79_reset),
    .io_stream1_ready(last_merger_79_io_stream1_ready),
    .io_stream1_valid(last_merger_79_io_stream1_valid),
    .io_stream1_bits(last_merger_79_io_stream1_bits),
    .io_stream2_ready(last_merger_79_io_stream2_ready),
    .io_stream2_valid(last_merger_79_io_stream2_valid),
    .io_stream2_bits(last_merger_79_io_stream2_bits),
    .io_result_ready(last_merger_79_io_result_ready),
    .io_result_valid(last_merger_79_io_result_valid),
    .io_result_bits(last_merger_79_io_result_bits)
  );
  Queue last_q_79 ( // @[Decoupled.scala 361:21]
    .clock(last_q_79_clock),
    .reset(last_q_79_reset),
    .io_enq_ready(last_q_79_io_enq_ready),
    .io_enq_valid(last_q_79_io_enq_valid),
    .io_enq_bits(last_q_79_io_enq_bits),
    .io_deq_ready(last_q_79_io_deq_ready),
    .io_deq_valid(last_q_79_io_deq_valid),
    .io_deq_bits(last_q_79_io_deq_bits)
  );
  StreamMerger_80 last_merger_80 ( // @[Stab.scala 175:24]
    .clock(last_merger_80_clock),
    .reset(last_merger_80_reset),
    .io_stream1_ready(last_merger_80_io_stream1_ready),
    .io_stream1_valid(last_merger_80_io_stream1_valid),
    .io_stream1_bits(last_merger_80_io_stream1_bits),
    .io_stream2_ready(last_merger_80_io_stream2_ready),
    .io_stream2_valid(last_merger_80_io_stream2_valid),
    .io_stream2_bits(last_merger_80_io_stream2_bits),
    .io_result_ready(last_merger_80_io_result_ready),
    .io_result_valid(last_merger_80_io_result_valid),
    .io_result_bits(last_merger_80_io_result_bits)
  );
  Queue last_q_80 ( // @[Decoupled.scala 361:21]
    .clock(last_q_80_clock),
    .reset(last_q_80_reset),
    .io_enq_ready(last_q_80_io_enq_ready),
    .io_enq_valid(last_q_80_io_enq_valid),
    .io_enq_bits(last_q_80_io_enq_bits),
    .io_deq_ready(last_q_80_io_deq_ready),
    .io_deq_valid(last_q_80_io_deq_valid),
    .io_deq_bits(last_q_80_io_deq_bits)
  );
  StreamMerger_81 last_merger_81 ( // @[Stab.scala 175:24]
    .clock(last_merger_81_clock),
    .reset(last_merger_81_reset),
    .io_stream1_ready(last_merger_81_io_stream1_ready),
    .io_stream1_valid(last_merger_81_io_stream1_valid),
    .io_stream1_bits(last_merger_81_io_stream1_bits),
    .io_stream2_ready(last_merger_81_io_stream2_ready),
    .io_stream2_valid(last_merger_81_io_stream2_valid),
    .io_stream2_bits(last_merger_81_io_stream2_bits),
    .io_result_ready(last_merger_81_io_result_ready),
    .io_result_valid(last_merger_81_io_result_valid),
    .io_result_bits(last_merger_81_io_result_bits)
  );
  Queue last_q_81 ( // @[Decoupled.scala 361:21]
    .clock(last_q_81_clock),
    .reset(last_q_81_reset),
    .io_enq_ready(last_q_81_io_enq_ready),
    .io_enq_valid(last_q_81_io_enq_valid),
    .io_enq_bits(last_q_81_io_enq_bits),
    .io_deq_ready(last_q_81_io_deq_ready),
    .io_deq_valid(last_q_81_io_deq_valid),
    .io_deq_bits(last_q_81_io_deq_bits)
  );
  StreamMerger_82 last_merger_82 ( // @[Stab.scala 175:24]
    .clock(last_merger_82_clock),
    .reset(last_merger_82_reset),
    .io_stream1_ready(last_merger_82_io_stream1_ready),
    .io_stream1_valid(last_merger_82_io_stream1_valid),
    .io_stream1_bits(last_merger_82_io_stream1_bits),
    .io_stream2_ready(last_merger_82_io_stream2_ready),
    .io_stream2_valid(last_merger_82_io_stream2_valid),
    .io_stream2_bits(last_merger_82_io_stream2_bits),
    .io_result_ready(last_merger_82_io_result_ready),
    .io_result_valid(last_merger_82_io_result_valid),
    .io_result_bits(last_merger_82_io_result_bits)
  );
  Queue last_q_82 ( // @[Decoupled.scala 361:21]
    .clock(last_q_82_clock),
    .reset(last_q_82_reset),
    .io_enq_ready(last_q_82_io_enq_ready),
    .io_enq_valid(last_q_82_io_enq_valid),
    .io_enq_bits(last_q_82_io_enq_bits),
    .io_deq_ready(last_q_82_io_deq_ready),
    .io_deq_valid(last_q_82_io_deq_valid),
    .io_deq_bits(last_q_82_io_deq_bits)
  );
  StreamMerger_83 last_merger_83 ( // @[Stab.scala 175:24]
    .clock(last_merger_83_clock),
    .reset(last_merger_83_reset),
    .io_stream1_ready(last_merger_83_io_stream1_ready),
    .io_stream1_valid(last_merger_83_io_stream1_valid),
    .io_stream1_bits(last_merger_83_io_stream1_bits),
    .io_stream2_ready(last_merger_83_io_stream2_ready),
    .io_stream2_valid(last_merger_83_io_stream2_valid),
    .io_stream2_bits(last_merger_83_io_stream2_bits),
    .io_result_ready(last_merger_83_io_result_ready),
    .io_result_valid(last_merger_83_io_result_valid),
    .io_result_bits(last_merger_83_io_result_bits)
  );
  Queue last_q_83 ( // @[Decoupled.scala 361:21]
    .clock(last_q_83_clock),
    .reset(last_q_83_reset),
    .io_enq_ready(last_q_83_io_enq_ready),
    .io_enq_valid(last_q_83_io_enq_valid),
    .io_enq_bits(last_q_83_io_enq_bits),
    .io_deq_ready(last_q_83_io_deq_ready),
    .io_deq_valid(last_q_83_io_deq_valid),
    .io_deq_bits(last_q_83_io_deq_bits)
  );
  StreamMerger_84 last_merger_84 ( // @[Stab.scala 175:24]
    .clock(last_merger_84_clock),
    .reset(last_merger_84_reset),
    .io_stream1_ready(last_merger_84_io_stream1_ready),
    .io_stream1_valid(last_merger_84_io_stream1_valid),
    .io_stream1_bits(last_merger_84_io_stream1_bits),
    .io_stream2_ready(last_merger_84_io_stream2_ready),
    .io_stream2_valid(last_merger_84_io_stream2_valid),
    .io_stream2_bits(last_merger_84_io_stream2_bits),
    .io_result_ready(last_merger_84_io_result_ready),
    .io_result_valid(last_merger_84_io_result_valid),
    .io_result_bits(last_merger_84_io_result_bits)
  );
  Queue last_q_84 ( // @[Decoupled.scala 361:21]
    .clock(last_q_84_clock),
    .reset(last_q_84_reset),
    .io_enq_ready(last_q_84_io_enq_ready),
    .io_enq_valid(last_q_84_io_enq_valid),
    .io_enq_bits(last_q_84_io_enq_bits),
    .io_deq_ready(last_q_84_io_deq_ready),
    .io_deq_valid(last_q_84_io_deq_valid),
    .io_deq_bits(last_q_84_io_deq_bits)
  );
  StreamMerger_85 last_merger_85 ( // @[Stab.scala 175:24]
    .clock(last_merger_85_clock),
    .reset(last_merger_85_reset),
    .io_stream1_ready(last_merger_85_io_stream1_ready),
    .io_stream1_valid(last_merger_85_io_stream1_valid),
    .io_stream1_bits(last_merger_85_io_stream1_bits),
    .io_stream2_ready(last_merger_85_io_stream2_ready),
    .io_stream2_valid(last_merger_85_io_stream2_valid),
    .io_stream2_bits(last_merger_85_io_stream2_bits),
    .io_result_ready(last_merger_85_io_result_ready),
    .io_result_valid(last_merger_85_io_result_valid),
    .io_result_bits(last_merger_85_io_result_bits)
  );
  Queue last_q_85 ( // @[Decoupled.scala 361:21]
    .clock(last_q_85_clock),
    .reset(last_q_85_reset),
    .io_enq_ready(last_q_85_io_enq_ready),
    .io_enq_valid(last_q_85_io_enq_valid),
    .io_enq_bits(last_q_85_io_enq_bits),
    .io_deq_ready(last_q_85_io_deq_ready),
    .io_deq_valid(last_q_85_io_deq_valid),
    .io_deq_bits(last_q_85_io_deq_bits)
  );
  StreamMerger_86 last_merger_86 ( // @[Stab.scala 175:24]
    .clock(last_merger_86_clock),
    .reset(last_merger_86_reset),
    .io_stream1_ready(last_merger_86_io_stream1_ready),
    .io_stream1_valid(last_merger_86_io_stream1_valid),
    .io_stream1_bits(last_merger_86_io_stream1_bits),
    .io_stream2_ready(last_merger_86_io_stream2_ready),
    .io_stream2_valid(last_merger_86_io_stream2_valid),
    .io_stream2_bits(last_merger_86_io_stream2_bits),
    .io_result_ready(last_merger_86_io_result_ready),
    .io_result_valid(last_merger_86_io_result_valid),
    .io_result_bits(last_merger_86_io_result_bits)
  );
  Queue last_q_86 ( // @[Decoupled.scala 361:21]
    .clock(last_q_86_clock),
    .reset(last_q_86_reset),
    .io_enq_ready(last_q_86_io_enq_ready),
    .io_enq_valid(last_q_86_io_enq_valid),
    .io_enq_bits(last_q_86_io_enq_bits),
    .io_deq_ready(last_q_86_io_deq_ready),
    .io_deq_valid(last_q_86_io_deq_valid),
    .io_deq_bits(last_q_86_io_deq_bits)
  );
  StreamMerger_87 last_merger_87 ( // @[Stab.scala 175:24]
    .clock(last_merger_87_clock),
    .reset(last_merger_87_reset),
    .io_stream1_ready(last_merger_87_io_stream1_ready),
    .io_stream1_valid(last_merger_87_io_stream1_valid),
    .io_stream1_bits(last_merger_87_io_stream1_bits),
    .io_stream2_ready(last_merger_87_io_stream2_ready),
    .io_stream2_valid(last_merger_87_io_stream2_valid),
    .io_stream2_bits(last_merger_87_io_stream2_bits),
    .io_result_ready(last_merger_87_io_result_ready),
    .io_result_valid(last_merger_87_io_result_valid),
    .io_result_bits(last_merger_87_io_result_bits)
  );
  Queue last_q_87 ( // @[Decoupled.scala 361:21]
    .clock(last_q_87_clock),
    .reset(last_q_87_reset),
    .io_enq_ready(last_q_87_io_enq_ready),
    .io_enq_valid(last_q_87_io_enq_valid),
    .io_enq_bits(last_q_87_io_enq_bits),
    .io_deq_ready(last_q_87_io_deq_ready),
    .io_deq_valid(last_q_87_io_deq_valid),
    .io_deq_bits(last_q_87_io_deq_bits)
  );
  StreamMerger_88 last_merger_88 ( // @[Stab.scala 175:24]
    .clock(last_merger_88_clock),
    .reset(last_merger_88_reset),
    .io_stream1_ready(last_merger_88_io_stream1_ready),
    .io_stream1_valid(last_merger_88_io_stream1_valid),
    .io_stream1_bits(last_merger_88_io_stream1_bits),
    .io_stream2_ready(last_merger_88_io_stream2_ready),
    .io_stream2_valid(last_merger_88_io_stream2_valid),
    .io_stream2_bits(last_merger_88_io_stream2_bits),
    .io_result_ready(last_merger_88_io_result_ready),
    .io_result_valid(last_merger_88_io_result_valid),
    .io_result_bits(last_merger_88_io_result_bits)
  );
  Queue last_q_88 ( // @[Decoupled.scala 361:21]
    .clock(last_q_88_clock),
    .reset(last_q_88_reset),
    .io_enq_ready(last_q_88_io_enq_ready),
    .io_enq_valid(last_q_88_io_enq_valid),
    .io_enq_bits(last_q_88_io_enq_bits),
    .io_deq_ready(last_q_88_io_deq_ready),
    .io_deq_valid(last_q_88_io_deq_valid),
    .io_deq_bits(last_q_88_io_deq_bits)
  );
  StreamMerger_89 last_merger_89 ( // @[Stab.scala 175:24]
    .clock(last_merger_89_clock),
    .reset(last_merger_89_reset),
    .io_stream1_ready(last_merger_89_io_stream1_ready),
    .io_stream1_valid(last_merger_89_io_stream1_valid),
    .io_stream1_bits(last_merger_89_io_stream1_bits),
    .io_stream2_ready(last_merger_89_io_stream2_ready),
    .io_stream2_valid(last_merger_89_io_stream2_valid),
    .io_stream2_bits(last_merger_89_io_stream2_bits),
    .io_result_ready(last_merger_89_io_result_ready),
    .io_result_valid(last_merger_89_io_result_valid),
    .io_result_bits(last_merger_89_io_result_bits)
  );
  Queue last_q_89 ( // @[Decoupled.scala 361:21]
    .clock(last_q_89_clock),
    .reset(last_q_89_reset),
    .io_enq_ready(last_q_89_io_enq_ready),
    .io_enq_valid(last_q_89_io_enq_valid),
    .io_enq_bits(last_q_89_io_enq_bits),
    .io_deq_ready(last_q_89_io_deq_ready),
    .io_deq_valid(last_q_89_io_deq_valid),
    .io_deq_bits(last_q_89_io_deq_bits)
  );
  StreamMerger_90 last_merger_90 ( // @[Stab.scala 175:24]
    .clock(last_merger_90_clock),
    .reset(last_merger_90_reset),
    .io_stream1_ready(last_merger_90_io_stream1_ready),
    .io_stream1_valid(last_merger_90_io_stream1_valid),
    .io_stream1_bits(last_merger_90_io_stream1_bits),
    .io_stream2_ready(last_merger_90_io_stream2_ready),
    .io_stream2_valid(last_merger_90_io_stream2_valid),
    .io_stream2_bits(last_merger_90_io_stream2_bits),
    .io_result_ready(last_merger_90_io_result_ready),
    .io_result_valid(last_merger_90_io_result_valid),
    .io_result_bits(last_merger_90_io_result_bits)
  );
  Queue last_q_90 ( // @[Decoupled.scala 361:21]
    .clock(last_q_90_clock),
    .reset(last_q_90_reset),
    .io_enq_ready(last_q_90_io_enq_ready),
    .io_enq_valid(last_q_90_io_enq_valid),
    .io_enq_bits(last_q_90_io_enq_bits),
    .io_deq_ready(last_q_90_io_deq_ready),
    .io_deq_valid(last_q_90_io_deq_valid),
    .io_deq_bits(last_q_90_io_deq_bits)
  );
  StreamMerger_91 last_merger_91 ( // @[Stab.scala 175:24]
    .clock(last_merger_91_clock),
    .reset(last_merger_91_reset),
    .io_stream1_ready(last_merger_91_io_stream1_ready),
    .io_stream1_valid(last_merger_91_io_stream1_valid),
    .io_stream1_bits(last_merger_91_io_stream1_bits),
    .io_stream2_ready(last_merger_91_io_stream2_ready),
    .io_stream2_valid(last_merger_91_io_stream2_valid),
    .io_stream2_bits(last_merger_91_io_stream2_bits),
    .io_result_ready(last_merger_91_io_result_ready),
    .io_result_valid(last_merger_91_io_result_valid),
    .io_result_bits(last_merger_91_io_result_bits)
  );
  Queue last_q_91 ( // @[Decoupled.scala 361:21]
    .clock(last_q_91_clock),
    .reset(last_q_91_reset),
    .io_enq_ready(last_q_91_io_enq_ready),
    .io_enq_valid(last_q_91_io_enq_valid),
    .io_enq_bits(last_q_91_io_enq_bits),
    .io_deq_ready(last_q_91_io_deq_ready),
    .io_deq_valid(last_q_91_io_deq_valid),
    .io_deq_bits(last_q_91_io_deq_bits)
  );
  StreamMerger_92 last_merger_92 ( // @[Stab.scala 175:24]
    .clock(last_merger_92_clock),
    .reset(last_merger_92_reset),
    .io_stream1_ready(last_merger_92_io_stream1_ready),
    .io_stream1_valid(last_merger_92_io_stream1_valid),
    .io_stream1_bits(last_merger_92_io_stream1_bits),
    .io_stream2_ready(last_merger_92_io_stream2_ready),
    .io_stream2_valid(last_merger_92_io_stream2_valid),
    .io_stream2_bits(last_merger_92_io_stream2_bits),
    .io_result_ready(last_merger_92_io_result_ready),
    .io_result_valid(last_merger_92_io_result_valid),
    .io_result_bits(last_merger_92_io_result_bits)
  );
  Queue last_q_92 ( // @[Decoupled.scala 361:21]
    .clock(last_q_92_clock),
    .reset(last_q_92_reset),
    .io_enq_ready(last_q_92_io_enq_ready),
    .io_enq_valid(last_q_92_io_enq_valid),
    .io_enq_bits(last_q_92_io_enq_bits),
    .io_deq_ready(last_q_92_io_deq_ready),
    .io_deq_valid(last_q_92_io_deq_valid),
    .io_deq_bits(last_q_92_io_deq_bits)
  );
  StreamMerger_93 last_merger_93 ( // @[Stab.scala 175:24]
    .clock(last_merger_93_clock),
    .reset(last_merger_93_reset),
    .io_stream1_ready(last_merger_93_io_stream1_ready),
    .io_stream1_valid(last_merger_93_io_stream1_valid),
    .io_stream1_bits(last_merger_93_io_stream1_bits),
    .io_stream2_ready(last_merger_93_io_stream2_ready),
    .io_stream2_valid(last_merger_93_io_stream2_valid),
    .io_stream2_bits(last_merger_93_io_stream2_bits),
    .io_result_ready(last_merger_93_io_result_ready),
    .io_result_valid(last_merger_93_io_result_valid),
    .io_result_bits(last_merger_93_io_result_bits)
  );
  Queue last_q_93 ( // @[Decoupled.scala 361:21]
    .clock(last_q_93_clock),
    .reset(last_q_93_reset),
    .io_enq_ready(last_q_93_io_enq_ready),
    .io_enq_valid(last_q_93_io_enq_valid),
    .io_enq_bits(last_q_93_io_enq_bits),
    .io_deq_ready(last_q_93_io_deq_ready),
    .io_deq_valid(last_q_93_io_deq_valid),
    .io_deq_bits(last_q_93_io_deq_bits)
  );
  StreamMerger_94 last_merger_94 ( // @[Stab.scala 175:24]
    .clock(last_merger_94_clock),
    .reset(last_merger_94_reset),
    .io_stream1_ready(last_merger_94_io_stream1_ready),
    .io_stream1_valid(last_merger_94_io_stream1_valid),
    .io_stream1_bits(last_merger_94_io_stream1_bits),
    .io_stream2_ready(last_merger_94_io_stream2_ready),
    .io_stream2_valid(last_merger_94_io_stream2_valid),
    .io_stream2_bits(last_merger_94_io_stream2_bits),
    .io_result_ready(last_merger_94_io_result_ready),
    .io_result_valid(last_merger_94_io_result_valid),
    .io_result_bits(last_merger_94_io_result_bits)
  );
  Queue last_q_94 ( // @[Decoupled.scala 361:21]
    .clock(last_q_94_clock),
    .reset(last_q_94_reset),
    .io_enq_ready(last_q_94_io_enq_ready),
    .io_enq_valid(last_q_94_io_enq_valid),
    .io_enq_bits(last_q_94_io_enq_bits),
    .io_deq_ready(last_q_94_io_deq_ready),
    .io_deq_valid(last_q_94_io_deq_valid),
    .io_deq_bits(last_q_94_io_deq_bits)
  );
  StreamMerger_95 last_merger_95 ( // @[Stab.scala 175:24]
    .clock(last_merger_95_clock),
    .reset(last_merger_95_reset),
    .io_stream1_ready(last_merger_95_io_stream1_ready),
    .io_stream1_valid(last_merger_95_io_stream1_valid),
    .io_stream1_bits(last_merger_95_io_stream1_bits),
    .io_stream2_ready(last_merger_95_io_stream2_ready),
    .io_stream2_valid(last_merger_95_io_stream2_valid),
    .io_stream2_bits(last_merger_95_io_stream2_bits),
    .io_result_ready(last_merger_95_io_result_ready),
    .io_result_valid(last_merger_95_io_result_valid),
    .io_result_bits(last_merger_95_io_result_bits)
  );
  Queue last_q_95 ( // @[Decoupled.scala 361:21]
    .clock(last_q_95_clock),
    .reset(last_q_95_reset),
    .io_enq_ready(last_q_95_io_enq_ready),
    .io_enq_valid(last_q_95_io_enq_valid),
    .io_enq_bits(last_q_95_io_enq_bits),
    .io_deq_ready(last_q_95_io_deq_ready),
    .io_deq_valid(last_q_95_io_deq_valid),
    .io_deq_bits(last_q_95_io_deq_bits)
  );
  StreamMerger_96 last_merger_96 ( // @[Stab.scala 175:24]
    .clock(last_merger_96_clock),
    .reset(last_merger_96_reset),
    .io_stream1_ready(last_merger_96_io_stream1_ready),
    .io_stream1_valid(last_merger_96_io_stream1_valid),
    .io_stream1_bits(last_merger_96_io_stream1_bits),
    .io_stream2_ready(last_merger_96_io_stream2_ready),
    .io_stream2_valid(last_merger_96_io_stream2_valid),
    .io_stream2_bits(last_merger_96_io_stream2_bits),
    .io_result_ready(last_merger_96_io_result_ready),
    .io_result_valid(last_merger_96_io_result_valid),
    .io_result_bits(last_merger_96_io_result_bits)
  );
  Queue last_q_96 ( // @[Decoupled.scala 361:21]
    .clock(last_q_96_clock),
    .reset(last_q_96_reset),
    .io_enq_ready(last_q_96_io_enq_ready),
    .io_enq_valid(last_q_96_io_enq_valid),
    .io_enq_bits(last_q_96_io_enq_bits),
    .io_deq_ready(last_q_96_io_deq_ready),
    .io_deq_valid(last_q_96_io_deq_valid),
    .io_deq_bits(last_q_96_io_deq_bits)
  );
  StreamMerger_97 last_merger_97 ( // @[Stab.scala 175:24]
    .clock(last_merger_97_clock),
    .reset(last_merger_97_reset),
    .io_stream1_ready(last_merger_97_io_stream1_ready),
    .io_stream1_valid(last_merger_97_io_stream1_valid),
    .io_stream1_bits(last_merger_97_io_stream1_bits),
    .io_stream2_ready(last_merger_97_io_stream2_ready),
    .io_stream2_valid(last_merger_97_io_stream2_valid),
    .io_stream2_bits(last_merger_97_io_stream2_bits),
    .io_result_ready(last_merger_97_io_result_ready),
    .io_result_valid(last_merger_97_io_result_valid),
    .io_result_bits(last_merger_97_io_result_bits)
  );
  Queue last_q_97 ( // @[Decoupled.scala 361:21]
    .clock(last_q_97_clock),
    .reset(last_q_97_reset),
    .io_enq_ready(last_q_97_io_enq_ready),
    .io_enq_valid(last_q_97_io_enq_valid),
    .io_enq_bits(last_q_97_io_enq_bits),
    .io_deq_ready(last_q_97_io_deq_ready),
    .io_deq_valid(last_q_97_io_deq_valid),
    .io_deq_bits(last_q_97_io_deq_bits)
  );
  StreamMerger_98 last_merger_98 ( // @[Stab.scala 175:24]
    .clock(last_merger_98_clock),
    .reset(last_merger_98_reset),
    .io_stream1_ready(last_merger_98_io_stream1_ready),
    .io_stream1_valid(last_merger_98_io_stream1_valid),
    .io_stream1_bits(last_merger_98_io_stream1_bits),
    .io_stream2_ready(last_merger_98_io_stream2_ready),
    .io_stream2_valid(last_merger_98_io_stream2_valid),
    .io_stream2_bits(last_merger_98_io_stream2_bits),
    .io_result_ready(last_merger_98_io_result_ready),
    .io_result_valid(last_merger_98_io_result_valid),
    .io_result_bits(last_merger_98_io_result_bits)
  );
  Queue last_q_98 ( // @[Decoupled.scala 361:21]
    .clock(last_q_98_clock),
    .reset(last_q_98_reset),
    .io_enq_ready(last_q_98_io_enq_ready),
    .io_enq_valid(last_q_98_io_enq_valid),
    .io_enq_bits(last_q_98_io_enq_bits),
    .io_deq_ready(last_q_98_io_deq_ready),
    .io_deq_valid(last_q_98_io_deq_valid),
    .io_deq_bits(last_q_98_io_deq_bits)
  );
  StreamMerger_99 last_merger_99 ( // @[Stab.scala 175:24]
    .clock(last_merger_99_clock),
    .reset(last_merger_99_reset),
    .io_stream1_ready(last_merger_99_io_stream1_ready),
    .io_stream1_valid(last_merger_99_io_stream1_valid),
    .io_stream1_bits(last_merger_99_io_stream1_bits),
    .io_stream2_ready(last_merger_99_io_stream2_ready),
    .io_stream2_valid(last_merger_99_io_stream2_valid),
    .io_stream2_bits(last_merger_99_io_stream2_bits),
    .io_result_ready(last_merger_99_io_result_ready),
    .io_result_valid(last_merger_99_io_result_valid),
    .io_result_bits(last_merger_99_io_result_bits)
  );
  Queue last_q_99 ( // @[Decoupled.scala 361:21]
    .clock(last_q_99_clock),
    .reset(last_q_99_reset),
    .io_enq_ready(last_q_99_io_enq_ready),
    .io_enq_valid(last_q_99_io_enq_valid),
    .io_enq_bits(last_q_99_io_enq_bits),
    .io_deq_ready(last_q_99_io_deq_ready),
    .io_deq_valid(last_q_99_io_deq_valid),
    .io_deq_bits(last_q_99_io_deq_bits)
  );
  StreamMerger_100 last_merger_100 ( // @[Stab.scala 175:24]
    .clock(last_merger_100_clock),
    .reset(last_merger_100_reset),
    .io_stream1_ready(last_merger_100_io_stream1_ready),
    .io_stream1_valid(last_merger_100_io_stream1_valid),
    .io_stream1_bits(last_merger_100_io_stream1_bits),
    .io_stream2_ready(last_merger_100_io_stream2_ready),
    .io_stream2_valid(last_merger_100_io_stream2_valid),
    .io_stream2_bits(last_merger_100_io_stream2_bits),
    .io_result_ready(last_merger_100_io_result_ready),
    .io_result_valid(last_merger_100_io_result_valid),
    .io_result_bits(last_merger_100_io_result_bits)
  );
  Queue last_q_100 ( // @[Decoupled.scala 361:21]
    .clock(last_q_100_clock),
    .reset(last_q_100_reset),
    .io_enq_ready(last_q_100_io_enq_ready),
    .io_enq_valid(last_q_100_io_enq_valid),
    .io_enq_bits(last_q_100_io_enq_bits),
    .io_deq_ready(last_q_100_io_deq_ready),
    .io_deq_valid(last_q_100_io_deq_valid),
    .io_deq_bits(last_q_100_io_deq_bits)
  );
  StreamMerger_101 last_merger_101 ( // @[Stab.scala 175:24]
    .clock(last_merger_101_clock),
    .reset(last_merger_101_reset),
    .io_stream1_ready(last_merger_101_io_stream1_ready),
    .io_stream1_valid(last_merger_101_io_stream1_valid),
    .io_stream1_bits(last_merger_101_io_stream1_bits),
    .io_stream2_ready(last_merger_101_io_stream2_ready),
    .io_stream2_valid(last_merger_101_io_stream2_valid),
    .io_stream2_bits(last_merger_101_io_stream2_bits),
    .io_result_ready(last_merger_101_io_result_ready),
    .io_result_valid(last_merger_101_io_result_valid),
    .io_result_bits(last_merger_101_io_result_bits)
  );
  Queue last_q_101 ( // @[Decoupled.scala 361:21]
    .clock(last_q_101_clock),
    .reset(last_q_101_reset),
    .io_enq_ready(last_q_101_io_enq_ready),
    .io_enq_valid(last_q_101_io_enq_valid),
    .io_enq_bits(last_q_101_io_enq_bits),
    .io_deq_ready(last_q_101_io_deq_ready),
    .io_deq_valid(last_q_101_io_deq_valid),
    .io_deq_bits(last_q_101_io_deq_bits)
  );
  StreamMerger_102 last_merger_102 ( // @[Stab.scala 175:24]
    .clock(last_merger_102_clock),
    .reset(last_merger_102_reset),
    .io_stream1_ready(last_merger_102_io_stream1_ready),
    .io_stream1_valid(last_merger_102_io_stream1_valid),
    .io_stream1_bits(last_merger_102_io_stream1_bits),
    .io_stream2_ready(last_merger_102_io_stream2_ready),
    .io_stream2_valid(last_merger_102_io_stream2_valid),
    .io_stream2_bits(last_merger_102_io_stream2_bits),
    .io_result_ready(last_merger_102_io_result_ready),
    .io_result_valid(last_merger_102_io_result_valid),
    .io_result_bits(last_merger_102_io_result_bits)
  );
  Queue last_q_102 ( // @[Decoupled.scala 361:21]
    .clock(last_q_102_clock),
    .reset(last_q_102_reset),
    .io_enq_ready(last_q_102_io_enq_ready),
    .io_enq_valid(last_q_102_io_enq_valid),
    .io_enq_bits(last_q_102_io_enq_bits),
    .io_deq_ready(last_q_102_io_deq_ready),
    .io_deq_valid(last_q_102_io_deq_valid),
    .io_deq_bits(last_q_102_io_deq_bits)
  );
  StreamMerger_103 last_merger_103 ( // @[Stab.scala 175:24]
    .clock(last_merger_103_clock),
    .reset(last_merger_103_reset),
    .io_stream1_ready(last_merger_103_io_stream1_ready),
    .io_stream1_valid(last_merger_103_io_stream1_valid),
    .io_stream1_bits(last_merger_103_io_stream1_bits),
    .io_stream2_ready(last_merger_103_io_stream2_ready),
    .io_stream2_valid(last_merger_103_io_stream2_valid),
    .io_stream2_bits(last_merger_103_io_stream2_bits),
    .io_result_ready(last_merger_103_io_result_ready),
    .io_result_valid(last_merger_103_io_result_valid),
    .io_result_bits(last_merger_103_io_result_bits)
  );
  Queue last_q_103 ( // @[Decoupled.scala 361:21]
    .clock(last_q_103_clock),
    .reset(last_q_103_reset),
    .io_enq_ready(last_q_103_io_enq_ready),
    .io_enq_valid(last_q_103_io_enq_valid),
    .io_enq_bits(last_q_103_io_enq_bits),
    .io_deq_ready(last_q_103_io_deq_ready),
    .io_deq_valid(last_q_103_io_deq_valid),
    .io_deq_bits(last_q_103_io_deq_bits)
  );
  StreamMerger_104 last_merger_104 ( // @[Stab.scala 175:24]
    .clock(last_merger_104_clock),
    .reset(last_merger_104_reset),
    .io_stream1_ready(last_merger_104_io_stream1_ready),
    .io_stream1_valid(last_merger_104_io_stream1_valid),
    .io_stream1_bits(last_merger_104_io_stream1_bits),
    .io_stream2_ready(last_merger_104_io_stream2_ready),
    .io_stream2_valid(last_merger_104_io_stream2_valid),
    .io_stream2_bits(last_merger_104_io_stream2_bits),
    .io_result_ready(last_merger_104_io_result_ready),
    .io_result_valid(last_merger_104_io_result_valid),
    .io_result_bits(last_merger_104_io_result_bits)
  );
  Queue last_q_104 ( // @[Decoupled.scala 361:21]
    .clock(last_q_104_clock),
    .reset(last_q_104_reset),
    .io_enq_ready(last_q_104_io_enq_ready),
    .io_enq_valid(last_q_104_io_enq_valid),
    .io_enq_bits(last_q_104_io_enq_bits),
    .io_deq_ready(last_q_104_io_deq_ready),
    .io_deq_valid(last_q_104_io_deq_valid),
    .io_deq_bits(last_q_104_io_deq_bits)
  );
  StreamMerger_105 last_merger_105 ( // @[Stab.scala 175:24]
    .clock(last_merger_105_clock),
    .reset(last_merger_105_reset),
    .io_stream1_ready(last_merger_105_io_stream1_ready),
    .io_stream1_valid(last_merger_105_io_stream1_valid),
    .io_stream1_bits(last_merger_105_io_stream1_bits),
    .io_stream2_ready(last_merger_105_io_stream2_ready),
    .io_stream2_valid(last_merger_105_io_stream2_valid),
    .io_stream2_bits(last_merger_105_io_stream2_bits),
    .io_result_ready(last_merger_105_io_result_ready),
    .io_result_valid(last_merger_105_io_result_valid),
    .io_result_bits(last_merger_105_io_result_bits)
  );
  Queue last_q_105 ( // @[Decoupled.scala 361:21]
    .clock(last_q_105_clock),
    .reset(last_q_105_reset),
    .io_enq_ready(last_q_105_io_enq_ready),
    .io_enq_valid(last_q_105_io_enq_valid),
    .io_enq_bits(last_q_105_io_enq_bits),
    .io_deq_ready(last_q_105_io_deq_ready),
    .io_deq_valid(last_q_105_io_deq_valid),
    .io_deq_bits(last_q_105_io_deq_bits)
  );
  StreamMerger_106 last_merger_106 ( // @[Stab.scala 175:24]
    .clock(last_merger_106_clock),
    .reset(last_merger_106_reset),
    .io_stream1_ready(last_merger_106_io_stream1_ready),
    .io_stream1_valid(last_merger_106_io_stream1_valid),
    .io_stream1_bits(last_merger_106_io_stream1_bits),
    .io_stream2_ready(last_merger_106_io_stream2_ready),
    .io_stream2_valid(last_merger_106_io_stream2_valid),
    .io_stream2_bits(last_merger_106_io_stream2_bits),
    .io_result_ready(last_merger_106_io_result_ready),
    .io_result_valid(last_merger_106_io_result_valid),
    .io_result_bits(last_merger_106_io_result_bits)
  );
  Queue last_q_106 ( // @[Decoupled.scala 361:21]
    .clock(last_q_106_clock),
    .reset(last_q_106_reset),
    .io_enq_ready(last_q_106_io_enq_ready),
    .io_enq_valid(last_q_106_io_enq_valid),
    .io_enq_bits(last_q_106_io_enq_bits),
    .io_deq_ready(last_q_106_io_deq_ready),
    .io_deq_valid(last_q_106_io_deq_valid),
    .io_deq_bits(last_q_106_io_deq_bits)
  );
  StreamMerger_107 last_merger_107 ( // @[Stab.scala 175:24]
    .clock(last_merger_107_clock),
    .reset(last_merger_107_reset),
    .io_stream1_ready(last_merger_107_io_stream1_ready),
    .io_stream1_valid(last_merger_107_io_stream1_valid),
    .io_stream1_bits(last_merger_107_io_stream1_bits),
    .io_stream2_ready(last_merger_107_io_stream2_ready),
    .io_stream2_valid(last_merger_107_io_stream2_valid),
    .io_stream2_bits(last_merger_107_io_stream2_bits),
    .io_result_ready(last_merger_107_io_result_ready),
    .io_result_valid(last_merger_107_io_result_valid),
    .io_result_bits(last_merger_107_io_result_bits)
  );
  Queue last_q_107 ( // @[Decoupled.scala 361:21]
    .clock(last_q_107_clock),
    .reset(last_q_107_reset),
    .io_enq_ready(last_q_107_io_enq_ready),
    .io_enq_valid(last_q_107_io_enq_valid),
    .io_enq_bits(last_q_107_io_enq_bits),
    .io_deq_ready(last_q_107_io_deq_ready),
    .io_deq_valid(last_q_107_io_deq_valid),
    .io_deq_bits(last_q_107_io_deq_bits)
  );
  StreamMerger_108 last_merger_108 ( // @[Stab.scala 175:24]
    .clock(last_merger_108_clock),
    .reset(last_merger_108_reset),
    .io_stream1_ready(last_merger_108_io_stream1_ready),
    .io_stream1_valid(last_merger_108_io_stream1_valid),
    .io_stream1_bits(last_merger_108_io_stream1_bits),
    .io_stream2_ready(last_merger_108_io_stream2_ready),
    .io_stream2_valid(last_merger_108_io_stream2_valid),
    .io_stream2_bits(last_merger_108_io_stream2_bits),
    .io_result_ready(last_merger_108_io_result_ready),
    .io_result_valid(last_merger_108_io_result_valid),
    .io_result_bits(last_merger_108_io_result_bits)
  );
  Queue last_q_108 ( // @[Decoupled.scala 361:21]
    .clock(last_q_108_clock),
    .reset(last_q_108_reset),
    .io_enq_ready(last_q_108_io_enq_ready),
    .io_enq_valid(last_q_108_io_enq_valid),
    .io_enq_bits(last_q_108_io_enq_bits),
    .io_deq_ready(last_q_108_io_deq_ready),
    .io_deq_valid(last_q_108_io_deq_valid),
    .io_deq_bits(last_q_108_io_deq_bits)
  );
  StreamMerger_109 last_merger_109 ( // @[Stab.scala 175:24]
    .clock(last_merger_109_clock),
    .reset(last_merger_109_reset),
    .io_stream1_ready(last_merger_109_io_stream1_ready),
    .io_stream1_valid(last_merger_109_io_stream1_valid),
    .io_stream1_bits(last_merger_109_io_stream1_bits),
    .io_stream2_ready(last_merger_109_io_stream2_ready),
    .io_stream2_valid(last_merger_109_io_stream2_valid),
    .io_stream2_bits(last_merger_109_io_stream2_bits),
    .io_result_ready(last_merger_109_io_result_ready),
    .io_result_valid(last_merger_109_io_result_valid),
    .io_result_bits(last_merger_109_io_result_bits)
  );
  Queue last_q_109 ( // @[Decoupled.scala 361:21]
    .clock(last_q_109_clock),
    .reset(last_q_109_reset),
    .io_enq_ready(last_q_109_io_enq_ready),
    .io_enq_valid(last_q_109_io_enq_valid),
    .io_enq_bits(last_q_109_io_enq_bits),
    .io_deq_ready(last_q_109_io_deq_ready),
    .io_deq_valid(last_q_109_io_deq_valid),
    .io_deq_bits(last_q_109_io_deq_bits)
  );
  StreamMerger_110 last_merger_110 ( // @[Stab.scala 175:24]
    .clock(last_merger_110_clock),
    .reset(last_merger_110_reset),
    .io_stream1_ready(last_merger_110_io_stream1_ready),
    .io_stream1_valid(last_merger_110_io_stream1_valid),
    .io_stream1_bits(last_merger_110_io_stream1_bits),
    .io_stream2_ready(last_merger_110_io_stream2_ready),
    .io_stream2_valid(last_merger_110_io_stream2_valid),
    .io_stream2_bits(last_merger_110_io_stream2_bits),
    .io_result_ready(last_merger_110_io_result_ready),
    .io_result_valid(last_merger_110_io_result_valid),
    .io_result_bits(last_merger_110_io_result_bits)
  );
  Queue last_q_110 ( // @[Decoupled.scala 361:21]
    .clock(last_q_110_clock),
    .reset(last_q_110_reset),
    .io_enq_ready(last_q_110_io_enq_ready),
    .io_enq_valid(last_q_110_io_enq_valid),
    .io_enq_bits(last_q_110_io_enq_bits),
    .io_deq_ready(last_q_110_io_deq_ready),
    .io_deq_valid(last_q_110_io_deq_valid),
    .io_deq_bits(last_q_110_io_deq_bits)
  );
  StreamMerger_111 last_merger_111 ( // @[Stab.scala 175:24]
    .clock(last_merger_111_clock),
    .reset(last_merger_111_reset),
    .io_stream1_ready(last_merger_111_io_stream1_ready),
    .io_stream1_valid(last_merger_111_io_stream1_valid),
    .io_stream1_bits(last_merger_111_io_stream1_bits),
    .io_stream2_ready(last_merger_111_io_stream2_ready),
    .io_stream2_valid(last_merger_111_io_stream2_valid),
    .io_stream2_bits(last_merger_111_io_stream2_bits),
    .io_result_ready(last_merger_111_io_result_ready),
    .io_result_valid(last_merger_111_io_result_valid),
    .io_result_bits(last_merger_111_io_result_bits)
  );
  Queue last_q_111 ( // @[Decoupled.scala 361:21]
    .clock(last_q_111_clock),
    .reset(last_q_111_reset),
    .io_enq_ready(last_q_111_io_enq_ready),
    .io_enq_valid(last_q_111_io_enq_valid),
    .io_enq_bits(last_q_111_io_enq_bits),
    .io_deq_ready(last_q_111_io_deq_ready),
    .io_deq_valid(last_q_111_io_deq_valid),
    .io_deq_bits(last_q_111_io_deq_bits)
  );
  StreamMerger_112 last_merger_112 ( // @[Stab.scala 175:24]
    .clock(last_merger_112_clock),
    .reset(last_merger_112_reset),
    .io_stream1_ready(last_merger_112_io_stream1_ready),
    .io_stream1_valid(last_merger_112_io_stream1_valid),
    .io_stream1_bits(last_merger_112_io_stream1_bits),
    .io_stream2_ready(last_merger_112_io_stream2_ready),
    .io_stream2_valid(last_merger_112_io_stream2_valid),
    .io_stream2_bits(last_merger_112_io_stream2_bits),
    .io_result_ready(last_merger_112_io_result_ready),
    .io_result_valid(last_merger_112_io_result_valid),
    .io_result_bits(last_merger_112_io_result_bits)
  );
  Queue last_q_112 ( // @[Decoupled.scala 361:21]
    .clock(last_q_112_clock),
    .reset(last_q_112_reset),
    .io_enq_ready(last_q_112_io_enq_ready),
    .io_enq_valid(last_q_112_io_enq_valid),
    .io_enq_bits(last_q_112_io_enq_bits),
    .io_deq_ready(last_q_112_io_deq_ready),
    .io_deq_valid(last_q_112_io_deq_valid),
    .io_deq_bits(last_q_112_io_deq_bits)
  );
  StreamMerger_113 last_merger_113 ( // @[Stab.scala 175:24]
    .clock(last_merger_113_clock),
    .reset(last_merger_113_reset),
    .io_stream1_ready(last_merger_113_io_stream1_ready),
    .io_stream1_valid(last_merger_113_io_stream1_valid),
    .io_stream1_bits(last_merger_113_io_stream1_bits),
    .io_stream2_ready(last_merger_113_io_stream2_ready),
    .io_stream2_valid(last_merger_113_io_stream2_valid),
    .io_stream2_bits(last_merger_113_io_stream2_bits),
    .io_result_ready(last_merger_113_io_result_ready),
    .io_result_valid(last_merger_113_io_result_valid),
    .io_result_bits(last_merger_113_io_result_bits)
  );
  Queue last_q_113 ( // @[Decoupled.scala 361:21]
    .clock(last_q_113_clock),
    .reset(last_q_113_reset),
    .io_enq_ready(last_q_113_io_enq_ready),
    .io_enq_valid(last_q_113_io_enq_valid),
    .io_enq_bits(last_q_113_io_enq_bits),
    .io_deq_ready(last_q_113_io_deq_ready),
    .io_deq_valid(last_q_113_io_deq_valid),
    .io_deq_bits(last_q_113_io_deq_bits)
  );
  StreamMerger_114 last_merger_114 ( // @[Stab.scala 175:24]
    .clock(last_merger_114_clock),
    .reset(last_merger_114_reset),
    .io_stream1_ready(last_merger_114_io_stream1_ready),
    .io_stream1_valid(last_merger_114_io_stream1_valid),
    .io_stream1_bits(last_merger_114_io_stream1_bits),
    .io_stream2_ready(last_merger_114_io_stream2_ready),
    .io_stream2_valid(last_merger_114_io_stream2_valid),
    .io_stream2_bits(last_merger_114_io_stream2_bits),
    .io_result_ready(last_merger_114_io_result_ready),
    .io_result_valid(last_merger_114_io_result_valid),
    .io_result_bits(last_merger_114_io_result_bits)
  );
  Queue last_q_114 ( // @[Decoupled.scala 361:21]
    .clock(last_q_114_clock),
    .reset(last_q_114_reset),
    .io_enq_ready(last_q_114_io_enq_ready),
    .io_enq_valid(last_q_114_io_enq_valid),
    .io_enq_bits(last_q_114_io_enq_bits),
    .io_deq_ready(last_q_114_io_deq_ready),
    .io_deq_valid(last_q_114_io_deq_valid),
    .io_deq_bits(last_q_114_io_deq_bits)
  );
  StreamMerger_115 last_merger_115 ( // @[Stab.scala 175:24]
    .clock(last_merger_115_clock),
    .reset(last_merger_115_reset),
    .io_stream1_ready(last_merger_115_io_stream1_ready),
    .io_stream1_valid(last_merger_115_io_stream1_valid),
    .io_stream1_bits(last_merger_115_io_stream1_bits),
    .io_stream2_ready(last_merger_115_io_stream2_ready),
    .io_stream2_valid(last_merger_115_io_stream2_valid),
    .io_stream2_bits(last_merger_115_io_stream2_bits),
    .io_result_ready(last_merger_115_io_result_ready),
    .io_result_valid(last_merger_115_io_result_valid),
    .io_result_bits(last_merger_115_io_result_bits)
  );
  Queue last_q_115 ( // @[Decoupled.scala 361:21]
    .clock(last_q_115_clock),
    .reset(last_q_115_reset),
    .io_enq_ready(last_q_115_io_enq_ready),
    .io_enq_valid(last_q_115_io_enq_valid),
    .io_enq_bits(last_q_115_io_enq_bits),
    .io_deq_ready(last_q_115_io_deq_ready),
    .io_deq_valid(last_q_115_io_deq_valid),
    .io_deq_bits(last_q_115_io_deq_bits)
  );
  StreamMerger_116 last_merger_116 ( // @[Stab.scala 175:24]
    .clock(last_merger_116_clock),
    .reset(last_merger_116_reset),
    .io_stream1_ready(last_merger_116_io_stream1_ready),
    .io_stream1_valid(last_merger_116_io_stream1_valid),
    .io_stream1_bits(last_merger_116_io_stream1_bits),
    .io_stream2_ready(last_merger_116_io_stream2_ready),
    .io_stream2_valid(last_merger_116_io_stream2_valid),
    .io_stream2_bits(last_merger_116_io_stream2_bits),
    .io_result_ready(last_merger_116_io_result_ready),
    .io_result_valid(last_merger_116_io_result_valid),
    .io_result_bits(last_merger_116_io_result_bits)
  );
  Queue last_q_116 ( // @[Decoupled.scala 361:21]
    .clock(last_q_116_clock),
    .reset(last_q_116_reset),
    .io_enq_ready(last_q_116_io_enq_ready),
    .io_enq_valid(last_q_116_io_enq_valid),
    .io_enq_bits(last_q_116_io_enq_bits),
    .io_deq_ready(last_q_116_io_deq_ready),
    .io_deq_valid(last_q_116_io_deq_valid),
    .io_deq_bits(last_q_116_io_deq_bits)
  );
  StreamMerger_117 last_merger_117 ( // @[Stab.scala 175:24]
    .clock(last_merger_117_clock),
    .reset(last_merger_117_reset),
    .io_stream1_ready(last_merger_117_io_stream1_ready),
    .io_stream1_valid(last_merger_117_io_stream1_valid),
    .io_stream1_bits(last_merger_117_io_stream1_bits),
    .io_stream2_ready(last_merger_117_io_stream2_ready),
    .io_stream2_valid(last_merger_117_io_stream2_valid),
    .io_stream2_bits(last_merger_117_io_stream2_bits),
    .io_result_ready(last_merger_117_io_result_ready),
    .io_result_valid(last_merger_117_io_result_valid),
    .io_result_bits(last_merger_117_io_result_bits)
  );
  Queue last_q_117 ( // @[Decoupled.scala 361:21]
    .clock(last_q_117_clock),
    .reset(last_q_117_reset),
    .io_enq_ready(last_q_117_io_enq_ready),
    .io_enq_valid(last_q_117_io_enq_valid),
    .io_enq_bits(last_q_117_io_enq_bits),
    .io_deq_ready(last_q_117_io_deq_ready),
    .io_deq_valid(last_q_117_io_deq_valid),
    .io_deq_bits(last_q_117_io_deq_bits)
  );
  StreamMerger_118 last_merger_118 ( // @[Stab.scala 175:24]
    .clock(last_merger_118_clock),
    .reset(last_merger_118_reset),
    .io_stream1_ready(last_merger_118_io_stream1_ready),
    .io_stream1_valid(last_merger_118_io_stream1_valid),
    .io_stream1_bits(last_merger_118_io_stream1_bits),
    .io_stream2_ready(last_merger_118_io_stream2_ready),
    .io_stream2_valid(last_merger_118_io_stream2_valid),
    .io_stream2_bits(last_merger_118_io_stream2_bits),
    .io_result_ready(last_merger_118_io_result_ready),
    .io_result_valid(last_merger_118_io_result_valid),
    .io_result_bits(last_merger_118_io_result_bits)
  );
  Queue last_q_118 ( // @[Decoupled.scala 361:21]
    .clock(last_q_118_clock),
    .reset(last_q_118_reset),
    .io_enq_ready(last_q_118_io_enq_ready),
    .io_enq_valid(last_q_118_io_enq_valid),
    .io_enq_bits(last_q_118_io_enq_bits),
    .io_deq_ready(last_q_118_io_deq_ready),
    .io_deq_valid(last_q_118_io_deq_valid),
    .io_deq_bits(last_q_118_io_deq_bits)
  );
  StreamMerger_119 last_merger_119 ( // @[Stab.scala 175:24]
    .clock(last_merger_119_clock),
    .reset(last_merger_119_reset),
    .io_stream1_ready(last_merger_119_io_stream1_ready),
    .io_stream1_valid(last_merger_119_io_stream1_valid),
    .io_stream1_bits(last_merger_119_io_stream1_bits),
    .io_stream2_ready(last_merger_119_io_stream2_ready),
    .io_stream2_valid(last_merger_119_io_stream2_valid),
    .io_stream2_bits(last_merger_119_io_stream2_bits),
    .io_result_ready(last_merger_119_io_result_ready),
    .io_result_valid(last_merger_119_io_result_valid),
    .io_result_bits(last_merger_119_io_result_bits)
  );
  Queue last_q_119 ( // @[Decoupled.scala 361:21]
    .clock(last_q_119_clock),
    .reset(last_q_119_reset),
    .io_enq_ready(last_q_119_io_enq_ready),
    .io_enq_valid(last_q_119_io_enq_valid),
    .io_enq_bits(last_q_119_io_enq_bits),
    .io_deq_ready(last_q_119_io_deq_ready),
    .io_deq_valid(last_q_119_io_deq_valid),
    .io_deq_bits(last_q_119_io_deq_bits)
  );
  StreamMerger_120 last_merger_120 ( // @[Stab.scala 175:24]
    .clock(last_merger_120_clock),
    .reset(last_merger_120_reset),
    .io_stream1_ready(last_merger_120_io_stream1_ready),
    .io_stream1_valid(last_merger_120_io_stream1_valid),
    .io_stream1_bits(last_merger_120_io_stream1_bits),
    .io_stream2_ready(last_merger_120_io_stream2_ready),
    .io_stream2_valid(last_merger_120_io_stream2_valid),
    .io_stream2_bits(last_merger_120_io_stream2_bits),
    .io_result_ready(last_merger_120_io_result_ready),
    .io_result_valid(last_merger_120_io_result_valid),
    .io_result_bits(last_merger_120_io_result_bits)
  );
  Queue last_q_120 ( // @[Decoupled.scala 361:21]
    .clock(last_q_120_clock),
    .reset(last_q_120_reset),
    .io_enq_ready(last_q_120_io_enq_ready),
    .io_enq_valid(last_q_120_io_enq_valid),
    .io_enq_bits(last_q_120_io_enq_bits),
    .io_deq_ready(last_q_120_io_deq_ready),
    .io_deq_valid(last_q_120_io_deq_valid),
    .io_deq_bits(last_q_120_io_deq_bits)
  );
  StreamMerger_121 last_merger_121 ( // @[Stab.scala 175:24]
    .clock(last_merger_121_clock),
    .reset(last_merger_121_reset),
    .io_stream1_ready(last_merger_121_io_stream1_ready),
    .io_stream1_valid(last_merger_121_io_stream1_valid),
    .io_stream1_bits(last_merger_121_io_stream1_bits),
    .io_stream2_ready(last_merger_121_io_stream2_ready),
    .io_stream2_valid(last_merger_121_io_stream2_valid),
    .io_stream2_bits(last_merger_121_io_stream2_bits),
    .io_result_ready(last_merger_121_io_result_ready),
    .io_result_valid(last_merger_121_io_result_valid),
    .io_result_bits(last_merger_121_io_result_bits)
  );
  Queue last_q_121 ( // @[Decoupled.scala 361:21]
    .clock(last_q_121_clock),
    .reset(last_q_121_reset),
    .io_enq_ready(last_q_121_io_enq_ready),
    .io_enq_valid(last_q_121_io_enq_valid),
    .io_enq_bits(last_q_121_io_enq_bits),
    .io_deq_ready(last_q_121_io_deq_ready),
    .io_deq_valid(last_q_121_io_deq_valid),
    .io_deq_bits(last_q_121_io_deq_bits)
  );
  StreamMerger_122 last_merger_122 ( // @[Stab.scala 175:24]
    .clock(last_merger_122_clock),
    .reset(last_merger_122_reset),
    .io_stream1_ready(last_merger_122_io_stream1_ready),
    .io_stream1_valid(last_merger_122_io_stream1_valid),
    .io_stream1_bits(last_merger_122_io_stream1_bits),
    .io_stream2_ready(last_merger_122_io_stream2_ready),
    .io_stream2_valid(last_merger_122_io_stream2_valid),
    .io_stream2_bits(last_merger_122_io_stream2_bits),
    .io_result_ready(last_merger_122_io_result_ready),
    .io_result_valid(last_merger_122_io_result_valid),
    .io_result_bits(last_merger_122_io_result_bits)
  );
  Queue last_q_122 ( // @[Decoupled.scala 361:21]
    .clock(last_q_122_clock),
    .reset(last_q_122_reset),
    .io_enq_ready(last_q_122_io_enq_ready),
    .io_enq_valid(last_q_122_io_enq_valid),
    .io_enq_bits(last_q_122_io_enq_bits),
    .io_deq_ready(last_q_122_io_deq_ready),
    .io_deq_valid(last_q_122_io_deq_valid),
    .io_deq_bits(last_q_122_io_deq_bits)
  );
  StreamMerger_123 last_merger_123 ( // @[Stab.scala 175:24]
    .clock(last_merger_123_clock),
    .reset(last_merger_123_reset),
    .io_stream1_ready(last_merger_123_io_stream1_ready),
    .io_stream1_valid(last_merger_123_io_stream1_valid),
    .io_stream1_bits(last_merger_123_io_stream1_bits),
    .io_stream2_ready(last_merger_123_io_stream2_ready),
    .io_stream2_valid(last_merger_123_io_stream2_valid),
    .io_stream2_bits(last_merger_123_io_stream2_bits),
    .io_result_ready(last_merger_123_io_result_ready),
    .io_result_valid(last_merger_123_io_result_valid),
    .io_result_bits(last_merger_123_io_result_bits)
  );
  Queue last_q_123 ( // @[Decoupled.scala 361:21]
    .clock(last_q_123_clock),
    .reset(last_q_123_reset),
    .io_enq_ready(last_q_123_io_enq_ready),
    .io_enq_valid(last_q_123_io_enq_valid),
    .io_enq_bits(last_q_123_io_enq_bits),
    .io_deq_ready(last_q_123_io_deq_ready),
    .io_deq_valid(last_q_123_io_deq_valid),
    .io_deq_bits(last_q_123_io_deq_bits)
  );
  StreamMerger_124 last_merger_124 ( // @[Stab.scala 175:24]
    .clock(last_merger_124_clock),
    .reset(last_merger_124_reset),
    .io_stream1_ready(last_merger_124_io_stream1_ready),
    .io_stream1_valid(last_merger_124_io_stream1_valid),
    .io_stream1_bits(last_merger_124_io_stream1_bits),
    .io_stream2_ready(last_merger_124_io_stream2_ready),
    .io_stream2_valid(last_merger_124_io_stream2_valid),
    .io_stream2_bits(last_merger_124_io_stream2_bits),
    .io_result_ready(last_merger_124_io_result_ready),
    .io_result_valid(last_merger_124_io_result_valid),
    .io_result_bits(last_merger_124_io_result_bits)
  );
  Queue last_q_124 ( // @[Decoupled.scala 361:21]
    .clock(last_q_124_clock),
    .reset(last_q_124_reset),
    .io_enq_ready(last_q_124_io_enq_ready),
    .io_enq_valid(last_q_124_io_enq_valid),
    .io_enq_bits(last_q_124_io_enq_bits),
    .io_deq_ready(last_q_124_io_deq_ready),
    .io_deq_valid(last_q_124_io_deq_valid),
    .io_deq_bits(last_q_124_io_deq_bits)
  );
  StreamMerger_125 last_merger_125 ( // @[Stab.scala 175:24]
    .clock(last_merger_125_clock),
    .reset(last_merger_125_reset),
    .io_stream1_ready(last_merger_125_io_stream1_ready),
    .io_stream1_valid(last_merger_125_io_stream1_valid),
    .io_stream1_bits(last_merger_125_io_stream1_bits),
    .io_stream2_ready(last_merger_125_io_stream2_ready),
    .io_stream2_valid(last_merger_125_io_stream2_valid),
    .io_stream2_bits(last_merger_125_io_stream2_bits),
    .io_result_ready(last_merger_125_io_result_ready),
    .io_result_valid(last_merger_125_io_result_valid),
    .io_result_bits(last_merger_125_io_result_bits)
  );
  Queue last_q_125 ( // @[Decoupled.scala 361:21]
    .clock(last_q_125_clock),
    .reset(last_q_125_reset),
    .io_enq_ready(last_q_125_io_enq_ready),
    .io_enq_valid(last_q_125_io_enq_valid),
    .io_enq_bits(last_q_125_io_enq_bits),
    .io_deq_ready(last_q_125_io_deq_ready),
    .io_deq_valid(last_q_125_io_deq_valid),
    .io_deq_bits(last_q_125_io_deq_bits)
  );
  StreamMerger_126 last_merger_126 ( // @[Stab.scala 175:24]
    .clock(last_merger_126_clock),
    .reset(last_merger_126_reset),
    .io_stream1_ready(last_merger_126_io_stream1_ready),
    .io_stream1_valid(last_merger_126_io_stream1_valid),
    .io_stream1_bits(last_merger_126_io_stream1_bits),
    .io_stream2_ready(last_merger_126_io_stream2_ready),
    .io_stream2_valid(last_merger_126_io_stream2_valid),
    .io_stream2_bits(last_merger_126_io_stream2_bits),
    .io_result_ready(last_merger_126_io_result_ready),
    .io_result_valid(last_merger_126_io_result_valid),
    .io_result_bits(last_merger_126_io_result_bits)
  );
  Queue last_q_126 ( // @[Decoupled.scala 361:21]
    .clock(last_q_126_clock),
    .reset(last_q_126_reset),
    .io_enq_ready(last_q_126_io_enq_ready),
    .io_enq_valid(last_q_126_io_enq_valid),
    .io_enq_bits(last_q_126_io_enq_bits),
    .io_deq_ready(last_q_126_io_deq_ready),
    .io_deq_valid(last_q_126_io_deq_valid),
    .io_deq_bits(last_q_126_io_deq_bits)
  );
  StreamMerger_127 last_merger_127 ( // @[Stab.scala 175:24]
    .clock(last_merger_127_clock),
    .reset(last_merger_127_reset),
    .io_stream1_ready(last_merger_127_io_stream1_ready),
    .io_stream1_valid(last_merger_127_io_stream1_valid),
    .io_stream1_bits(last_merger_127_io_stream1_bits),
    .io_stream2_ready(last_merger_127_io_stream2_ready),
    .io_stream2_valid(last_merger_127_io_stream2_valid),
    .io_stream2_bits(last_merger_127_io_stream2_bits),
    .io_result_ready(last_merger_127_io_result_ready),
    .io_result_valid(last_merger_127_io_result_valid),
    .io_result_bits(last_merger_127_io_result_bits)
  );
  Queue last_q_127 ( // @[Decoupled.scala 361:21]
    .clock(last_q_127_clock),
    .reset(last_q_127_reset),
    .io_enq_ready(last_q_127_io_enq_ready),
    .io_enq_valid(last_q_127_io_enq_valid),
    .io_enq_bits(last_q_127_io_enq_bits),
    .io_deq_ready(last_q_127_io_deq_ready),
    .io_deq_valid(last_q_127_io_deq_valid),
    .io_deq_bits(last_q_127_io_deq_bits)
  );
  StreamMerger_128 last_merger_128 ( // @[Stab.scala 175:24]
    .clock(last_merger_128_clock),
    .reset(last_merger_128_reset),
    .io_stream1_ready(last_merger_128_io_stream1_ready),
    .io_stream1_valid(last_merger_128_io_stream1_valid),
    .io_stream1_bits(last_merger_128_io_stream1_bits),
    .io_stream2_ready(last_merger_128_io_stream2_ready),
    .io_stream2_valid(last_merger_128_io_stream2_valid),
    .io_stream2_bits(last_merger_128_io_stream2_bits),
    .io_result_ready(last_merger_128_io_result_ready),
    .io_result_valid(last_merger_128_io_result_valid),
    .io_result_bits(last_merger_128_io_result_bits)
  );
  Queue last_q_128 ( // @[Decoupled.scala 361:21]
    .clock(last_q_128_clock),
    .reset(last_q_128_reset),
    .io_enq_ready(last_q_128_io_enq_ready),
    .io_enq_valid(last_q_128_io_enq_valid),
    .io_enq_bits(last_q_128_io_enq_bits),
    .io_deq_ready(last_q_128_io_deq_ready),
    .io_deq_valid(last_q_128_io_deq_valid),
    .io_deq_bits(last_q_128_io_deq_bits)
  );
  StreamMerger_129 last_merger_129 ( // @[Stab.scala 175:24]
    .clock(last_merger_129_clock),
    .reset(last_merger_129_reset),
    .io_stream1_ready(last_merger_129_io_stream1_ready),
    .io_stream1_valid(last_merger_129_io_stream1_valid),
    .io_stream1_bits(last_merger_129_io_stream1_bits),
    .io_stream2_ready(last_merger_129_io_stream2_ready),
    .io_stream2_valid(last_merger_129_io_stream2_valid),
    .io_stream2_bits(last_merger_129_io_stream2_bits),
    .io_result_ready(last_merger_129_io_result_ready),
    .io_result_valid(last_merger_129_io_result_valid),
    .io_result_bits(last_merger_129_io_result_bits)
  );
  Queue last_q_129 ( // @[Decoupled.scala 361:21]
    .clock(last_q_129_clock),
    .reset(last_q_129_reset),
    .io_enq_ready(last_q_129_io_enq_ready),
    .io_enq_valid(last_q_129_io_enq_valid),
    .io_enq_bits(last_q_129_io_enq_bits),
    .io_deq_ready(last_q_129_io_deq_ready),
    .io_deq_valid(last_q_129_io_deq_valid),
    .io_deq_bits(last_q_129_io_deq_bits)
  );
  StreamMerger_130 last_merger_130 ( // @[Stab.scala 175:24]
    .clock(last_merger_130_clock),
    .reset(last_merger_130_reset),
    .io_stream1_ready(last_merger_130_io_stream1_ready),
    .io_stream1_valid(last_merger_130_io_stream1_valid),
    .io_stream1_bits(last_merger_130_io_stream1_bits),
    .io_stream2_ready(last_merger_130_io_stream2_ready),
    .io_stream2_valid(last_merger_130_io_stream2_valid),
    .io_stream2_bits(last_merger_130_io_stream2_bits),
    .io_result_ready(last_merger_130_io_result_ready),
    .io_result_valid(last_merger_130_io_result_valid),
    .io_result_bits(last_merger_130_io_result_bits)
  );
  Queue last_q_130 ( // @[Decoupled.scala 361:21]
    .clock(last_q_130_clock),
    .reset(last_q_130_reset),
    .io_enq_ready(last_q_130_io_enq_ready),
    .io_enq_valid(last_q_130_io_enq_valid),
    .io_enq_bits(last_q_130_io_enq_bits),
    .io_deq_ready(last_q_130_io_deq_ready),
    .io_deq_valid(last_q_130_io_deq_valid),
    .io_deq_bits(last_q_130_io_deq_bits)
  );
  StreamMerger_131 last_merger_131 ( // @[Stab.scala 175:24]
    .clock(last_merger_131_clock),
    .reset(last_merger_131_reset),
    .io_stream1_ready(last_merger_131_io_stream1_ready),
    .io_stream1_valid(last_merger_131_io_stream1_valid),
    .io_stream1_bits(last_merger_131_io_stream1_bits),
    .io_stream2_ready(last_merger_131_io_stream2_ready),
    .io_stream2_valid(last_merger_131_io_stream2_valid),
    .io_stream2_bits(last_merger_131_io_stream2_bits),
    .io_result_ready(last_merger_131_io_result_ready),
    .io_result_valid(last_merger_131_io_result_valid),
    .io_result_bits(last_merger_131_io_result_bits)
  );
  Queue last_q_131 ( // @[Decoupled.scala 361:21]
    .clock(last_q_131_clock),
    .reset(last_q_131_reset),
    .io_enq_ready(last_q_131_io_enq_ready),
    .io_enq_valid(last_q_131_io_enq_valid),
    .io_enq_bits(last_q_131_io_enq_bits),
    .io_deq_ready(last_q_131_io_deq_ready),
    .io_deq_valid(last_q_131_io_deq_valid),
    .io_deq_bits(last_q_131_io_deq_bits)
  );
  StreamMerger_132 last_merger_132 ( // @[Stab.scala 175:24]
    .clock(last_merger_132_clock),
    .reset(last_merger_132_reset),
    .io_stream1_ready(last_merger_132_io_stream1_ready),
    .io_stream1_valid(last_merger_132_io_stream1_valid),
    .io_stream1_bits(last_merger_132_io_stream1_bits),
    .io_stream2_ready(last_merger_132_io_stream2_ready),
    .io_stream2_valid(last_merger_132_io_stream2_valid),
    .io_stream2_bits(last_merger_132_io_stream2_bits),
    .io_result_ready(last_merger_132_io_result_ready),
    .io_result_valid(last_merger_132_io_result_valid),
    .io_result_bits(last_merger_132_io_result_bits)
  );
  Queue last_q_132 ( // @[Decoupled.scala 361:21]
    .clock(last_q_132_clock),
    .reset(last_q_132_reset),
    .io_enq_ready(last_q_132_io_enq_ready),
    .io_enq_valid(last_q_132_io_enq_valid),
    .io_enq_bits(last_q_132_io_enq_bits),
    .io_deq_ready(last_q_132_io_deq_ready),
    .io_deq_valid(last_q_132_io_deq_valid),
    .io_deq_bits(last_q_132_io_deq_bits)
  );
  StreamMerger_133 last_merger_133 ( // @[Stab.scala 175:24]
    .clock(last_merger_133_clock),
    .reset(last_merger_133_reset),
    .io_stream1_ready(last_merger_133_io_stream1_ready),
    .io_stream1_valid(last_merger_133_io_stream1_valid),
    .io_stream1_bits(last_merger_133_io_stream1_bits),
    .io_stream2_ready(last_merger_133_io_stream2_ready),
    .io_stream2_valid(last_merger_133_io_stream2_valid),
    .io_stream2_bits(last_merger_133_io_stream2_bits),
    .io_result_ready(last_merger_133_io_result_ready),
    .io_result_valid(last_merger_133_io_result_valid),
    .io_result_bits(last_merger_133_io_result_bits)
  );
  Queue last_q_133 ( // @[Decoupled.scala 361:21]
    .clock(last_q_133_clock),
    .reset(last_q_133_reset),
    .io_enq_ready(last_q_133_io_enq_ready),
    .io_enq_valid(last_q_133_io_enq_valid),
    .io_enq_bits(last_q_133_io_enq_bits),
    .io_deq_ready(last_q_133_io_deq_ready),
    .io_deq_valid(last_q_133_io_deq_valid),
    .io_deq_bits(last_q_133_io_deq_bits)
  );
  StreamMerger_134 last_merger_134 ( // @[Stab.scala 175:24]
    .clock(last_merger_134_clock),
    .reset(last_merger_134_reset),
    .io_stream1_ready(last_merger_134_io_stream1_ready),
    .io_stream1_valid(last_merger_134_io_stream1_valid),
    .io_stream1_bits(last_merger_134_io_stream1_bits),
    .io_stream2_ready(last_merger_134_io_stream2_ready),
    .io_stream2_valid(last_merger_134_io_stream2_valid),
    .io_stream2_bits(last_merger_134_io_stream2_bits),
    .io_result_ready(last_merger_134_io_result_ready),
    .io_result_valid(last_merger_134_io_result_valid),
    .io_result_bits(last_merger_134_io_result_bits)
  );
  Queue last_q_134 ( // @[Decoupled.scala 361:21]
    .clock(last_q_134_clock),
    .reset(last_q_134_reset),
    .io_enq_ready(last_q_134_io_enq_ready),
    .io_enq_valid(last_q_134_io_enq_valid),
    .io_enq_bits(last_q_134_io_enq_bits),
    .io_deq_ready(last_q_134_io_deq_ready),
    .io_deq_valid(last_q_134_io_deq_valid),
    .io_deq_bits(last_q_134_io_deq_bits)
  );
  StreamMerger_135 last_merger_135 ( // @[Stab.scala 175:24]
    .clock(last_merger_135_clock),
    .reset(last_merger_135_reset),
    .io_stream1_ready(last_merger_135_io_stream1_ready),
    .io_stream1_valid(last_merger_135_io_stream1_valid),
    .io_stream1_bits(last_merger_135_io_stream1_bits),
    .io_stream2_ready(last_merger_135_io_stream2_ready),
    .io_stream2_valid(last_merger_135_io_stream2_valid),
    .io_stream2_bits(last_merger_135_io_stream2_bits),
    .io_result_ready(last_merger_135_io_result_ready),
    .io_result_valid(last_merger_135_io_result_valid),
    .io_result_bits(last_merger_135_io_result_bits)
  );
  Queue last_q_135 ( // @[Decoupled.scala 361:21]
    .clock(last_q_135_clock),
    .reset(last_q_135_reset),
    .io_enq_ready(last_q_135_io_enq_ready),
    .io_enq_valid(last_q_135_io_enq_valid),
    .io_enq_bits(last_q_135_io_enq_bits),
    .io_deq_ready(last_q_135_io_deq_ready),
    .io_deq_valid(last_q_135_io_deq_valid),
    .io_deq_bits(last_q_135_io_deq_bits)
  );
  StreamMerger_136 last_merger_136 ( // @[Stab.scala 175:24]
    .clock(last_merger_136_clock),
    .reset(last_merger_136_reset),
    .io_stream1_ready(last_merger_136_io_stream1_ready),
    .io_stream1_valid(last_merger_136_io_stream1_valid),
    .io_stream1_bits(last_merger_136_io_stream1_bits),
    .io_stream2_ready(last_merger_136_io_stream2_ready),
    .io_stream2_valid(last_merger_136_io_stream2_valid),
    .io_stream2_bits(last_merger_136_io_stream2_bits),
    .io_result_ready(last_merger_136_io_result_ready),
    .io_result_valid(last_merger_136_io_result_valid),
    .io_result_bits(last_merger_136_io_result_bits)
  );
  Queue last_q_136 ( // @[Decoupled.scala 361:21]
    .clock(last_q_136_clock),
    .reset(last_q_136_reset),
    .io_enq_ready(last_q_136_io_enq_ready),
    .io_enq_valid(last_q_136_io_enq_valid),
    .io_enq_bits(last_q_136_io_enq_bits),
    .io_deq_ready(last_q_136_io_deq_ready),
    .io_deq_valid(last_q_136_io_deq_valid),
    .io_deq_bits(last_q_136_io_deq_bits)
  );
  StreamMerger_137 last_merger_137 ( // @[Stab.scala 175:24]
    .clock(last_merger_137_clock),
    .reset(last_merger_137_reset),
    .io_stream1_ready(last_merger_137_io_stream1_ready),
    .io_stream1_valid(last_merger_137_io_stream1_valid),
    .io_stream1_bits(last_merger_137_io_stream1_bits),
    .io_stream2_ready(last_merger_137_io_stream2_ready),
    .io_stream2_valid(last_merger_137_io_stream2_valid),
    .io_stream2_bits(last_merger_137_io_stream2_bits),
    .io_result_ready(last_merger_137_io_result_ready),
    .io_result_valid(last_merger_137_io_result_valid),
    .io_result_bits(last_merger_137_io_result_bits)
  );
  Queue last_q_137 ( // @[Decoupled.scala 361:21]
    .clock(last_q_137_clock),
    .reset(last_q_137_reset),
    .io_enq_ready(last_q_137_io_enq_ready),
    .io_enq_valid(last_q_137_io_enq_valid),
    .io_enq_bits(last_q_137_io_enq_bits),
    .io_deq_ready(last_q_137_io_deq_ready),
    .io_deq_valid(last_q_137_io_deq_valid),
    .io_deq_bits(last_q_137_io_deq_bits)
  );
  StreamMerger_138 last_merger_138 ( // @[Stab.scala 175:24]
    .clock(last_merger_138_clock),
    .reset(last_merger_138_reset),
    .io_stream1_ready(last_merger_138_io_stream1_ready),
    .io_stream1_valid(last_merger_138_io_stream1_valid),
    .io_stream1_bits(last_merger_138_io_stream1_bits),
    .io_stream2_ready(last_merger_138_io_stream2_ready),
    .io_stream2_valid(last_merger_138_io_stream2_valid),
    .io_stream2_bits(last_merger_138_io_stream2_bits),
    .io_result_ready(last_merger_138_io_result_ready),
    .io_result_valid(last_merger_138_io_result_valid),
    .io_result_bits(last_merger_138_io_result_bits)
  );
  Queue last_q_138 ( // @[Decoupled.scala 361:21]
    .clock(last_q_138_clock),
    .reset(last_q_138_reset),
    .io_enq_ready(last_q_138_io_enq_ready),
    .io_enq_valid(last_q_138_io_enq_valid),
    .io_enq_bits(last_q_138_io_enq_bits),
    .io_deq_ready(last_q_138_io_deq_ready),
    .io_deq_valid(last_q_138_io_deq_valid),
    .io_deq_bits(last_q_138_io_deq_bits)
  );
  StreamMerger_139 last_merger_139 ( // @[Stab.scala 175:24]
    .clock(last_merger_139_clock),
    .reset(last_merger_139_reset),
    .io_stream1_ready(last_merger_139_io_stream1_ready),
    .io_stream1_valid(last_merger_139_io_stream1_valid),
    .io_stream1_bits(last_merger_139_io_stream1_bits),
    .io_stream2_ready(last_merger_139_io_stream2_ready),
    .io_stream2_valid(last_merger_139_io_stream2_valid),
    .io_stream2_bits(last_merger_139_io_stream2_bits),
    .io_result_ready(last_merger_139_io_result_ready),
    .io_result_valid(last_merger_139_io_result_valid),
    .io_result_bits(last_merger_139_io_result_bits)
  );
  Queue last_q_139 ( // @[Decoupled.scala 361:21]
    .clock(last_q_139_clock),
    .reset(last_q_139_reset),
    .io_enq_ready(last_q_139_io_enq_ready),
    .io_enq_valid(last_q_139_io_enq_valid),
    .io_enq_bits(last_q_139_io_enq_bits),
    .io_deq_ready(last_q_139_io_deq_ready),
    .io_deq_valid(last_q_139_io_deq_valid),
    .io_deq_bits(last_q_139_io_deq_bits)
  );
  StreamMerger_140 last_merger_140 ( // @[Stab.scala 175:24]
    .clock(last_merger_140_clock),
    .reset(last_merger_140_reset),
    .io_stream1_ready(last_merger_140_io_stream1_ready),
    .io_stream1_valid(last_merger_140_io_stream1_valid),
    .io_stream1_bits(last_merger_140_io_stream1_bits),
    .io_stream2_ready(last_merger_140_io_stream2_ready),
    .io_stream2_valid(last_merger_140_io_stream2_valid),
    .io_stream2_bits(last_merger_140_io_stream2_bits),
    .io_result_ready(last_merger_140_io_result_ready),
    .io_result_valid(last_merger_140_io_result_valid),
    .io_result_bits(last_merger_140_io_result_bits)
  );
  Queue last_q_140 ( // @[Decoupled.scala 361:21]
    .clock(last_q_140_clock),
    .reset(last_q_140_reset),
    .io_enq_ready(last_q_140_io_enq_ready),
    .io_enq_valid(last_q_140_io_enq_valid),
    .io_enq_bits(last_q_140_io_enq_bits),
    .io_deq_ready(last_q_140_io_deq_ready),
    .io_deq_valid(last_q_140_io_deq_valid),
    .io_deq_bits(last_q_140_io_deq_bits)
  );
  StreamMerger_141 last_merger_141 ( // @[Stab.scala 175:24]
    .clock(last_merger_141_clock),
    .reset(last_merger_141_reset),
    .io_stream1_ready(last_merger_141_io_stream1_ready),
    .io_stream1_valid(last_merger_141_io_stream1_valid),
    .io_stream1_bits(last_merger_141_io_stream1_bits),
    .io_stream2_ready(last_merger_141_io_stream2_ready),
    .io_stream2_valid(last_merger_141_io_stream2_valid),
    .io_stream2_bits(last_merger_141_io_stream2_bits),
    .io_result_ready(last_merger_141_io_result_ready),
    .io_result_valid(last_merger_141_io_result_valid),
    .io_result_bits(last_merger_141_io_result_bits)
  );
  Queue last_q_141 ( // @[Decoupled.scala 361:21]
    .clock(last_q_141_clock),
    .reset(last_q_141_reset),
    .io_enq_ready(last_q_141_io_enq_ready),
    .io_enq_valid(last_q_141_io_enq_valid),
    .io_enq_bits(last_q_141_io_enq_bits),
    .io_deq_ready(last_q_141_io_deq_ready),
    .io_deq_valid(last_q_141_io_deq_valid),
    .io_deq_bits(last_q_141_io_deq_bits)
  );
  StreamMerger_142 last_merger_142 ( // @[Stab.scala 175:24]
    .clock(last_merger_142_clock),
    .reset(last_merger_142_reset),
    .io_stream1_ready(last_merger_142_io_stream1_ready),
    .io_stream1_valid(last_merger_142_io_stream1_valid),
    .io_stream1_bits(last_merger_142_io_stream1_bits),
    .io_stream2_ready(last_merger_142_io_stream2_ready),
    .io_stream2_valid(last_merger_142_io_stream2_valid),
    .io_stream2_bits(last_merger_142_io_stream2_bits),
    .io_result_ready(last_merger_142_io_result_ready),
    .io_result_valid(last_merger_142_io_result_valid),
    .io_result_bits(last_merger_142_io_result_bits)
  );
  Queue last_q_142 ( // @[Decoupled.scala 361:21]
    .clock(last_q_142_clock),
    .reset(last_q_142_reset),
    .io_enq_ready(last_q_142_io_enq_ready),
    .io_enq_valid(last_q_142_io_enq_valid),
    .io_enq_bits(last_q_142_io_enq_bits),
    .io_deq_ready(last_q_142_io_deq_ready),
    .io_deq_valid(last_q_142_io_deq_valid),
    .io_deq_bits(last_q_142_io_deq_bits)
  );
  StreamMerger_143 last_merger_143 ( // @[Stab.scala 175:24]
    .clock(last_merger_143_clock),
    .reset(last_merger_143_reset),
    .io_stream1_ready(last_merger_143_io_stream1_ready),
    .io_stream1_valid(last_merger_143_io_stream1_valid),
    .io_stream1_bits(last_merger_143_io_stream1_bits),
    .io_stream2_ready(last_merger_143_io_stream2_ready),
    .io_stream2_valid(last_merger_143_io_stream2_valid),
    .io_stream2_bits(last_merger_143_io_stream2_bits),
    .io_result_ready(last_merger_143_io_result_ready),
    .io_result_valid(last_merger_143_io_result_valid),
    .io_result_bits(last_merger_143_io_result_bits)
  );
  Queue last_q_143 ( // @[Decoupled.scala 361:21]
    .clock(last_q_143_clock),
    .reset(last_q_143_reset),
    .io_enq_ready(last_q_143_io_enq_ready),
    .io_enq_valid(last_q_143_io_enq_valid),
    .io_enq_bits(last_q_143_io_enq_bits),
    .io_deq_ready(last_q_143_io_deq_ready),
    .io_deq_valid(last_q_143_io_deq_valid),
    .io_deq_bits(last_q_143_io_deq_bits)
  );
  StreamMerger_144 last_merger_144 ( // @[Stab.scala 175:24]
    .clock(last_merger_144_clock),
    .reset(last_merger_144_reset),
    .io_stream1_ready(last_merger_144_io_stream1_ready),
    .io_stream1_valid(last_merger_144_io_stream1_valid),
    .io_stream1_bits(last_merger_144_io_stream1_bits),
    .io_stream2_ready(last_merger_144_io_stream2_ready),
    .io_stream2_valid(last_merger_144_io_stream2_valid),
    .io_stream2_bits(last_merger_144_io_stream2_bits),
    .io_result_ready(last_merger_144_io_result_ready),
    .io_result_valid(last_merger_144_io_result_valid),
    .io_result_bits(last_merger_144_io_result_bits)
  );
  Queue last_q_144 ( // @[Decoupled.scala 361:21]
    .clock(last_q_144_clock),
    .reset(last_q_144_reset),
    .io_enq_ready(last_q_144_io_enq_ready),
    .io_enq_valid(last_q_144_io_enq_valid),
    .io_enq_bits(last_q_144_io_enq_bits),
    .io_deq_ready(last_q_144_io_deq_ready),
    .io_deq_valid(last_q_144_io_deq_valid),
    .io_deq_bits(last_q_144_io_deq_bits)
  );
  StreamMerger_145 last_merger_145 ( // @[Stab.scala 175:24]
    .clock(last_merger_145_clock),
    .reset(last_merger_145_reset),
    .io_stream1_ready(last_merger_145_io_stream1_ready),
    .io_stream1_valid(last_merger_145_io_stream1_valid),
    .io_stream1_bits(last_merger_145_io_stream1_bits),
    .io_stream2_ready(last_merger_145_io_stream2_ready),
    .io_stream2_valid(last_merger_145_io_stream2_valid),
    .io_stream2_bits(last_merger_145_io_stream2_bits),
    .io_result_ready(last_merger_145_io_result_ready),
    .io_result_valid(last_merger_145_io_result_valid),
    .io_result_bits(last_merger_145_io_result_bits)
  );
  Queue last_q_145 ( // @[Decoupled.scala 361:21]
    .clock(last_q_145_clock),
    .reset(last_q_145_reset),
    .io_enq_ready(last_q_145_io_enq_ready),
    .io_enq_valid(last_q_145_io_enq_valid),
    .io_enq_bits(last_q_145_io_enq_bits),
    .io_deq_ready(last_q_145_io_deq_ready),
    .io_deq_valid(last_q_145_io_deq_valid),
    .io_deq_bits(last_q_145_io_deq_bits)
  );
  StreamMerger_146 last_merger_146 ( // @[Stab.scala 175:24]
    .clock(last_merger_146_clock),
    .reset(last_merger_146_reset),
    .io_stream1_ready(last_merger_146_io_stream1_ready),
    .io_stream1_valid(last_merger_146_io_stream1_valid),
    .io_stream1_bits(last_merger_146_io_stream1_bits),
    .io_stream2_ready(last_merger_146_io_stream2_ready),
    .io_stream2_valid(last_merger_146_io_stream2_valid),
    .io_stream2_bits(last_merger_146_io_stream2_bits),
    .io_result_ready(last_merger_146_io_result_ready),
    .io_result_valid(last_merger_146_io_result_valid),
    .io_result_bits(last_merger_146_io_result_bits)
  );
  Queue last_q_146 ( // @[Decoupled.scala 361:21]
    .clock(last_q_146_clock),
    .reset(last_q_146_reset),
    .io_enq_ready(last_q_146_io_enq_ready),
    .io_enq_valid(last_q_146_io_enq_valid),
    .io_enq_bits(last_q_146_io_enq_bits),
    .io_deq_ready(last_q_146_io_deq_ready),
    .io_deq_valid(last_q_146_io_deq_valid),
    .io_deq_bits(last_q_146_io_deq_bits)
  );
  StreamMerger_147 last_merger_147 ( // @[Stab.scala 175:24]
    .clock(last_merger_147_clock),
    .reset(last_merger_147_reset),
    .io_stream1_ready(last_merger_147_io_stream1_ready),
    .io_stream1_valid(last_merger_147_io_stream1_valid),
    .io_stream1_bits(last_merger_147_io_stream1_bits),
    .io_stream2_ready(last_merger_147_io_stream2_ready),
    .io_stream2_valid(last_merger_147_io_stream2_valid),
    .io_stream2_bits(last_merger_147_io_stream2_bits),
    .io_result_ready(last_merger_147_io_result_ready),
    .io_result_valid(last_merger_147_io_result_valid),
    .io_result_bits(last_merger_147_io_result_bits)
  );
  Queue last_q_147 ( // @[Decoupled.scala 361:21]
    .clock(last_q_147_clock),
    .reset(last_q_147_reset),
    .io_enq_ready(last_q_147_io_enq_ready),
    .io_enq_valid(last_q_147_io_enq_valid),
    .io_enq_bits(last_q_147_io_enq_bits),
    .io_deq_ready(last_q_147_io_deq_ready),
    .io_deq_valid(last_q_147_io_deq_valid),
    .io_deq_bits(last_q_147_io_deq_bits)
  );
  StreamMerger_148 last_merger_148 ( // @[Stab.scala 175:24]
    .clock(last_merger_148_clock),
    .reset(last_merger_148_reset),
    .io_stream1_ready(last_merger_148_io_stream1_ready),
    .io_stream1_valid(last_merger_148_io_stream1_valid),
    .io_stream1_bits(last_merger_148_io_stream1_bits),
    .io_stream2_ready(last_merger_148_io_stream2_ready),
    .io_stream2_valid(last_merger_148_io_stream2_valid),
    .io_stream2_bits(last_merger_148_io_stream2_bits),
    .io_result_ready(last_merger_148_io_result_ready),
    .io_result_valid(last_merger_148_io_result_valid),
    .io_result_bits(last_merger_148_io_result_bits)
  );
  Queue last_q_148 ( // @[Decoupled.scala 361:21]
    .clock(last_q_148_clock),
    .reset(last_q_148_reset),
    .io_enq_ready(last_q_148_io_enq_ready),
    .io_enq_valid(last_q_148_io_enq_valid),
    .io_enq_bits(last_q_148_io_enq_bits),
    .io_deq_ready(last_q_148_io_deq_ready),
    .io_deq_valid(last_q_148_io_deq_valid),
    .io_deq_bits(last_q_148_io_deq_bits)
  );
  StreamMerger_149 last_merger_149 ( // @[Stab.scala 175:24]
    .clock(last_merger_149_clock),
    .reset(last_merger_149_reset),
    .io_stream1_ready(last_merger_149_io_stream1_ready),
    .io_stream1_valid(last_merger_149_io_stream1_valid),
    .io_stream1_bits(last_merger_149_io_stream1_bits),
    .io_stream2_ready(last_merger_149_io_stream2_ready),
    .io_stream2_valid(last_merger_149_io_stream2_valid),
    .io_stream2_bits(last_merger_149_io_stream2_bits),
    .io_result_ready(last_merger_149_io_result_ready),
    .io_result_valid(last_merger_149_io_result_valid),
    .io_result_bits(last_merger_149_io_result_bits)
  );
  Queue last_q_149 ( // @[Decoupled.scala 361:21]
    .clock(last_q_149_clock),
    .reset(last_q_149_reset),
    .io_enq_ready(last_q_149_io_enq_ready),
    .io_enq_valid(last_q_149_io_enq_valid),
    .io_enq_bits(last_q_149_io_enq_bits),
    .io_deq_ready(last_q_149_io_deq_ready),
    .io_deq_valid(last_q_149_io_deq_valid),
    .io_deq_bits(last_q_149_io_deq_bits)
  );
  StreamMerger_150 last_merger_150 ( // @[Stab.scala 175:24]
    .clock(last_merger_150_clock),
    .reset(last_merger_150_reset),
    .io_stream1_ready(last_merger_150_io_stream1_ready),
    .io_stream1_valid(last_merger_150_io_stream1_valid),
    .io_stream1_bits(last_merger_150_io_stream1_bits),
    .io_stream2_ready(last_merger_150_io_stream2_ready),
    .io_stream2_valid(last_merger_150_io_stream2_valid),
    .io_stream2_bits(last_merger_150_io_stream2_bits),
    .io_result_ready(last_merger_150_io_result_ready),
    .io_result_valid(last_merger_150_io_result_valid),
    .io_result_bits(last_merger_150_io_result_bits)
  );
  Queue last_q_150 ( // @[Decoupled.scala 361:21]
    .clock(last_q_150_clock),
    .reset(last_q_150_reset),
    .io_enq_ready(last_q_150_io_enq_ready),
    .io_enq_valid(last_q_150_io_enq_valid),
    .io_enq_bits(last_q_150_io_enq_bits),
    .io_deq_ready(last_q_150_io_deq_ready),
    .io_deq_valid(last_q_150_io_deq_valid),
    .io_deq_bits(last_q_150_io_deq_bits)
  );
  StreamMerger_151 last_merger_151 ( // @[Stab.scala 175:24]
    .clock(last_merger_151_clock),
    .reset(last_merger_151_reset),
    .io_stream1_ready(last_merger_151_io_stream1_ready),
    .io_stream1_valid(last_merger_151_io_stream1_valid),
    .io_stream1_bits(last_merger_151_io_stream1_bits),
    .io_stream2_ready(last_merger_151_io_stream2_ready),
    .io_stream2_valid(last_merger_151_io_stream2_valid),
    .io_stream2_bits(last_merger_151_io_stream2_bits),
    .io_result_ready(last_merger_151_io_result_ready),
    .io_result_valid(last_merger_151_io_result_valid),
    .io_result_bits(last_merger_151_io_result_bits)
  );
  Queue last_q_151 ( // @[Decoupled.scala 361:21]
    .clock(last_q_151_clock),
    .reset(last_q_151_reset),
    .io_enq_ready(last_q_151_io_enq_ready),
    .io_enq_valid(last_q_151_io_enq_valid),
    .io_enq_bits(last_q_151_io_enq_bits),
    .io_deq_ready(last_q_151_io_deq_ready),
    .io_deq_valid(last_q_151_io_deq_valid),
    .io_deq_bits(last_q_151_io_deq_bits)
  );
  StreamMerger_152 last_merger_152 ( // @[Stab.scala 175:24]
    .clock(last_merger_152_clock),
    .reset(last_merger_152_reset),
    .io_stream1_ready(last_merger_152_io_stream1_ready),
    .io_stream1_valid(last_merger_152_io_stream1_valid),
    .io_stream1_bits(last_merger_152_io_stream1_bits),
    .io_stream2_ready(last_merger_152_io_stream2_ready),
    .io_stream2_valid(last_merger_152_io_stream2_valid),
    .io_stream2_bits(last_merger_152_io_stream2_bits),
    .io_result_ready(last_merger_152_io_result_ready),
    .io_result_valid(last_merger_152_io_result_valid),
    .io_result_bits(last_merger_152_io_result_bits)
  );
  Queue last_q_152 ( // @[Decoupled.scala 361:21]
    .clock(last_q_152_clock),
    .reset(last_q_152_reset),
    .io_enq_ready(last_q_152_io_enq_ready),
    .io_enq_valid(last_q_152_io_enq_valid),
    .io_enq_bits(last_q_152_io_enq_bits),
    .io_deq_ready(last_q_152_io_deq_ready),
    .io_deq_valid(last_q_152_io_deq_valid),
    .io_deq_bits(last_q_152_io_deq_bits)
  );
  StreamMerger_153 last_merger_153 ( // @[Stab.scala 175:24]
    .clock(last_merger_153_clock),
    .reset(last_merger_153_reset),
    .io_stream1_ready(last_merger_153_io_stream1_ready),
    .io_stream1_valid(last_merger_153_io_stream1_valid),
    .io_stream1_bits(last_merger_153_io_stream1_bits),
    .io_stream2_ready(last_merger_153_io_stream2_ready),
    .io_stream2_valid(last_merger_153_io_stream2_valid),
    .io_stream2_bits(last_merger_153_io_stream2_bits),
    .io_result_ready(last_merger_153_io_result_ready),
    .io_result_valid(last_merger_153_io_result_valid),
    .io_result_bits(last_merger_153_io_result_bits)
  );
  Queue last_q_153 ( // @[Decoupled.scala 361:21]
    .clock(last_q_153_clock),
    .reset(last_q_153_reset),
    .io_enq_ready(last_q_153_io_enq_ready),
    .io_enq_valid(last_q_153_io_enq_valid),
    .io_enq_bits(last_q_153_io_enq_bits),
    .io_deq_ready(last_q_153_io_deq_ready),
    .io_deq_valid(last_q_153_io_deq_valid),
    .io_deq_bits(last_q_153_io_deq_bits)
  );
  StreamMerger_154 last_merger_154 ( // @[Stab.scala 175:24]
    .clock(last_merger_154_clock),
    .reset(last_merger_154_reset),
    .io_stream1_ready(last_merger_154_io_stream1_ready),
    .io_stream1_valid(last_merger_154_io_stream1_valid),
    .io_stream1_bits(last_merger_154_io_stream1_bits),
    .io_stream2_ready(last_merger_154_io_stream2_ready),
    .io_stream2_valid(last_merger_154_io_stream2_valid),
    .io_stream2_bits(last_merger_154_io_stream2_bits),
    .io_result_ready(last_merger_154_io_result_ready),
    .io_result_valid(last_merger_154_io_result_valid),
    .io_result_bits(last_merger_154_io_result_bits)
  );
  Queue last_q_154 ( // @[Decoupled.scala 361:21]
    .clock(last_q_154_clock),
    .reset(last_q_154_reset),
    .io_enq_ready(last_q_154_io_enq_ready),
    .io_enq_valid(last_q_154_io_enq_valid),
    .io_enq_bits(last_q_154_io_enq_bits),
    .io_deq_ready(last_q_154_io_deq_ready),
    .io_deq_valid(last_q_154_io_deq_valid),
    .io_deq_bits(last_q_154_io_deq_bits)
  );
  StreamMerger_155 last_merger_155 ( // @[Stab.scala 175:24]
    .clock(last_merger_155_clock),
    .reset(last_merger_155_reset),
    .io_stream1_ready(last_merger_155_io_stream1_ready),
    .io_stream1_valid(last_merger_155_io_stream1_valid),
    .io_stream1_bits(last_merger_155_io_stream1_bits),
    .io_stream2_ready(last_merger_155_io_stream2_ready),
    .io_stream2_valid(last_merger_155_io_stream2_valid),
    .io_stream2_bits(last_merger_155_io_stream2_bits),
    .io_result_ready(last_merger_155_io_result_ready),
    .io_result_valid(last_merger_155_io_result_valid),
    .io_result_bits(last_merger_155_io_result_bits)
  );
  Queue last_q_155 ( // @[Decoupled.scala 361:21]
    .clock(last_q_155_clock),
    .reset(last_q_155_reset),
    .io_enq_ready(last_q_155_io_enq_ready),
    .io_enq_valid(last_q_155_io_enq_valid),
    .io_enq_bits(last_q_155_io_enq_bits),
    .io_deq_ready(last_q_155_io_deq_ready),
    .io_deq_valid(last_q_155_io_deq_valid),
    .io_deq_bits(last_q_155_io_deq_bits)
  );
  StreamMerger_156 last_merger_156 ( // @[Stab.scala 175:24]
    .clock(last_merger_156_clock),
    .reset(last_merger_156_reset),
    .io_stream1_ready(last_merger_156_io_stream1_ready),
    .io_stream1_valid(last_merger_156_io_stream1_valid),
    .io_stream1_bits(last_merger_156_io_stream1_bits),
    .io_stream2_ready(last_merger_156_io_stream2_ready),
    .io_stream2_valid(last_merger_156_io_stream2_valid),
    .io_stream2_bits(last_merger_156_io_stream2_bits),
    .io_result_ready(last_merger_156_io_result_ready),
    .io_result_valid(last_merger_156_io_result_valid),
    .io_result_bits(last_merger_156_io_result_bits)
  );
  Queue last_q_156 ( // @[Decoupled.scala 361:21]
    .clock(last_q_156_clock),
    .reset(last_q_156_reset),
    .io_enq_ready(last_q_156_io_enq_ready),
    .io_enq_valid(last_q_156_io_enq_valid),
    .io_enq_bits(last_q_156_io_enq_bits),
    .io_deq_ready(last_q_156_io_deq_ready),
    .io_deq_valid(last_q_156_io_deq_valid),
    .io_deq_bits(last_q_156_io_deq_bits)
  );
  StreamMerger_157 last_merger_157 ( // @[Stab.scala 175:24]
    .clock(last_merger_157_clock),
    .reset(last_merger_157_reset),
    .io_stream1_ready(last_merger_157_io_stream1_ready),
    .io_stream1_valid(last_merger_157_io_stream1_valid),
    .io_stream1_bits(last_merger_157_io_stream1_bits),
    .io_stream2_ready(last_merger_157_io_stream2_ready),
    .io_stream2_valid(last_merger_157_io_stream2_valid),
    .io_stream2_bits(last_merger_157_io_stream2_bits),
    .io_result_ready(last_merger_157_io_result_ready),
    .io_result_valid(last_merger_157_io_result_valid),
    .io_result_bits(last_merger_157_io_result_bits)
  );
  Queue last_q_157 ( // @[Decoupled.scala 361:21]
    .clock(last_q_157_clock),
    .reset(last_q_157_reset),
    .io_enq_ready(last_q_157_io_enq_ready),
    .io_enq_valid(last_q_157_io_enq_valid),
    .io_enq_bits(last_q_157_io_enq_bits),
    .io_deq_ready(last_q_157_io_deq_ready),
    .io_deq_valid(last_q_157_io_deq_valid),
    .io_deq_bits(last_q_157_io_deq_bits)
  );
  StreamMerger_158 last_merger_158 ( // @[Stab.scala 175:24]
    .clock(last_merger_158_clock),
    .reset(last_merger_158_reset),
    .io_stream1_ready(last_merger_158_io_stream1_ready),
    .io_stream1_valid(last_merger_158_io_stream1_valid),
    .io_stream1_bits(last_merger_158_io_stream1_bits),
    .io_stream2_ready(last_merger_158_io_stream2_ready),
    .io_stream2_valid(last_merger_158_io_stream2_valid),
    .io_stream2_bits(last_merger_158_io_stream2_bits),
    .io_result_ready(last_merger_158_io_result_ready),
    .io_result_valid(last_merger_158_io_result_valid),
    .io_result_bits(last_merger_158_io_result_bits)
  );
  Queue last_q_158 ( // @[Decoupled.scala 361:21]
    .clock(last_q_158_clock),
    .reset(last_q_158_reset),
    .io_enq_ready(last_q_158_io_enq_ready),
    .io_enq_valid(last_q_158_io_enq_valid),
    .io_enq_bits(last_q_158_io_enq_bits),
    .io_deq_ready(last_q_158_io_deq_ready),
    .io_deq_valid(last_q_158_io_deq_valid),
    .io_deq_bits(last_q_158_io_deq_bits)
  );
  StreamMerger_159 last_merger_159 ( // @[Stab.scala 175:24]
    .clock(last_merger_159_clock),
    .reset(last_merger_159_reset),
    .io_stream1_ready(last_merger_159_io_stream1_ready),
    .io_stream1_valid(last_merger_159_io_stream1_valid),
    .io_stream1_bits(last_merger_159_io_stream1_bits),
    .io_stream2_ready(last_merger_159_io_stream2_ready),
    .io_stream2_valid(last_merger_159_io_stream2_valid),
    .io_stream2_bits(last_merger_159_io_stream2_bits),
    .io_result_ready(last_merger_159_io_result_ready),
    .io_result_valid(last_merger_159_io_result_valid),
    .io_result_bits(last_merger_159_io_result_bits)
  );
  Queue last_q_159 ( // @[Decoupled.scala 361:21]
    .clock(last_q_159_clock),
    .reset(last_q_159_reset),
    .io_enq_ready(last_q_159_io_enq_ready),
    .io_enq_valid(last_q_159_io_enq_valid),
    .io_enq_bits(last_q_159_io_enq_bits),
    .io_deq_ready(last_q_159_io_deq_ready),
    .io_deq_valid(last_q_159_io_deq_valid),
    .io_deq_bits(last_q_159_io_deq_bits)
  );
  StreamMerger_160 last_merger_160 ( // @[Stab.scala 175:24]
    .clock(last_merger_160_clock),
    .reset(last_merger_160_reset),
    .io_stream1_ready(last_merger_160_io_stream1_ready),
    .io_stream1_valid(last_merger_160_io_stream1_valid),
    .io_stream1_bits(last_merger_160_io_stream1_bits),
    .io_stream2_ready(last_merger_160_io_stream2_ready),
    .io_stream2_valid(last_merger_160_io_stream2_valid),
    .io_stream2_bits(last_merger_160_io_stream2_bits),
    .io_result_ready(last_merger_160_io_result_ready),
    .io_result_valid(last_merger_160_io_result_valid),
    .io_result_bits(last_merger_160_io_result_bits)
  );
  Queue last_q_160 ( // @[Decoupled.scala 361:21]
    .clock(last_q_160_clock),
    .reset(last_q_160_reset),
    .io_enq_ready(last_q_160_io_enq_ready),
    .io_enq_valid(last_q_160_io_enq_valid),
    .io_enq_bits(last_q_160_io_enq_bits),
    .io_deq_ready(last_q_160_io_deq_ready),
    .io_deq_valid(last_q_160_io_deq_valid),
    .io_deq_bits(last_q_160_io_deq_bits)
  );
  StreamMerger_161 last_merger_161 ( // @[Stab.scala 175:24]
    .clock(last_merger_161_clock),
    .reset(last_merger_161_reset),
    .io_stream1_ready(last_merger_161_io_stream1_ready),
    .io_stream1_valid(last_merger_161_io_stream1_valid),
    .io_stream1_bits(last_merger_161_io_stream1_bits),
    .io_stream2_ready(last_merger_161_io_stream2_ready),
    .io_stream2_valid(last_merger_161_io_stream2_valid),
    .io_stream2_bits(last_merger_161_io_stream2_bits),
    .io_result_ready(last_merger_161_io_result_ready),
    .io_result_valid(last_merger_161_io_result_valid),
    .io_result_bits(last_merger_161_io_result_bits)
  );
  Queue last_q_161 ( // @[Decoupled.scala 361:21]
    .clock(last_q_161_clock),
    .reset(last_q_161_reset),
    .io_enq_ready(last_q_161_io_enq_ready),
    .io_enq_valid(last_q_161_io_enq_valid),
    .io_enq_bits(last_q_161_io_enq_bits),
    .io_deq_ready(last_q_161_io_deq_ready),
    .io_deq_valid(last_q_161_io_deq_valid),
    .io_deq_bits(last_q_161_io_deq_bits)
  );
  StreamMerger_162 last_merger_162 ( // @[Stab.scala 175:24]
    .clock(last_merger_162_clock),
    .reset(last_merger_162_reset),
    .io_stream1_ready(last_merger_162_io_stream1_ready),
    .io_stream1_valid(last_merger_162_io_stream1_valid),
    .io_stream1_bits(last_merger_162_io_stream1_bits),
    .io_stream2_ready(last_merger_162_io_stream2_ready),
    .io_stream2_valid(last_merger_162_io_stream2_valid),
    .io_stream2_bits(last_merger_162_io_stream2_bits),
    .io_result_ready(last_merger_162_io_result_ready),
    .io_result_valid(last_merger_162_io_result_valid),
    .io_result_bits(last_merger_162_io_result_bits)
  );
  Queue last_q_162 ( // @[Decoupled.scala 361:21]
    .clock(last_q_162_clock),
    .reset(last_q_162_reset),
    .io_enq_ready(last_q_162_io_enq_ready),
    .io_enq_valid(last_q_162_io_enq_valid),
    .io_enq_bits(last_q_162_io_enq_bits),
    .io_deq_ready(last_q_162_io_deq_ready),
    .io_deq_valid(last_q_162_io_deq_valid),
    .io_deq_bits(last_q_162_io_deq_bits)
  );
  StreamMerger_163 last_merger_163 ( // @[Stab.scala 175:24]
    .clock(last_merger_163_clock),
    .reset(last_merger_163_reset),
    .io_stream1_ready(last_merger_163_io_stream1_ready),
    .io_stream1_valid(last_merger_163_io_stream1_valid),
    .io_stream1_bits(last_merger_163_io_stream1_bits),
    .io_stream2_ready(last_merger_163_io_stream2_ready),
    .io_stream2_valid(last_merger_163_io_stream2_valid),
    .io_stream2_bits(last_merger_163_io_stream2_bits),
    .io_result_ready(last_merger_163_io_result_ready),
    .io_result_valid(last_merger_163_io_result_valid),
    .io_result_bits(last_merger_163_io_result_bits)
  );
  Queue last_q_163 ( // @[Decoupled.scala 361:21]
    .clock(last_q_163_clock),
    .reset(last_q_163_reset),
    .io_enq_ready(last_q_163_io_enq_ready),
    .io_enq_valid(last_q_163_io_enq_valid),
    .io_enq_bits(last_q_163_io_enq_bits),
    .io_deq_ready(last_q_163_io_deq_ready),
    .io_deq_valid(last_q_163_io_deq_valid),
    .io_deq_bits(last_q_163_io_deq_bits)
  );
  StreamMerger_164 last_merger_164 ( // @[Stab.scala 175:24]
    .clock(last_merger_164_clock),
    .reset(last_merger_164_reset),
    .io_stream1_ready(last_merger_164_io_stream1_ready),
    .io_stream1_valid(last_merger_164_io_stream1_valid),
    .io_stream1_bits(last_merger_164_io_stream1_bits),
    .io_stream2_ready(last_merger_164_io_stream2_ready),
    .io_stream2_valid(last_merger_164_io_stream2_valid),
    .io_stream2_bits(last_merger_164_io_stream2_bits),
    .io_result_ready(last_merger_164_io_result_ready),
    .io_result_valid(last_merger_164_io_result_valid),
    .io_result_bits(last_merger_164_io_result_bits)
  );
  Queue last_q_164 ( // @[Decoupled.scala 361:21]
    .clock(last_q_164_clock),
    .reset(last_q_164_reset),
    .io_enq_ready(last_q_164_io_enq_ready),
    .io_enq_valid(last_q_164_io_enq_valid),
    .io_enq_bits(last_q_164_io_enq_bits),
    .io_deq_ready(last_q_164_io_deq_ready),
    .io_deq_valid(last_q_164_io_deq_valid),
    .io_deq_bits(last_q_164_io_deq_bits)
  );
  StreamMerger_165 last_merger_165 ( // @[Stab.scala 175:24]
    .clock(last_merger_165_clock),
    .reset(last_merger_165_reset),
    .io_stream1_ready(last_merger_165_io_stream1_ready),
    .io_stream1_valid(last_merger_165_io_stream1_valid),
    .io_stream1_bits(last_merger_165_io_stream1_bits),
    .io_stream2_ready(last_merger_165_io_stream2_ready),
    .io_stream2_valid(last_merger_165_io_stream2_valid),
    .io_stream2_bits(last_merger_165_io_stream2_bits),
    .io_result_ready(last_merger_165_io_result_ready),
    .io_result_valid(last_merger_165_io_result_valid),
    .io_result_bits(last_merger_165_io_result_bits)
  );
  Queue last_q_165 ( // @[Decoupled.scala 361:21]
    .clock(last_q_165_clock),
    .reset(last_q_165_reset),
    .io_enq_ready(last_q_165_io_enq_ready),
    .io_enq_valid(last_q_165_io_enq_valid),
    .io_enq_bits(last_q_165_io_enq_bits),
    .io_deq_ready(last_q_165_io_deq_ready),
    .io_deq_valid(last_q_165_io_deq_valid),
    .io_deq_bits(last_q_165_io_deq_bits)
  );
  StreamMerger_166 last_merger_166 ( // @[Stab.scala 175:24]
    .clock(last_merger_166_clock),
    .reset(last_merger_166_reset),
    .io_stream1_ready(last_merger_166_io_stream1_ready),
    .io_stream1_valid(last_merger_166_io_stream1_valid),
    .io_stream1_bits(last_merger_166_io_stream1_bits),
    .io_stream2_ready(last_merger_166_io_stream2_ready),
    .io_stream2_valid(last_merger_166_io_stream2_valid),
    .io_stream2_bits(last_merger_166_io_stream2_bits),
    .io_result_ready(last_merger_166_io_result_ready),
    .io_result_valid(last_merger_166_io_result_valid),
    .io_result_bits(last_merger_166_io_result_bits)
  );
  Queue last_q_166 ( // @[Decoupled.scala 361:21]
    .clock(last_q_166_clock),
    .reset(last_q_166_reset),
    .io_enq_ready(last_q_166_io_enq_ready),
    .io_enq_valid(last_q_166_io_enq_valid),
    .io_enq_bits(last_q_166_io_enq_bits),
    .io_deq_ready(last_q_166_io_deq_ready),
    .io_deq_valid(last_q_166_io_deq_valid),
    .io_deq_bits(last_q_166_io_deq_bits)
  );
  StreamMerger_167 last_merger_167 ( // @[Stab.scala 175:24]
    .clock(last_merger_167_clock),
    .reset(last_merger_167_reset),
    .io_stream1_ready(last_merger_167_io_stream1_ready),
    .io_stream1_valid(last_merger_167_io_stream1_valid),
    .io_stream1_bits(last_merger_167_io_stream1_bits),
    .io_stream2_ready(last_merger_167_io_stream2_ready),
    .io_stream2_valid(last_merger_167_io_stream2_valid),
    .io_stream2_bits(last_merger_167_io_stream2_bits),
    .io_result_ready(last_merger_167_io_result_ready),
    .io_result_valid(last_merger_167_io_result_valid),
    .io_result_bits(last_merger_167_io_result_bits)
  );
  Queue last_q_167 ( // @[Decoupled.scala 361:21]
    .clock(last_q_167_clock),
    .reset(last_q_167_reset),
    .io_enq_ready(last_q_167_io_enq_ready),
    .io_enq_valid(last_q_167_io_enq_valid),
    .io_enq_bits(last_q_167_io_enq_bits),
    .io_deq_ready(last_q_167_io_deq_ready),
    .io_deq_valid(last_q_167_io_deq_valid),
    .io_deq_bits(last_q_167_io_deq_bits)
  );
  StreamMerger_168 last_merger_168 ( // @[Stab.scala 175:24]
    .clock(last_merger_168_clock),
    .reset(last_merger_168_reset),
    .io_stream1_ready(last_merger_168_io_stream1_ready),
    .io_stream1_valid(last_merger_168_io_stream1_valid),
    .io_stream1_bits(last_merger_168_io_stream1_bits),
    .io_stream2_ready(last_merger_168_io_stream2_ready),
    .io_stream2_valid(last_merger_168_io_stream2_valid),
    .io_stream2_bits(last_merger_168_io_stream2_bits),
    .io_result_ready(last_merger_168_io_result_ready),
    .io_result_valid(last_merger_168_io_result_valid),
    .io_result_bits(last_merger_168_io_result_bits)
  );
  Queue last_q_168 ( // @[Decoupled.scala 361:21]
    .clock(last_q_168_clock),
    .reset(last_q_168_reset),
    .io_enq_ready(last_q_168_io_enq_ready),
    .io_enq_valid(last_q_168_io_enq_valid),
    .io_enq_bits(last_q_168_io_enq_bits),
    .io_deq_ready(last_q_168_io_deq_ready),
    .io_deq_valid(last_q_168_io_deq_valid),
    .io_deq_bits(last_q_168_io_deq_bits)
  );
  StreamMerger_169 last_merger_169 ( // @[Stab.scala 175:24]
    .clock(last_merger_169_clock),
    .reset(last_merger_169_reset),
    .io_stream1_ready(last_merger_169_io_stream1_ready),
    .io_stream1_valid(last_merger_169_io_stream1_valid),
    .io_stream1_bits(last_merger_169_io_stream1_bits),
    .io_stream2_ready(last_merger_169_io_stream2_ready),
    .io_stream2_valid(last_merger_169_io_stream2_valid),
    .io_stream2_bits(last_merger_169_io_stream2_bits),
    .io_result_ready(last_merger_169_io_result_ready),
    .io_result_valid(last_merger_169_io_result_valid),
    .io_result_bits(last_merger_169_io_result_bits)
  );
  Queue last_q_169 ( // @[Decoupled.scala 361:21]
    .clock(last_q_169_clock),
    .reset(last_q_169_reset),
    .io_enq_ready(last_q_169_io_enq_ready),
    .io_enq_valid(last_q_169_io_enq_valid),
    .io_enq_bits(last_q_169_io_enq_bits),
    .io_deq_ready(last_q_169_io_deq_ready),
    .io_deq_valid(last_q_169_io_deq_valid),
    .io_deq_bits(last_q_169_io_deq_bits)
  );
  StreamMerger_170 last_merger_170 ( // @[Stab.scala 175:24]
    .clock(last_merger_170_clock),
    .reset(last_merger_170_reset),
    .io_stream1_ready(last_merger_170_io_stream1_ready),
    .io_stream1_valid(last_merger_170_io_stream1_valid),
    .io_stream1_bits(last_merger_170_io_stream1_bits),
    .io_stream2_ready(last_merger_170_io_stream2_ready),
    .io_stream2_valid(last_merger_170_io_stream2_valid),
    .io_stream2_bits(last_merger_170_io_stream2_bits),
    .io_result_ready(last_merger_170_io_result_ready),
    .io_result_valid(last_merger_170_io_result_valid),
    .io_result_bits(last_merger_170_io_result_bits)
  );
  Queue last_q_170 ( // @[Decoupled.scala 361:21]
    .clock(last_q_170_clock),
    .reset(last_q_170_reset),
    .io_enq_ready(last_q_170_io_enq_ready),
    .io_enq_valid(last_q_170_io_enq_valid),
    .io_enq_bits(last_q_170_io_enq_bits),
    .io_deq_ready(last_q_170_io_deq_ready),
    .io_deq_valid(last_q_170_io_deq_valid),
    .io_deq_bits(last_q_170_io_deq_bits)
  );
  StreamMerger_171 last_merger_171 ( // @[Stab.scala 175:24]
    .clock(last_merger_171_clock),
    .reset(last_merger_171_reset),
    .io_stream1_ready(last_merger_171_io_stream1_ready),
    .io_stream1_valid(last_merger_171_io_stream1_valid),
    .io_stream1_bits(last_merger_171_io_stream1_bits),
    .io_stream2_ready(last_merger_171_io_stream2_ready),
    .io_stream2_valid(last_merger_171_io_stream2_valid),
    .io_stream2_bits(last_merger_171_io_stream2_bits),
    .io_result_ready(last_merger_171_io_result_ready),
    .io_result_valid(last_merger_171_io_result_valid),
    .io_result_bits(last_merger_171_io_result_bits)
  );
  Queue last_q_171 ( // @[Decoupled.scala 361:21]
    .clock(last_q_171_clock),
    .reset(last_q_171_reset),
    .io_enq_ready(last_q_171_io_enq_ready),
    .io_enq_valid(last_q_171_io_enq_valid),
    .io_enq_bits(last_q_171_io_enq_bits),
    .io_deq_ready(last_q_171_io_deq_ready),
    .io_deq_valid(last_q_171_io_deq_valid),
    .io_deq_bits(last_q_171_io_deq_bits)
  );
  StreamMerger_172 last_merger_172 ( // @[Stab.scala 175:24]
    .clock(last_merger_172_clock),
    .reset(last_merger_172_reset),
    .io_stream1_ready(last_merger_172_io_stream1_ready),
    .io_stream1_valid(last_merger_172_io_stream1_valid),
    .io_stream1_bits(last_merger_172_io_stream1_bits),
    .io_stream2_ready(last_merger_172_io_stream2_ready),
    .io_stream2_valid(last_merger_172_io_stream2_valid),
    .io_stream2_bits(last_merger_172_io_stream2_bits),
    .io_result_ready(last_merger_172_io_result_ready),
    .io_result_valid(last_merger_172_io_result_valid),
    .io_result_bits(last_merger_172_io_result_bits)
  );
  Queue last_q_172 ( // @[Decoupled.scala 361:21]
    .clock(last_q_172_clock),
    .reset(last_q_172_reset),
    .io_enq_ready(last_q_172_io_enq_ready),
    .io_enq_valid(last_q_172_io_enq_valid),
    .io_enq_bits(last_q_172_io_enq_bits),
    .io_deq_ready(last_q_172_io_deq_ready),
    .io_deq_valid(last_q_172_io_deq_valid),
    .io_deq_bits(last_q_172_io_deq_bits)
  );
  StreamMerger_173 last_merger_173 ( // @[Stab.scala 175:24]
    .clock(last_merger_173_clock),
    .reset(last_merger_173_reset),
    .io_stream1_ready(last_merger_173_io_stream1_ready),
    .io_stream1_valid(last_merger_173_io_stream1_valid),
    .io_stream1_bits(last_merger_173_io_stream1_bits),
    .io_stream2_ready(last_merger_173_io_stream2_ready),
    .io_stream2_valid(last_merger_173_io_stream2_valid),
    .io_stream2_bits(last_merger_173_io_stream2_bits),
    .io_result_ready(last_merger_173_io_result_ready),
    .io_result_valid(last_merger_173_io_result_valid),
    .io_result_bits(last_merger_173_io_result_bits)
  );
  Queue last_q_173 ( // @[Decoupled.scala 361:21]
    .clock(last_q_173_clock),
    .reset(last_q_173_reset),
    .io_enq_ready(last_q_173_io_enq_ready),
    .io_enq_valid(last_q_173_io_enq_valid),
    .io_enq_bits(last_q_173_io_enq_bits),
    .io_deq_ready(last_q_173_io_deq_ready),
    .io_deq_valid(last_q_173_io_deq_valid),
    .io_deq_bits(last_q_173_io_deq_bits)
  );
  StreamMerger_174 last_merger_174 ( // @[Stab.scala 175:24]
    .clock(last_merger_174_clock),
    .reset(last_merger_174_reset),
    .io_stream1_ready(last_merger_174_io_stream1_ready),
    .io_stream1_valid(last_merger_174_io_stream1_valid),
    .io_stream1_bits(last_merger_174_io_stream1_bits),
    .io_stream2_ready(last_merger_174_io_stream2_ready),
    .io_stream2_valid(last_merger_174_io_stream2_valid),
    .io_stream2_bits(last_merger_174_io_stream2_bits),
    .io_result_ready(last_merger_174_io_result_ready),
    .io_result_valid(last_merger_174_io_result_valid),
    .io_result_bits(last_merger_174_io_result_bits)
  );
  Queue last_q_174 ( // @[Decoupled.scala 361:21]
    .clock(last_q_174_clock),
    .reset(last_q_174_reset),
    .io_enq_ready(last_q_174_io_enq_ready),
    .io_enq_valid(last_q_174_io_enq_valid),
    .io_enq_bits(last_q_174_io_enq_bits),
    .io_deq_ready(last_q_174_io_deq_ready),
    .io_deq_valid(last_q_174_io_deq_valid),
    .io_deq_bits(last_q_174_io_deq_bits)
  );
  StreamMerger_175 last_merger_175 ( // @[Stab.scala 175:24]
    .clock(last_merger_175_clock),
    .reset(last_merger_175_reset),
    .io_stream1_ready(last_merger_175_io_stream1_ready),
    .io_stream1_valid(last_merger_175_io_stream1_valid),
    .io_stream1_bits(last_merger_175_io_stream1_bits),
    .io_stream2_ready(last_merger_175_io_stream2_ready),
    .io_stream2_valid(last_merger_175_io_stream2_valid),
    .io_stream2_bits(last_merger_175_io_stream2_bits),
    .io_result_ready(last_merger_175_io_result_ready),
    .io_result_valid(last_merger_175_io_result_valid),
    .io_result_bits(last_merger_175_io_result_bits)
  );
  Queue last_q_175 ( // @[Decoupled.scala 361:21]
    .clock(last_q_175_clock),
    .reset(last_q_175_reset),
    .io_enq_ready(last_q_175_io_enq_ready),
    .io_enq_valid(last_q_175_io_enq_valid),
    .io_enq_bits(last_q_175_io_enq_bits),
    .io_deq_ready(last_q_175_io_deq_ready),
    .io_deq_valid(last_q_175_io_deq_valid),
    .io_deq_bits(last_q_175_io_deq_bits)
  );
  StreamMerger_176 last_merger_176 ( // @[Stab.scala 175:24]
    .clock(last_merger_176_clock),
    .reset(last_merger_176_reset),
    .io_stream1_ready(last_merger_176_io_stream1_ready),
    .io_stream1_valid(last_merger_176_io_stream1_valid),
    .io_stream1_bits(last_merger_176_io_stream1_bits),
    .io_stream2_ready(last_merger_176_io_stream2_ready),
    .io_stream2_valid(last_merger_176_io_stream2_valid),
    .io_stream2_bits(last_merger_176_io_stream2_bits),
    .io_result_ready(last_merger_176_io_result_ready),
    .io_result_valid(last_merger_176_io_result_valid),
    .io_result_bits(last_merger_176_io_result_bits)
  );
  Queue last_q_176 ( // @[Decoupled.scala 361:21]
    .clock(last_q_176_clock),
    .reset(last_q_176_reset),
    .io_enq_ready(last_q_176_io_enq_ready),
    .io_enq_valid(last_q_176_io_enq_valid),
    .io_enq_bits(last_q_176_io_enq_bits),
    .io_deq_ready(last_q_176_io_deq_ready),
    .io_deq_valid(last_q_176_io_deq_valid),
    .io_deq_bits(last_q_176_io_deq_bits)
  );
  StreamMerger_177 last_merger_177 ( // @[Stab.scala 175:24]
    .clock(last_merger_177_clock),
    .reset(last_merger_177_reset),
    .io_stream1_ready(last_merger_177_io_stream1_ready),
    .io_stream1_valid(last_merger_177_io_stream1_valid),
    .io_stream1_bits(last_merger_177_io_stream1_bits),
    .io_stream2_ready(last_merger_177_io_stream2_ready),
    .io_stream2_valid(last_merger_177_io_stream2_valid),
    .io_stream2_bits(last_merger_177_io_stream2_bits),
    .io_result_ready(last_merger_177_io_result_ready),
    .io_result_valid(last_merger_177_io_result_valid),
    .io_result_bits(last_merger_177_io_result_bits)
  );
  Queue last_q_177 ( // @[Decoupled.scala 361:21]
    .clock(last_q_177_clock),
    .reset(last_q_177_reset),
    .io_enq_ready(last_q_177_io_enq_ready),
    .io_enq_valid(last_q_177_io_enq_valid),
    .io_enq_bits(last_q_177_io_enq_bits),
    .io_deq_ready(last_q_177_io_deq_ready),
    .io_deq_valid(last_q_177_io_deq_valid),
    .io_deq_bits(last_q_177_io_deq_bits)
  );
  StreamMerger_178 last_merger_178 ( // @[Stab.scala 175:24]
    .clock(last_merger_178_clock),
    .reset(last_merger_178_reset),
    .io_stream1_ready(last_merger_178_io_stream1_ready),
    .io_stream1_valid(last_merger_178_io_stream1_valid),
    .io_stream1_bits(last_merger_178_io_stream1_bits),
    .io_stream2_ready(last_merger_178_io_stream2_ready),
    .io_stream2_valid(last_merger_178_io_stream2_valid),
    .io_stream2_bits(last_merger_178_io_stream2_bits),
    .io_result_ready(last_merger_178_io_result_ready),
    .io_result_valid(last_merger_178_io_result_valid),
    .io_result_bits(last_merger_178_io_result_bits)
  );
  Queue last_q_178 ( // @[Decoupled.scala 361:21]
    .clock(last_q_178_clock),
    .reset(last_q_178_reset),
    .io_enq_ready(last_q_178_io_enq_ready),
    .io_enq_valid(last_q_178_io_enq_valid),
    .io_enq_bits(last_q_178_io_enq_bits),
    .io_deq_ready(last_q_178_io_deq_ready),
    .io_deq_valid(last_q_178_io_deq_valid),
    .io_deq_bits(last_q_178_io_deq_bits)
  );
  StreamMerger_179 last_merger_179 ( // @[Stab.scala 175:24]
    .clock(last_merger_179_clock),
    .reset(last_merger_179_reset),
    .io_stream1_ready(last_merger_179_io_stream1_ready),
    .io_stream1_valid(last_merger_179_io_stream1_valid),
    .io_stream1_bits(last_merger_179_io_stream1_bits),
    .io_stream2_ready(last_merger_179_io_stream2_ready),
    .io_stream2_valid(last_merger_179_io_stream2_valid),
    .io_stream2_bits(last_merger_179_io_stream2_bits),
    .io_result_ready(last_merger_179_io_result_ready),
    .io_result_valid(last_merger_179_io_result_valid),
    .io_result_bits(last_merger_179_io_result_bits)
  );
  Queue last_q_179 ( // @[Decoupled.scala 361:21]
    .clock(last_q_179_clock),
    .reset(last_q_179_reset),
    .io_enq_ready(last_q_179_io_enq_ready),
    .io_enq_valid(last_q_179_io_enq_valid),
    .io_enq_bits(last_q_179_io_enq_bits),
    .io_deq_ready(last_q_179_io_deq_ready),
    .io_deq_valid(last_q_179_io_deq_valid),
    .io_deq_bits(last_q_179_io_deq_bits)
  );
  StreamMerger_180 last_merger_180 ( // @[Stab.scala 175:24]
    .clock(last_merger_180_clock),
    .reset(last_merger_180_reset),
    .io_stream1_ready(last_merger_180_io_stream1_ready),
    .io_stream1_valid(last_merger_180_io_stream1_valid),
    .io_stream1_bits(last_merger_180_io_stream1_bits),
    .io_stream2_ready(last_merger_180_io_stream2_ready),
    .io_stream2_valid(last_merger_180_io_stream2_valid),
    .io_stream2_bits(last_merger_180_io_stream2_bits),
    .io_result_ready(last_merger_180_io_result_ready),
    .io_result_valid(last_merger_180_io_result_valid),
    .io_result_bits(last_merger_180_io_result_bits)
  );
  Queue last_q_180 ( // @[Decoupled.scala 361:21]
    .clock(last_q_180_clock),
    .reset(last_q_180_reset),
    .io_enq_ready(last_q_180_io_enq_ready),
    .io_enq_valid(last_q_180_io_enq_valid),
    .io_enq_bits(last_q_180_io_enq_bits),
    .io_deq_ready(last_q_180_io_deq_ready),
    .io_deq_valid(last_q_180_io_deq_valid),
    .io_deq_bits(last_q_180_io_deq_bits)
  );
  StreamMerger_181 last_merger_181 ( // @[Stab.scala 175:24]
    .clock(last_merger_181_clock),
    .reset(last_merger_181_reset),
    .io_stream1_ready(last_merger_181_io_stream1_ready),
    .io_stream1_valid(last_merger_181_io_stream1_valid),
    .io_stream1_bits(last_merger_181_io_stream1_bits),
    .io_stream2_ready(last_merger_181_io_stream2_ready),
    .io_stream2_valid(last_merger_181_io_stream2_valid),
    .io_stream2_bits(last_merger_181_io_stream2_bits),
    .io_result_ready(last_merger_181_io_result_ready),
    .io_result_valid(last_merger_181_io_result_valid),
    .io_result_bits(last_merger_181_io_result_bits)
  );
  Queue last_q_181 ( // @[Decoupled.scala 361:21]
    .clock(last_q_181_clock),
    .reset(last_q_181_reset),
    .io_enq_ready(last_q_181_io_enq_ready),
    .io_enq_valid(last_q_181_io_enq_valid),
    .io_enq_bits(last_q_181_io_enq_bits),
    .io_deq_ready(last_q_181_io_deq_ready),
    .io_deq_valid(last_q_181_io_deq_valid),
    .io_deq_bits(last_q_181_io_deq_bits)
  );
  StreamMerger_182 last_merger_182 ( // @[Stab.scala 175:24]
    .clock(last_merger_182_clock),
    .reset(last_merger_182_reset),
    .io_stream1_ready(last_merger_182_io_stream1_ready),
    .io_stream1_valid(last_merger_182_io_stream1_valid),
    .io_stream1_bits(last_merger_182_io_stream1_bits),
    .io_stream2_ready(last_merger_182_io_stream2_ready),
    .io_stream2_valid(last_merger_182_io_stream2_valid),
    .io_stream2_bits(last_merger_182_io_stream2_bits),
    .io_result_ready(last_merger_182_io_result_ready),
    .io_result_valid(last_merger_182_io_result_valid),
    .io_result_bits(last_merger_182_io_result_bits)
  );
  Queue last_q_182 ( // @[Decoupled.scala 361:21]
    .clock(last_q_182_clock),
    .reset(last_q_182_reset),
    .io_enq_ready(last_q_182_io_enq_ready),
    .io_enq_valid(last_q_182_io_enq_valid),
    .io_enq_bits(last_q_182_io_enq_bits),
    .io_deq_ready(last_q_182_io_deq_ready),
    .io_deq_valid(last_q_182_io_deq_valid),
    .io_deq_bits(last_q_182_io_deq_bits)
  );
  StreamMerger_183 last_merger_183 ( // @[Stab.scala 175:24]
    .clock(last_merger_183_clock),
    .reset(last_merger_183_reset),
    .io_stream1_ready(last_merger_183_io_stream1_ready),
    .io_stream1_valid(last_merger_183_io_stream1_valid),
    .io_stream1_bits(last_merger_183_io_stream1_bits),
    .io_stream2_ready(last_merger_183_io_stream2_ready),
    .io_stream2_valid(last_merger_183_io_stream2_valid),
    .io_stream2_bits(last_merger_183_io_stream2_bits),
    .io_result_ready(last_merger_183_io_result_ready),
    .io_result_valid(last_merger_183_io_result_valid),
    .io_result_bits(last_merger_183_io_result_bits)
  );
  Queue last_q_183 ( // @[Decoupled.scala 361:21]
    .clock(last_q_183_clock),
    .reset(last_q_183_reset),
    .io_enq_ready(last_q_183_io_enq_ready),
    .io_enq_valid(last_q_183_io_enq_valid),
    .io_enq_bits(last_q_183_io_enq_bits),
    .io_deq_ready(last_q_183_io_deq_ready),
    .io_deq_valid(last_q_183_io_deq_valid),
    .io_deq_bits(last_q_183_io_deq_bits)
  );
  StreamMerger_184 last_merger_184 ( // @[Stab.scala 175:24]
    .clock(last_merger_184_clock),
    .reset(last_merger_184_reset),
    .io_stream1_ready(last_merger_184_io_stream1_ready),
    .io_stream1_valid(last_merger_184_io_stream1_valid),
    .io_stream1_bits(last_merger_184_io_stream1_bits),
    .io_stream2_ready(last_merger_184_io_stream2_ready),
    .io_stream2_valid(last_merger_184_io_stream2_valid),
    .io_stream2_bits(last_merger_184_io_stream2_bits),
    .io_result_ready(last_merger_184_io_result_ready),
    .io_result_valid(last_merger_184_io_result_valid),
    .io_result_bits(last_merger_184_io_result_bits)
  );
  Queue last_q_184 ( // @[Decoupled.scala 361:21]
    .clock(last_q_184_clock),
    .reset(last_q_184_reset),
    .io_enq_ready(last_q_184_io_enq_ready),
    .io_enq_valid(last_q_184_io_enq_valid),
    .io_enq_bits(last_q_184_io_enq_bits),
    .io_deq_ready(last_q_184_io_deq_ready),
    .io_deq_valid(last_q_184_io_deq_valid),
    .io_deq_bits(last_q_184_io_deq_bits)
  );
  StreamMerger_185 last_merger_185 ( // @[Stab.scala 175:24]
    .clock(last_merger_185_clock),
    .reset(last_merger_185_reset),
    .io_stream1_ready(last_merger_185_io_stream1_ready),
    .io_stream1_valid(last_merger_185_io_stream1_valid),
    .io_stream1_bits(last_merger_185_io_stream1_bits),
    .io_stream2_ready(last_merger_185_io_stream2_ready),
    .io_stream2_valid(last_merger_185_io_stream2_valid),
    .io_stream2_bits(last_merger_185_io_stream2_bits),
    .io_result_ready(last_merger_185_io_result_ready),
    .io_result_valid(last_merger_185_io_result_valid),
    .io_result_bits(last_merger_185_io_result_bits)
  );
  Queue last_q_185 ( // @[Decoupled.scala 361:21]
    .clock(last_q_185_clock),
    .reset(last_q_185_reset),
    .io_enq_ready(last_q_185_io_enq_ready),
    .io_enq_valid(last_q_185_io_enq_valid),
    .io_enq_bits(last_q_185_io_enq_bits),
    .io_deq_ready(last_q_185_io_deq_ready),
    .io_deq_valid(last_q_185_io_deq_valid),
    .io_deq_bits(last_q_185_io_deq_bits)
  );
  StreamMerger_186 last_merger_186 ( // @[Stab.scala 175:24]
    .clock(last_merger_186_clock),
    .reset(last_merger_186_reset),
    .io_stream1_ready(last_merger_186_io_stream1_ready),
    .io_stream1_valid(last_merger_186_io_stream1_valid),
    .io_stream1_bits(last_merger_186_io_stream1_bits),
    .io_stream2_ready(last_merger_186_io_stream2_ready),
    .io_stream2_valid(last_merger_186_io_stream2_valid),
    .io_stream2_bits(last_merger_186_io_stream2_bits),
    .io_result_ready(last_merger_186_io_result_ready),
    .io_result_valid(last_merger_186_io_result_valid),
    .io_result_bits(last_merger_186_io_result_bits)
  );
  Queue last_q_186 ( // @[Decoupled.scala 361:21]
    .clock(last_q_186_clock),
    .reset(last_q_186_reset),
    .io_enq_ready(last_q_186_io_enq_ready),
    .io_enq_valid(last_q_186_io_enq_valid),
    .io_enq_bits(last_q_186_io_enq_bits),
    .io_deq_ready(last_q_186_io_deq_ready),
    .io_deq_valid(last_q_186_io_deq_valid),
    .io_deq_bits(last_q_186_io_deq_bits)
  );
  StreamMerger_187 last_merger_187 ( // @[Stab.scala 175:24]
    .clock(last_merger_187_clock),
    .reset(last_merger_187_reset),
    .io_stream1_ready(last_merger_187_io_stream1_ready),
    .io_stream1_valid(last_merger_187_io_stream1_valid),
    .io_stream1_bits(last_merger_187_io_stream1_bits),
    .io_stream2_ready(last_merger_187_io_stream2_ready),
    .io_stream2_valid(last_merger_187_io_stream2_valid),
    .io_stream2_bits(last_merger_187_io_stream2_bits),
    .io_result_ready(last_merger_187_io_result_ready),
    .io_result_valid(last_merger_187_io_result_valid),
    .io_result_bits(last_merger_187_io_result_bits)
  );
  Queue last_q_187 ( // @[Decoupled.scala 361:21]
    .clock(last_q_187_clock),
    .reset(last_q_187_reset),
    .io_enq_ready(last_q_187_io_enq_ready),
    .io_enq_valid(last_q_187_io_enq_valid),
    .io_enq_bits(last_q_187_io_enq_bits),
    .io_deq_ready(last_q_187_io_deq_ready),
    .io_deq_valid(last_q_187_io_deq_valid),
    .io_deq_bits(last_q_187_io_deq_bits)
  );
  StreamMerger_188 last_merger_188 ( // @[Stab.scala 175:24]
    .clock(last_merger_188_clock),
    .reset(last_merger_188_reset),
    .io_stream1_ready(last_merger_188_io_stream1_ready),
    .io_stream1_valid(last_merger_188_io_stream1_valid),
    .io_stream1_bits(last_merger_188_io_stream1_bits),
    .io_stream2_ready(last_merger_188_io_stream2_ready),
    .io_stream2_valid(last_merger_188_io_stream2_valid),
    .io_stream2_bits(last_merger_188_io_stream2_bits),
    .io_result_ready(last_merger_188_io_result_ready),
    .io_result_valid(last_merger_188_io_result_valid),
    .io_result_bits(last_merger_188_io_result_bits)
  );
  Queue last_q_188 ( // @[Decoupled.scala 361:21]
    .clock(last_q_188_clock),
    .reset(last_q_188_reset),
    .io_enq_ready(last_q_188_io_enq_ready),
    .io_enq_valid(last_q_188_io_enq_valid),
    .io_enq_bits(last_q_188_io_enq_bits),
    .io_deq_ready(last_q_188_io_deq_ready),
    .io_deq_valid(last_q_188_io_deq_valid),
    .io_deq_bits(last_q_188_io_deq_bits)
  );
  StreamMerger_189 last_merger_189 ( // @[Stab.scala 175:24]
    .clock(last_merger_189_clock),
    .reset(last_merger_189_reset),
    .io_stream1_ready(last_merger_189_io_stream1_ready),
    .io_stream1_valid(last_merger_189_io_stream1_valid),
    .io_stream1_bits(last_merger_189_io_stream1_bits),
    .io_stream2_ready(last_merger_189_io_stream2_ready),
    .io_stream2_valid(last_merger_189_io_stream2_valid),
    .io_stream2_bits(last_merger_189_io_stream2_bits),
    .io_result_ready(last_merger_189_io_result_ready),
    .io_result_valid(last_merger_189_io_result_valid),
    .io_result_bits(last_merger_189_io_result_bits)
  );
  Queue last_q_189 ( // @[Decoupled.scala 361:21]
    .clock(last_q_189_clock),
    .reset(last_q_189_reset),
    .io_enq_ready(last_q_189_io_enq_ready),
    .io_enq_valid(last_q_189_io_enq_valid),
    .io_enq_bits(last_q_189_io_enq_bits),
    .io_deq_ready(last_q_189_io_deq_ready),
    .io_deq_valid(last_q_189_io_deq_valid),
    .io_deq_bits(last_q_189_io_deq_bits)
  );
  StreamMerger_190 last_merger_190 ( // @[Stab.scala 175:24]
    .clock(last_merger_190_clock),
    .reset(last_merger_190_reset),
    .io_stream1_ready(last_merger_190_io_stream1_ready),
    .io_stream1_valid(last_merger_190_io_stream1_valid),
    .io_stream1_bits(last_merger_190_io_stream1_bits),
    .io_stream2_ready(last_merger_190_io_stream2_ready),
    .io_stream2_valid(last_merger_190_io_stream2_valid),
    .io_stream2_bits(last_merger_190_io_stream2_bits),
    .io_result_ready(last_merger_190_io_result_ready),
    .io_result_valid(last_merger_190_io_result_valid),
    .io_result_bits(last_merger_190_io_result_bits)
  );
  Queue last_q_190 ( // @[Decoupled.scala 361:21]
    .clock(last_q_190_clock),
    .reset(last_q_190_reset),
    .io_enq_ready(last_q_190_io_enq_ready),
    .io_enq_valid(last_q_190_io_enq_valid),
    .io_enq_bits(last_q_190_io_enq_bits),
    .io_deq_ready(last_q_190_io_deq_ready),
    .io_deq_valid(last_q_190_io_deq_valid),
    .io_deq_bits(last_q_190_io_deq_bits)
  );
  StreamMerger_191 last_merger_191 ( // @[Stab.scala 175:24]
    .clock(last_merger_191_clock),
    .reset(last_merger_191_reset),
    .io_stream1_ready(last_merger_191_io_stream1_ready),
    .io_stream1_valid(last_merger_191_io_stream1_valid),
    .io_stream1_bits(last_merger_191_io_stream1_bits),
    .io_stream2_ready(last_merger_191_io_stream2_ready),
    .io_stream2_valid(last_merger_191_io_stream2_valid),
    .io_stream2_bits(last_merger_191_io_stream2_bits),
    .io_result_ready(last_merger_191_io_result_ready),
    .io_result_valid(last_merger_191_io_result_valid),
    .io_result_bits(last_merger_191_io_result_bits)
  );
  Queue last_q_191 ( // @[Decoupled.scala 361:21]
    .clock(last_q_191_clock),
    .reset(last_q_191_reset),
    .io_enq_ready(last_q_191_io_enq_ready),
    .io_enq_valid(last_q_191_io_enq_valid),
    .io_enq_bits(last_q_191_io_enq_bits),
    .io_deq_ready(last_q_191_io_deq_ready),
    .io_deq_valid(last_q_191_io_deq_valid),
    .io_deq_bits(last_q_191_io_deq_bits)
  );
  StreamMerger_192 last_merger_192 ( // @[Stab.scala 175:24]
    .clock(last_merger_192_clock),
    .reset(last_merger_192_reset),
    .io_stream1_ready(last_merger_192_io_stream1_ready),
    .io_stream1_valid(last_merger_192_io_stream1_valid),
    .io_stream1_bits(last_merger_192_io_stream1_bits),
    .io_stream2_ready(last_merger_192_io_stream2_ready),
    .io_stream2_valid(last_merger_192_io_stream2_valid),
    .io_stream2_bits(last_merger_192_io_stream2_bits),
    .io_result_ready(last_merger_192_io_result_ready),
    .io_result_valid(last_merger_192_io_result_valid),
    .io_result_bits(last_merger_192_io_result_bits)
  );
  Queue last_q_192 ( // @[Decoupled.scala 361:21]
    .clock(last_q_192_clock),
    .reset(last_q_192_reset),
    .io_enq_ready(last_q_192_io_enq_ready),
    .io_enq_valid(last_q_192_io_enq_valid),
    .io_enq_bits(last_q_192_io_enq_bits),
    .io_deq_ready(last_q_192_io_deq_ready),
    .io_deq_valid(last_q_192_io_deq_valid),
    .io_deq_bits(last_q_192_io_deq_bits)
  );
  StreamMerger_193 last_merger_193 ( // @[Stab.scala 175:24]
    .clock(last_merger_193_clock),
    .reset(last_merger_193_reset),
    .io_stream1_ready(last_merger_193_io_stream1_ready),
    .io_stream1_valid(last_merger_193_io_stream1_valid),
    .io_stream1_bits(last_merger_193_io_stream1_bits),
    .io_stream2_ready(last_merger_193_io_stream2_ready),
    .io_stream2_valid(last_merger_193_io_stream2_valid),
    .io_stream2_bits(last_merger_193_io_stream2_bits),
    .io_result_ready(last_merger_193_io_result_ready),
    .io_result_valid(last_merger_193_io_result_valid),
    .io_result_bits(last_merger_193_io_result_bits)
  );
  Queue last_q_193 ( // @[Decoupled.scala 361:21]
    .clock(last_q_193_clock),
    .reset(last_q_193_reset),
    .io_enq_ready(last_q_193_io_enq_ready),
    .io_enq_valid(last_q_193_io_enq_valid),
    .io_enq_bits(last_q_193_io_enq_bits),
    .io_deq_ready(last_q_193_io_deq_ready),
    .io_deq_valid(last_q_193_io_deq_valid),
    .io_deq_bits(last_q_193_io_deq_bits)
  );
  StreamMerger_194 last_merger_194 ( // @[Stab.scala 175:24]
    .clock(last_merger_194_clock),
    .reset(last_merger_194_reset),
    .io_stream1_ready(last_merger_194_io_stream1_ready),
    .io_stream1_valid(last_merger_194_io_stream1_valid),
    .io_stream1_bits(last_merger_194_io_stream1_bits),
    .io_stream2_ready(last_merger_194_io_stream2_ready),
    .io_stream2_valid(last_merger_194_io_stream2_valid),
    .io_stream2_bits(last_merger_194_io_stream2_bits),
    .io_result_ready(last_merger_194_io_result_ready),
    .io_result_valid(last_merger_194_io_result_valid),
    .io_result_bits(last_merger_194_io_result_bits)
  );
  Queue last_q_194 ( // @[Decoupled.scala 361:21]
    .clock(last_q_194_clock),
    .reset(last_q_194_reset),
    .io_enq_ready(last_q_194_io_enq_ready),
    .io_enq_valid(last_q_194_io_enq_valid),
    .io_enq_bits(last_q_194_io_enq_bits),
    .io_deq_ready(last_q_194_io_deq_ready),
    .io_deq_valid(last_q_194_io_deq_valid),
    .io_deq_bits(last_q_194_io_deq_bits)
  );
  StreamMerger_195 last_merger_195 ( // @[Stab.scala 175:24]
    .clock(last_merger_195_clock),
    .reset(last_merger_195_reset),
    .io_stream1_ready(last_merger_195_io_stream1_ready),
    .io_stream1_valid(last_merger_195_io_stream1_valid),
    .io_stream1_bits(last_merger_195_io_stream1_bits),
    .io_stream2_ready(last_merger_195_io_stream2_ready),
    .io_stream2_valid(last_merger_195_io_stream2_valid),
    .io_stream2_bits(last_merger_195_io_stream2_bits),
    .io_result_ready(last_merger_195_io_result_ready),
    .io_result_valid(last_merger_195_io_result_valid),
    .io_result_bits(last_merger_195_io_result_bits)
  );
  Queue last_q_195 ( // @[Decoupled.scala 361:21]
    .clock(last_q_195_clock),
    .reset(last_q_195_reset),
    .io_enq_ready(last_q_195_io_enq_ready),
    .io_enq_valid(last_q_195_io_enq_valid),
    .io_enq_bits(last_q_195_io_enq_bits),
    .io_deq_ready(last_q_195_io_deq_ready),
    .io_deq_valid(last_q_195_io_deq_valid),
    .io_deq_bits(last_q_195_io_deq_bits)
  );
  StreamMerger_196 last_merger_196 ( // @[Stab.scala 175:24]
    .clock(last_merger_196_clock),
    .reset(last_merger_196_reset),
    .io_stream1_ready(last_merger_196_io_stream1_ready),
    .io_stream1_valid(last_merger_196_io_stream1_valid),
    .io_stream1_bits(last_merger_196_io_stream1_bits),
    .io_stream2_ready(last_merger_196_io_stream2_ready),
    .io_stream2_valid(last_merger_196_io_stream2_valid),
    .io_stream2_bits(last_merger_196_io_stream2_bits),
    .io_result_ready(last_merger_196_io_result_ready),
    .io_result_valid(last_merger_196_io_result_valid),
    .io_result_bits(last_merger_196_io_result_bits)
  );
  Queue last_q_196 ( // @[Decoupled.scala 361:21]
    .clock(last_q_196_clock),
    .reset(last_q_196_reset),
    .io_enq_ready(last_q_196_io_enq_ready),
    .io_enq_valid(last_q_196_io_enq_valid),
    .io_enq_bits(last_q_196_io_enq_bits),
    .io_deq_ready(last_q_196_io_deq_ready),
    .io_deq_valid(last_q_196_io_deq_valid),
    .io_deq_bits(last_q_196_io_deq_bits)
  );
  StreamMerger_197 last_merger_197 ( // @[Stab.scala 175:24]
    .clock(last_merger_197_clock),
    .reset(last_merger_197_reset),
    .io_stream1_ready(last_merger_197_io_stream1_ready),
    .io_stream1_valid(last_merger_197_io_stream1_valid),
    .io_stream1_bits(last_merger_197_io_stream1_bits),
    .io_stream2_ready(last_merger_197_io_stream2_ready),
    .io_stream2_valid(last_merger_197_io_stream2_valid),
    .io_stream2_bits(last_merger_197_io_stream2_bits),
    .io_result_ready(last_merger_197_io_result_ready),
    .io_result_valid(last_merger_197_io_result_valid),
    .io_result_bits(last_merger_197_io_result_bits)
  );
  Queue last_q_197 ( // @[Decoupled.scala 361:21]
    .clock(last_q_197_clock),
    .reset(last_q_197_reset),
    .io_enq_ready(last_q_197_io_enq_ready),
    .io_enq_valid(last_q_197_io_enq_valid),
    .io_enq_bits(last_q_197_io_enq_bits),
    .io_deq_ready(last_q_197_io_deq_ready),
    .io_deq_valid(last_q_197_io_deq_valid),
    .io_deq_bits(last_q_197_io_deq_bits)
  );
  StreamMerger_198 last_merger_198 ( // @[Stab.scala 175:24]
    .clock(last_merger_198_clock),
    .reset(last_merger_198_reset),
    .io_stream1_ready(last_merger_198_io_stream1_ready),
    .io_stream1_valid(last_merger_198_io_stream1_valid),
    .io_stream1_bits(last_merger_198_io_stream1_bits),
    .io_stream2_ready(last_merger_198_io_stream2_ready),
    .io_stream2_valid(last_merger_198_io_stream2_valid),
    .io_stream2_bits(last_merger_198_io_stream2_bits),
    .io_result_ready(last_merger_198_io_result_ready),
    .io_result_valid(last_merger_198_io_result_valid),
    .io_result_bits(last_merger_198_io_result_bits)
  );
  Queue last_q_198 ( // @[Decoupled.scala 361:21]
    .clock(last_q_198_clock),
    .reset(last_q_198_reset),
    .io_enq_ready(last_q_198_io_enq_ready),
    .io_enq_valid(last_q_198_io_enq_valid),
    .io_enq_bits(last_q_198_io_enq_bits),
    .io_deq_ready(last_q_198_io_deq_ready),
    .io_deq_valid(last_q_198_io_deq_valid),
    .io_deq_bits(last_q_198_io_deq_bits)
  );
  StreamMerger_199 last_merger_199 ( // @[Stab.scala 175:24]
    .clock(last_merger_199_clock),
    .reset(last_merger_199_reset),
    .io_stream1_ready(last_merger_199_io_stream1_ready),
    .io_stream1_valid(last_merger_199_io_stream1_valid),
    .io_stream1_bits(last_merger_199_io_stream1_bits),
    .io_stream2_ready(last_merger_199_io_stream2_ready),
    .io_stream2_valid(last_merger_199_io_stream2_valid),
    .io_stream2_bits(last_merger_199_io_stream2_bits),
    .io_result_ready(last_merger_199_io_result_ready),
    .io_result_valid(last_merger_199_io_result_valid),
    .io_result_bits(last_merger_199_io_result_bits)
  );
  Queue last_q_199 ( // @[Decoupled.scala 361:21]
    .clock(last_q_199_clock),
    .reset(last_q_199_reset),
    .io_enq_ready(last_q_199_io_enq_ready),
    .io_enq_valid(last_q_199_io_enq_valid),
    .io_enq_bits(last_q_199_io_enq_bits),
    .io_deq_ready(last_q_199_io_deq_ready),
    .io_deq_valid(last_q_199_io_deq_valid),
    .io_deq_bits(last_q_199_io_deq_bits)
  );
  StreamMerger_200 last_merger_200 ( // @[Stab.scala 175:24]
    .clock(last_merger_200_clock),
    .reset(last_merger_200_reset),
    .io_stream1_ready(last_merger_200_io_stream1_ready),
    .io_stream1_valid(last_merger_200_io_stream1_valid),
    .io_stream1_bits(last_merger_200_io_stream1_bits),
    .io_stream2_ready(last_merger_200_io_stream2_ready),
    .io_stream2_valid(last_merger_200_io_stream2_valid),
    .io_stream2_bits(last_merger_200_io_stream2_bits),
    .io_result_ready(last_merger_200_io_result_ready),
    .io_result_valid(last_merger_200_io_result_valid),
    .io_result_bits(last_merger_200_io_result_bits)
  );
  Queue last_q_200 ( // @[Decoupled.scala 361:21]
    .clock(last_q_200_clock),
    .reset(last_q_200_reset),
    .io_enq_ready(last_q_200_io_enq_ready),
    .io_enq_valid(last_q_200_io_enq_valid),
    .io_enq_bits(last_q_200_io_enq_bits),
    .io_deq_ready(last_q_200_io_deq_ready),
    .io_deq_valid(last_q_200_io_deq_valid),
    .io_deq_bits(last_q_200_io_deq_bits)
  );
  StreamMerger_201 last_merger_201 ( // @[Stab.scala 175:24]
    .clock(last_merger_201_clock),
    .reset(last_merger_201_reset),
    .io_stream1_ready(last_merger_201_io_stream1_ready),
    .io_stream1_valid(last_merger_201_io_stream1_valid),
    .io_stream1_bits(last_merger_201_io_stream1_bits),
    .io_stream2_ready(last_merger_201_io_stream2_ready),
    .io_stream2_valid(last_merger_201_io_stream2_valid),
    .io_stream2_bits(last_merger_201_io_stream2_bits),
    .io_result_ready(last_merger_201_io_result_ready),
    .io_result_valid(last_merger_201_io_result_valid),
    .io_result_bits(last_merger_201_io_result_bits)
  );
  Queue last_q_201 ( // @[Decoupled.scala 361:21]
    .clock(last_q_201_clock),
    .reset(last_q_201_reset),
    .io_enq_ready(last_q_201_io_enq_ready),
    .io_enq_valid(last_q_201_io_enq_valid),
    .io_enq_bits(last_q_201_io_enq_bits),
    .io_deq_ready(last_q_201_io_deq_ready),
    .io_deq_valid(last_q_201_io_deq_valid),
    .io_deq_bits(last_q_201_io_deq_bits)
  );
  StreamMerger_202 last_merger_202 ( // @[Stab.scala 175:24]
    .clock(last_merger_202_clock),
    .reset(last_merger_202_reset),
    .io_stream1_ready(last_merger_202_io_stream1_ready),
    .io_stream1_valid(last_merger_202_io_stream1_valid),
    .io_stream1_bits(last_merger_202_io_stream1_bits),
    .io_stream2_ready(last_merger_202_io_stream2_ready),
    .io_stream2_valid(last_merger_202_io_stream2_valid),
    .io_stream2_bits(last_merger_202_io_stream2_bits),
    .io_result_ready(last_merger_202_io_result_ready),
    .io_result_valid(last_merger_202_io_result_valid),
    .io_result_bits(last_merger_202_io_result_bits)
  );
  Queue last_q_202 ( // @[Decoupled.scala 361:21]
    .clock(last_q_202_clock),
    .reset(last_q_202_reset),
    .io_enq_ready(last_q_202_io_enq_ready),
    .io_enq_valid(last_q_202_io_enq_valid),
    .io_enq_bits(last_q_202_io_enq_bits),
    .io_deq_ready(last_q_202_io_deq_ready),
    .io_deq_valid(last_q_202_io_deq_valid),
    .io_deq_bits(last_q_202_io_deq_bits)
  );
  StreamMerger_203 last_merger_203 ( // @[Stab.scala 175:24]
    .clock(last_merger_203_clock),
    .reset(last_merger_203_reset),
    .io_stream1_ready(last_merger_203_io_stream1_ready),
    .io_stream1_valid(last_merger_203_io_stream1_valid),
    .io_stream1_bits(last_merger_203_io_stream1_bits),
    .io_stream2_ready(last_merger_203_io_stream2_ready),
    .io_stream2_valid(last_merger_203_io_stream2_valid),
    .io_stream2_bits(last_merger_203_io_stream2_bits),
    .io_result_ready(last_merger_203_io_result_ready),
    .io_result_valid(last_merger_203_io_result_valid),
    .io_result_bits(last_merger_203_io_result_bits)
  );
  Queue last_q_203 ( // @[Decoupled.scala 361:21]
    .clock(last_q_203_clock),
    .reset(last_q_203_reset),
    .io_enq_ready(last_q_203_io_enq_ready),
    .io_enq_valid(last_q_203_io_enq_valid),
    .io_enq_bits(last_q_203_io_enq_bits),
    .io_deq_ready(last_q_203_io_deq_ready),
    .io_deq_valid(last_q_203_io_deq_valid),
    .io_deq_bits(last_q_203_io_deq_bits)
  );
  StreamMerger_204 last_merger_204 ( // @[Stab.scala 175:24]
    .clock(last_merger_204_clock),
    .reset(last_merger_204_reset),
    .io_stream1_ready(last_merger_204_io_stream1_ready),
    .io_stream1_valid(last_merger_204_io_stream1_valid),
    .io_stream1_bits(last_merger_204_io_stream1_bits),
    .io_stream2_ready(last_merger_204_io_stream2_ready),
    .io_stream2_valid(last_merger_204_io_stream2_valid),
    .io_stream2_bits(last_merger_204_io_stream2_bits),
    .io_result_ready(last_merger_204_io_result_ready),
    .io_result_valid(last_merger_204_io_result_valid),
    .io_result_bits(last_merger_204_io_result_bits)
  );
  Queue last_q_204 ( // @[Decoupled.scala 361:21]
    .clock(last_q_204_clock),
    .reset(last_q_204_reset),
    .io_enq_ready(last_q_204_io_enq_ready),
    .io_enq_valid(last_q_204_io_enq_valid),
    .io_enq_bits(last_q_204_io_enq_bits),
    .io_deq_ready(last_q_204_io_deq_ready),
    .io_deq_valid(last_q_204_io_deq_valid),
    .io_deq_bits(last_q_204_io_deq_bits)
  );
  StreamMerger_205 last_merger_205 ( // @[Stab.scala 175:24]
    .clock(last_merger_205_clock),
    .reset(last_merger_205_reset),
    .io_stream1_ready(last_merger_205_io_stream1_ready),
    .io_stream1_valid(last_merger_205_io_stream1_valid),
    .io_stream1_bits(last_merger_205_io_stream1_bits),
    .io_stream2_ready(last_merger_205_io_stream2_ready),
    .io_stream2_valid(last_merger_205_io_stream2_valid),
    .io_stream2_bits(last_merger_205_io_stream2_bits),
    .io_result_ready(last_merger_205_io_result_ready),
    .io_result_valid(last_merger_205_io_result_valid),
    .io_result_bits(last_merger_205_io_result_bits)
  );
  Queue last_q_205 ( // @[Decoupled.scala 361:21]
    .clock(last_q_205_clock),
    .reset(last_q_205_reset),
    .io_enq_ready(last_q_205_io_enq_ready),
    .io_enq_valid(last_q_205_io_enq_valid),
    .io_enq_bits(last_q_205_io_enq_bits),
    .io_deq_ready(last_q_205_io_deq_ready),
    .io_deq_valid(last_q_205_io_deq_valid),
    .io_deq_bits(last_q_205_io_deq_bits)
  );
  StreamMerger_206 last_merger_206 ( // @[Stab.scala 175:24]
    .clock(last_merger_206_clock),
    .reset(last_merger_206_reset),
    .io_stream1_ready(last_merger_206_io_stream1_ready),
    .io_stream1_valid(last_merger_206_io_stream1_valid),
    .io_stream1_bits(last_merger_206_io_stream1_bits),
    .io_stream2_ready(last_merger_206_io_stream2_ready),
    .io_stream2_valid(last_merger_206_io_stream2_valid),
    .io_stream2_bits(last_merger_206_io_stream2_bits),
    .io_result_ready(last_merger_206_io_result_ready),
    .io_result_valid(last_merger_206_io_result_valid),
    .io_result_bits(last_merger_206_io_result_bits)
  );
  Queue last_q_206 ( // @[Decoupled.scala 361:21]
    .clock(last_q_206_clock),
    .reset(last_q_206_reset),
    .io_enq_ready(last_q_206_io_enq_ready),
    .io_enq_valid(last_q_206_io_enq_valid),
    .io_enq_bits(last_q_206_io_enq_bits),
    .io_deq_ready(last_q_206_io_deq_ready),
    .io_deq_valid(last_q_206_io_deq_valid),
    .io_deq_bits(last_q_206_io_deq_bits)
  );
  StreamMerger_207 last_merger_207 ( // @[Stab.scala 175:24]
    .clock(last_merger_207_clock),
    .reset(last_merger_207_reset),
    .io_stream1_ready(last_merger_207_io_stream1_ready),
    .io_stream1_valid(last_merger_207_io_stream1_valid),
    .io_stream1_bits(last_merger_207_io_stream1_bits),
    .io_stream2_ready(last_merger_207_io_stream2_ready),
    .io_stream2_valid(last_merger_207_io_stream2_valid),
    .io_stream2_bits(last_merger_207_io_stream2_bits),
    .io_result_ready(last_merger_207_io_result_ready),
    .io_result_valid(last_merger_207_io_result_valid),
    .io_result_bits(last_merger_207_io_result_bits)
  );
  Queue last_q_207 ( // @[Decoupled.scala 361:21]
    .clock(last_q_207_clock),
    .reset(last_q_207_reset),
    .io_enq_ready(last_q_207_io_enq_ready),
    .io_enq_valid(last_q_207_io_enq_valid),
    .io_enq_bits(last_q_207_io_enq_bits),
    .io_deq_ready(last_q_207_io_deq_ready),
    .io_deq_valid(last_q_207_io_deq_valid),
    .io_deq_bits(last_q_207_io_deq_bits)
  );
  StreamMerger_208 last_merger_208 ( // @[Stab.scala 175:24]
    .clock(last_merger_208_clock),
    .reset(last_merger_208_reset),
    .io_stream1_ready(last_merger_208_io_stream1_ready),
    .io_stream1_valid(last_merger_208_io_stream1_valid),
    .io_stream1_bits(last_merger_208_io_stream1_bits),
    .io_stream2_ready(last_merger_208_io_stream2_ready),
    .io_stream2_valid(last_merger_208_io_stream2_valid),
    .io_stream2_bits(last_merger_208_io_stream2_bits),
    .io_result_ready(last_merger_208_io_result_ready),
    .io_result_valid(last_merger_208_io_result_valid),
    .io_result_bits(last_merger_208_io_result_bits)
  );
  Queue last_q_208 ( // @[Decoupled.scala 361:21]
    .clock(last_q_208_clock),
    .reset(last_q_208_reset),
    .io_enq_ready(last_q_208_io_enq_ready),
    .io_enq_valid(last_q_208_io_enq_valid),
    .io_enq_bits(last_q_208_io_enq_bits),
    .io_deq_ready(last_q_208_io_deq_ready),
    .io_deq_valid(last_q_208_io_deq_valid),
    .io_deq_bits(last_q_208_io_deq_bits)
  );
  StreamMerger_209 last_merger_209 ( // @[Stab.scala 175:24]
    .clock(last_merger_209_clock),
    .reset(last_merger_209_reset),
    .io_stream1_ready(last_merger_209_io_stream1_ready),
    .io_stream1_valid(last_merger_209_io_stream1_valid),
    .io_stream1_bits(last_merger_209_io_stream1_bits),
    .io_stream2_ready(last_merger_209_io_stream2_ready),
    .io_stream2_valid(last_merger_209_io_stream2_valid),
    .io_stream2_bits(last_merger_209_io_stream2_bits),
    .io_result_ready(last_merger_209_io_result_ready),
    .io_result_valid(last_merger_209_io_result_valid),
    .io_result_bits(last_merger_209_io_result_bits)
  );
  Queue last_q_209 ( // @[Decoupled.scala 361:21]
    .clock(last_q_209_clock),
    .reset(last_q_209_reset),
    .io_enq_ready(last_q_209_io_enq_ready),
    .io_enq_valid(last_q_209_io_enq_valid),
    .io_enq_bits(last_q_209_io_enq_bits),
    .io_deq_ready(last_q_209_io_deq_ready),
    .io_deq_valid(last_q_209_io_deq_valid),
    .io_deq_bits(last_q_209_io_deq_bits)
  );
  StreamMerger_210 last_merger_210 ( // @[Stab.scala 175:24]
    .clock(last_merger_210_clock),
    .reset(last_merger_210_reset),
    .io_stream1_ready(last_merger_210_io_stream1_ready),
    .io_stream1_valid(last_merger_210_io_stream1_valid),
    .io_stream1_bits(last_merger_210_io_stream1_bits),
    .io_stream2_ready(last_merger_210_io_stream2_ready),
    .io_stream2_valid(last_merger_210_io_stream2_valid),
    .io_stream2_bits(last_merger_210_io_stream2_bits),
    .io_result_ready(last_merger_210_io_result_ready),
    .io_result_valid(last_merger_210_io_result_valid),
    .io_result_bits(last_merger_210_io_result_bits)
  );
  Queue last_q_210 ( // @[Decoupled.scala 361:21]
    .clock(last_q_210_clock),
    .reset(last_q_210_reset),
    .io_enq_ready(last_q_210_io_enq_ready),
    .io_enq_valid(last_q_210_io_enq_valid),
    .io_enq_bits(last_q_210_io_enq_bits),
    .io_deq_ready(last_q_210_io_deq_ready),
    .io_deq_valid(last_q_210_io_deq_valid),
    .io_deq_bits(last_q_210_io_deq_bits)
  );
  StreamMerger_211 last_merger_211 ( // @[Stab.scala 175:24]
    .clock(last_merger_211_clock),
    .reset(last_merger_211_reset),
    .io_stream1_ready(last_merger_211_io_stream1_ready),
    .io_stream1_valid(last_merger_211_io_stream1_valid),
    .io_stream1_bits(last_merger_211_io_stream1_bits),
    .io_stream2_ready(last_merger_211_io_stream2_ready),
    .io_stream2_valid(last_merger_211_io_stream2_valid),
    .io_stream2_bits(last_merger_211_io_stream2_bits),
    .io_result_ready(last_merger_211_io_result_ready),
    .io_result_valid(last_merger_211_io_result_valid),
    .io_result_bits(last_merger_211_io_result_bits)
  );
  Queue last_q_211 ( // @[Decoupled.scala 361:21]
    .clock(last_q_211_clock),
    .reset(last_q_211_reset),
    .io_enq_ready(last_q_211_io_enq_ready),
    .io_enq_valid(last_q_211_io_enq_valid),
    .io_enq_bits(last_q_211_io_enq_bits),
    .io_deq_ready(last_q_211_io_deq_ready),
    .io_deq_valid(last_q_211_io_deq_valid),
    .io_deq_bits(last_q_211_io_deq_bits)
  );
  StreamMerger_212 last_merger_212 ( // @[Stab.scala 175:24]
    .clock(last_merger_212_clock),
    .reset(last_merger_212_reset),
    .io_stream1_ready(last_merger_212_io_stream1_ready),
    .io_stream1_valid(last_merger_212_io_stream1_valid),
    .io_stream1_bits(last_merger_212_io_stream1_bits),
    .io_stream2_ready(last_merger_212_io_stream2_ready),
    .io_stream2_valid(last_merger_212_io_stream2_valid),
    .io_stream2_bits(last_merger_212_io_stream2_bits),
    .io_result_ready(last_merger_212_io_result_ready),
    .io_result_valid(last_merger_212_io_result_valid),
    .io_result_bits(last_merger_212_io_result_bits)
  );
  Queue last_q_212 ( // @[Decoupled.scala 361:21]
    .clock(last_q_212_clock),
    .reset(last_q_212_reset),
    .io_enq_ready(last_q_212_io_enq_ready),
    .io_enq_valid(last_q_212_io_enq_valid),
    .io_enq_bits(last_q_212_io_enq_bits),
    .io_deq_ready(last_q_212_io_deq_ready),
    .io_deq_valid(last_q_212_io_deq_valid),
    .io_deq_bits(last_q_212_io_deq_bits)
  );
  StreamMerger_213 last_merger_213 ( // @[Stab.scala 175:24]
    .clock(last_merger_213_clock),
    .reset(last_merger_213_reset),
    .io_stream1_ready(last_merger_213_io_stream1_ready),
    .io_stream1_valid(last_merger_213_io_stream1_valid),
    .io_stream1_bits(last_merger_213_io_stream1_bits),
    .io_stream2_ready(last_merger_213_io_stream2_ready),
    .io_stream2_valid(last_merger_213_io_stream2_valid),
    .io_stream2_bits(last_merger_213_io_stream2_bits),
    .io_result_ready(last_merger_213_io_result_ready),
    .io_result_valid(last_merger_213_io_result_valid),
    .io_result_bits(last_merger_213_io_result_bits)
  );
  Queue last_q_213 ( // @[Decoupled.scala 361:21]
    .clock(last_q_213_clock),
    .reset(last_q_213_reset),
    .io_enq_ready(last_q_213_io_enq_ready),
    .io_enq_valid(last_q_213_io_enq_valid),
    .io_enq_bits(last_q_213_io_enq_bits),
    .io_deq_ready(last_q_213_io_deq_ready),
    .io_deq_valid(last_q_213_io_deq_valid),
    .io_deq_bits(last_q_213_io_deq_bits)
  );
  StreamMerger_214 last_merger_214 ( // @[Stab.scala 175:24]
    .clock(last_merger_214_clock),
    .reset(last_merger_214_reset),
    .io_stream1_ready(last_merger_214_io_stream1_ready),
    .io_stream1_valid(last_merger_214_io_stream1_valid),
    .io_stream1_bits(last_merger_214_io_stream1_bits),
    .io_stream2_ready(last_merger_214_io_stream2_ready),
    .io_stream2_valid(last_merger_214_io_stream2_valid),
    .io_stream2_bits(last_merger_214_io_stream2_bits),
    .io_result_ready(last_merger_214_io_result_ready),
    .io_result_valid(last_merger_214_io_result_valid),
    .io_result_bits(last_merger_214_io_result_bits)
  );
  Queue last_q_214 ( // @[Decoupled.scala 361:21]
    .clock(last_q_214_clock),
    .reset(last_q_214_reset),
    .io_enq_ready(last_q_214_io_enq_ready),
    .io_enq_valid(last_q_214_io_enq_valid),
    .io_enq_bits(last_q_214_io_enq_bits),
    .io_deq_ready(last_q_214_io_deq_ready),
    .io_deq_valid(last_q_214_io_deq_valid),
    .io_deq_bits(last_q_214_io_deq_bits)
  );
  StreamMerger_215 last_merger_215 ( // @[Stab.scala 175:24]
    .clock(last_merger_215_clock),
    .reset(last_merger_215_reset),
    .io_stream1_ready(last_merger_215_io_stream1_ready),
    .io_stream1_valid(last_merger_215_io_stream1_valid),
    .io_stream1_bits(last_merger_215_io_stream1_bits),
    .io_stream2_ready(last_merger_215_io_stream2_ready),
    .io_stream2_valid(last_merger_215_io_stream2_valid),
    .io_stream2_bits(last_merger_215_io_stream2_bits),
    .io_result_ready(last_merger_215_io_result_ready),
    .io_result_valid(last_merger_215_io_result_valid),
    .io_result_bits(last_merger_215_io_result_bits)
  );
  Queue last_q_215 ( // @[Decoupled.scala 361:21]
    .clock(last_q_215_clock),
    .reset(last_q_215_reset),
    .io_enq_ready(last_q_215_io_enq_ready),
    .io_enq_valid(last_q_215_io_enq_valid),
    .io_enq_bits(last_q_215_io_enq_bits),
    .io_deq_ready(last_q_215_io_deq_ready),
    .io_deq_valid(last_q_215_io_deq_valid),
    .io_deq_bits(last_q_215_io_deq_bits)
  );
  StreamMerger_216 last_merger_216 ( // @[Stab.scala 175:24]
    .clock(last_merger_216_clock),
    .reset(last_merger_216_reset),
    .io_stream1_ready(last_merger_216_io_stream1_ready),
    .io_stream1_valid(last_merger_216_io_stream1_valid),
    .io_stream1_bits(last_merger_216_io_stream1_bits),
    .io_stream2_ready(last_merger_216_io_stream2_ready),
    .io_stream2_valid(last_merger_216_io_stream2_valid),
    .io_stream2_bits(last_merger_216_io_stream2_bits),
    .io_result_ready(last_merger_216_io_result_ready),
    .io_result_valid(last_merger_216_io_result_valid),
    .io_result_bits(last_merger_216_io_result_bits)
  );
  Queue last_q_216 ( // @[Decoupled.scala 361:21]
    .clock(last_q_216_clock),
    .reset(last_q_216_reset),
    .io_enq_ready(last_q_216_io_enq_ready),
    .io_enq_valid(last_q_216_io_enq_valid),
    .io_enq_bits(last_q_216_io_enq_bits),
    .io_deq_ready(last_q_216_io_deq_ready),
    .io_deq_valid(last_q_216_io_deq_valid),
    .io_deq_bits(last_q_216_io_deq_bits)
  );
  StreamMerger_217 last_merger_217 ( // @[Stab.scala 175:24]
    .clock(last_merger_217_clock),
    .reset(last_merger_217_reset),
    .io_stream1_ready(last_merger_217_io_stream1_ready),
    .io_stream1_valid(last_merger_217_io_stream1_valid),
    .io_stream1_bits(last_merger_217_io_stream1_bits),
    .io_stream2_ready(last_merger_217_io_stream2_ready),
    .io_stream2_valid(last_merger_217_io_stream2_valid),
    .io_stream2_bits(last_merger_217_io_stream2_bits),
    .io_result_ready(last_merger_217_io_result_ready),
    .io_result_valid(last_merger_217_io_result_valid),
    .io_result_bits(last_merger_217_io_result_bits)
  );
  Queue last_q_217 ( // @[Decoupled.scala 361:21]
    .clock(last_q_217_clock),
    .reset(last_q_217_reset),
    .io_enq_ready(last_q_217_io_enq_ready),
    .io_enq_valid(last_q_217_io_enq_valid),
    .io_enq_bits(last_q_217_io_enq_bits),
    .io_deq_ready(last_q_217_io_deq_ready),
    .io_deq_valid(last_q_217_io_deq_valid),
    .io_deq_bits(last_q_217_io_deq_bits)
  );
  StreamMerger_218 last_merger_218 ( // @[Stab.scala 175:24]
    .clock(last_merger_218_clock),
    .reset(last_merger_218_reset),
    .io_stream1_ready(last_merger_218_io_stream1_ready),
    .io_stream1_valid(last_merger_218_io_stream1_valid),
    .io_stream1_bits(last_merger_218_io_stream1_bits),
    .io_stream2_ready(last_merger_218_io_stream2_ready),
    .io_stream2_valid(last_merger_218_io_stream2_valid),
    .io_stream2_bits(last_merger_218_io_stream2_bits),
    .io_result_ready(last_merger_218_io_result_ready),
    .io_result_valid(last_merger_218_io_result_valid),
    .io_result_bits(last_merger_218_io_result_bits)
  );
  Queue last_q_218 ( // @[Decoupled.scala 361:21]
    .clock(last_q_218_clock),
    .reset(last_q_218_reset),
    .io_enq_ready(last_q_218_io_enq_ready),
    .io_enq_valid(last_q_218_io_enq_valid),
    .io_enq_bits(last_q_218_io_enq_bits),
    .io_deq_ready(last_q_218_io_deq_ready),
    .io_deq_valid(last_q_218_io_deq_valid),
    .io_deq_bits(last_q_218_io_deq_bits)
  );
  StreamMerger_219 last_merger_219 ( // @[Stab.scala 175:24]
    .clock(last_merger_219_clock),
    .reset(last_merger_219_reset),
    .io_stream1_ready(last_merger_219_io_stream1_ready),
    .io_stream1_valid(last_merger_219_io_stream1_valid),
    .io_stream1_bits(last_merger_219_io_stream1_bits),
    .io_stream2_ready(last_merger_219_io_stream2_ready),
    .io_stream2_valid(last_merger_219_io_stream2_valid),
    .io_stream2_bits(last_merger_219_io_stream2_bits),
    .io_result_ready(last_merger_219_io_result_ready),
    .io_result_valid(last_merger_219_io_result_valid),
    .io_result_bits(last_merger_219_io_result_bits)
  );
  Queue last_q_219 ( // @[Decoupled.scala 361:21]
    .clock(last_q_219_clock),
    .reset(last_q_219_reset),
    .io_enq_ready(last_q_219_io_enq_ready),
    .io_enq_valid(last_q_219_io_enq_valid),
    .io_enq_bits(last_q_219_io_enq_bits),
    .io_deq_ready(last_q_219_io_deq_ready),
    .io_deq_valid(last_q_219_io_deq_valid),
    .io_deq_bits(last_q_219_io_deq_bits)
  );
  StreamMerger_220 last_merger_220 ( // @[Stab.scala 175:24]
    .clock(last_merger_220_clock),
    .reset(last_merger_220_reset),
    .io_stream1_ready(last_merger_220_io_stream1_ready),
    .io_stream1_valid(last_merger_220_io_stream1_valid),
    .io_stream1_bits(last_merger_220_io_stream1_bits),
    .io_stream2_ready(last_merger_220_io_stream2_ready),
    .io_stream2_valid(last_merger_220_io_stream2_valid),
    .io_stream2_bits(last_merger_220_io_stream2_bits),
    .io_result_ready(last_merger_220_io_result_ready),
    .io_result_valid(last_merger_220_io_result_valid),
    .io_result_bits(last_merger_220_io_result_bits)
  );
  Queue last_q_220 ( // @[Decoupled.scala 361:21]
    .clock(last_q_220_clock),
    .reset(last_q_220_reset),
    .io_enq_ready(last_q_220_io_enq_ready),
    .io_enq_valid(last_q_220_io_enq_valid),
    .io_enq_bits(last_q_220_io_enq_bits),
    .io_deq_ready(last_q_220_io_deq_ready),
    .io_deq_valid(last_q_220_io_deq_valid),
    .io_deq_bits(last_q_220_io_deq_bits)
  );
  StreamMerger_221 last_merger_221 ( // @[Stab.scala 175:24]
    .clock(last_merger_221_clock),
    .reset(last_merger_221_reset),
    .io_stream1_ready(last_merger_221_io_stream1_ready),
    .io_stream1_valid(last_merger_221_io_stream1_valid),
    .io_stream1_bits(last_merger_221_io_stream1_bits),
    .io_stream2_ready(last_merger_221_io_stream2_ready),
    .io_stream2_valid(last_merger_221_io_stream2_valid),
    .io_stream2_bits(last_merger_221_io_stream2_bits),
    .io_result_ready(last_merger_221_io_result_ready),
    .io_result_valid(last_merger_221_io_result_valid),
    .io_result_bits(last_merger_221_io_result_bits)
  );
  Queue last_q_221 ( // @[Decoupled.scala 361:21]
    .clock(last_q_221_clock),
    .reset(last_q_221_reset),
    .io_enq_ready(last_q_221_io_enq_ready),
    .io_enq_valid(last_q_221_io_enq_valid),
    .io_enq_bits(last_q_221_io_enq_bits),
    .io_deq_ready(last_q_221_io_deq_ready),
    .io_deq_valid(last_q_221_io_deq_valid),
    .io_deq_bits(last_q_221_io_deq_bits)
  );
  StreamMerger_222 last_merger_222 ( // @[Stab.scala 175:24]
    .clock(last_merger_222_clock),
    .reset(last_merger_222_reset),
    .io_stream1_ready(last_merger_222_io_stream1_ready),
    .io_stream1_valid(last_merger_222_io_stream1_valid),
    .io_stream1_bits(last_merger_222_io_stream1_bits),
    .io_stream2_ready(last_merger_222_io_stream2_ready),
    .io_stream2_valid(last_merger_222_io_stream2_valid),
    .io_stream2_bits(last_merger_222_io_stream2_bits),
    .io_result_ready(last_merger_222_io_result_ready),
    .io_result_valid(last_merger_222_io_result_valid),
    .io_result_bits(last_merger_222_io_result_bits)
  );
  Queue last_q_222 ( // @[Decoupled.scala 361:21]
    .clock(last_q_222_clock),
    .reset(last_q_222_reset),
    .io_enq_ready(last_q_222_io_enq_ready),
    .io_enq_valid(last_q_222_io_enq_valid),
    .io_enq_bits(last_q_222_io_enq_bits),
    .io_deq_ready(last_q_222_io_deq_ready),
    .io_deq_valid(last_q_222_io_deq_valid),
    .io_deq_bits(last_q_222_io_deq_bits)
  );
  StreamMerger_223 last_merger_223 ( // @[Stab.scala 175:24]
    .clock(last_merger_223_clock),
    .reset(last_merger_223_reset),
    .io_stream1_ready(last_merger_223_io_stream1_ready),
    .io_stream1_valid(last_merger_223_io_stream1_valid),
    .io_stream1_bits(last_merger_223_io_stream1_bits),
    .io_stream2_ready(last_merger_223_io_stream2_ready),
    .io_stream2_valid(last_merger_223_io_stream2_valid),
    .io_stream2_bits(last_merger_223_io_stream2_bits),
    .io_result_ready(last_merger_223_io_result_ready),
    .io_result_valid(last_merger_223_io_result_valid),
    .io_result_bits(last_merger_223_io_result_bits)
  );
  Queue last_q_223 ( // @[Decoupled.scala 361:21]
    .clock(last_q_223_clock),
    .reset(last_q_223_reset),
    .io_enq_ready(last_q_223_io_enq_ready),
    .io_enq_valid(last_q_223_io_enq_valid),
    .io_enq_bits(last_q_223_io_enq_bits),
    .io_deq_ready(last_q_223_io_deq_ready),
    .io_deq_valid(last_q_223_io_deq_valid),
    .io_deq_bits(last_q_223_io_deq_bits)
  );
  StreamMerger_224 last_merger_224 ( // @[Stab.scala 175:24]
    .clock(last_merger_224_clock),
    .reset(last_merger_224_reset),
    .io_stream1_ready(last_merger_224_io_stream1_ready),
    .io_stream1_valid(last_merger_224_io_stream1_valid),
    .io_stream1_bits(last_merger_224_io_stream1_bits),
    .io_stream2_ready(last_merger_224_io_stream2_ready),
    .io_stream2_valid(last_merger_224_io_stream2_valid),
    .io_stream2_bits(last_merger_224_io_stream2_bits),
    .io_result_ready(last_merger_224_io_result_ready),
    .io_result_valid(last_merger_224_io_result_valid),
    .io_result_bits(last_merger_224_io_result_bits)
  );
  Queue last_q_224 ( // @[Decoupled.scala 361:21]
    .clock(last_q_224_clock),
    .reset(last_q_224_reset),
    .io_enq_ready(last_q_224_io_enq_ready),
    .io_enq_valid(last_q_224_io_enq_valid),
    .io_enq_bits(last_q_224_io_enq_bits),
    .io_deq_ready(last_q_224_io_deq_ready),
    .io_deq_valid(last_q_224_io_deq_valid),
    .io_deq_bits(last_q_224_io_deq_bits)
  );
  StreamMerger_225 last_merger_225 ( // @[Stab.scala 175:24]
    .clock(last_merger_225_clock),
    .reset(last_merger_225_reset),
    .io_stream1_ready(last_merger_225_io_stream1_ready),
    .io_stream1_valid(last_merger_225_io_stream1_valid),
    .io_stream1_bits(last_merger_225_io_stream1_bits),
    .io_stream2_ready(last_merger_225_io_stream2_ready),
    .io_stream2_valid(last_merger_225_io_stream2_valid),
    .io_stream2_bits(last_merger_225_io_stream2_bits),
    .io_result_ready(last_merger_225_io_result_ready),
    .io_result_valid(last_merger_225_io_result_valid),
    .io_result_bits(last_merger_225_io_result_bits)
  );
  Queue last_q_225 ( // @[Decoupled.scala 361:21]
    .clock(last_q_225_clock),
    .reset(last_q_225_reset),
    .io_enq_ready(last_q_225_io_enq_ready),
    .io_enq_valid(last_q_225_io_enq_valid),
    .io_enq_bits(last_q_225_io_enq_bits),
    .io_deq_ready(last_q_225_io_deq_ready),
    .io_deq_valid(last_q_225_io_deq_valid),
    .io_deq_bits(last_q_225_io_deq_bits)
  );
  StreamMerger_226 last_merger_226 ( // @[Stab.scala 175:24]
    .clock(last_merger_226_clock),
    .reset(last_merger_226_reset),
    .io_stream1_ready(last_merger_226_io_stream1_ready),
    .io_stream1_valid(last_merger_226_io_stream1_valid),
    .io_stream1_bits(last_merger_226_io_stream1_bits),
    .io_stream2_ready(last_merger_226_io_stream2_ready),
    .io_stream2_valid(last_merger_226_io_stream2_valid),
    .io_stream2_bits(last_merger_226_io_stream2_bits),
    .io_result_ready(last_merger_226_io_result_ready),
    .io_result_valid(last_merger_226_io_result_valid),
    .io_result_bits(last_merger_226_io_result_bits)
  );
  Queue last_q_226 ( // @[Decoupled.scala 361:21]
    .clock(last_q_226_clock),
    .reset(last_q_226_reset),
    .io_enq_ready(last_q_226_io_enq_ready),
    .io_enq_valid(last_q_226_io_enq_valid),
    .io_enq_bits(last_q_226_io_enq_bits),
    .io_deq_ready(last_q_226_io_deq_ready),
    .io_deq_valid(last_q_226_io_deq_valid),
    .io_deq_bits(last_q_226_io_deq_bits)
  );
  StreamMerger_227 last_merger_227 ( // @[Stab.scala 175:24]
    .clock(last_merger_227_clock),
    .reset(last_merger_227_reset),
    .io_stream1_ready(last_merger_227_io_stream1_ready),
    .io_stream1_valid(last_merger_227_io_stream1_valid),
    .io_stream1_bits(last_merger_227_io_stream1_bits),
    .io_stream2_ready(last_merger_227_io_stream2_ready),
    .io_stream2_valid(last_merger_227_io_stream2_valid),
    .io_stream2_bits(last_merger_227_io_stream2_bits),
    .io_result_ready(last_merger_227_io_result_ready),
    .io_result_valid(last_merger_227_io_result_valid),
    .io_result_bits(last_merger_227_io_result_bits)
  );
  Queue last_q_227 ( // @[Decoupled.scala 361:21]
    .clock(last_q_227_clock),
    .reset(last_q_227_reset),
    .io_enq_ready(last_q_227_io_enq_ready),
    .io_enq_valid(last_q_227_io_enq_valid),
    .io_enq_bits(last_q_227_io_enq_bits),
    .io_deq_ready(last_q_227_io_deq_ready),
    .io_deq_valid(last_q_227_io_deq_valid),
    .io_deq_bits(last_q_227_io_deq_bits)
  );
  StreamMerger_228 last_merger_228 ( // @[Stab.scala 175:24]
    .clock(last_merger_228_clock),
    .reset(last_merger_228_reset),
    .io_stream1_ready(last_merger_228_io_stream1_ready),
    .io_stream1_valid(last_merger_228_io_stream1_valid),
    .io_stream1_bits(last_merger_228_io_stream1_bits),
    .io_stream2_ready(last_merger_228_io_stream2_ready),
    .io_stream2_valid(last_merger_228_io_stream2_valid),
    .io_stream2_bits(last_merger_228_io_stream2_bits),
    .io_result_ready(last_merger_228_io_result_ready),
    .io_result_valid(last_merger_228_io_result_valid),
    .io_result_bits(last_merger_228_io_result_bits)
  );
  Queue last_q_228 ( // @[Decoupled.scala 361:21]
    .clock(last_q_228_clock),
    .reset(last_q_228_reset),
    .io_enq_ready(last_q_228_io_enq_ready),
    .io_enq_valid(last_q_228_io_enq_valid),
    .io_enq_bits(last_q_228_io_enq_bits),
    .io_deq_ready(last_q_228_io_deq_ready),
    .io_deq_valid(last_q_228_io_deq_valid),
    .io_deq_bits(last_q_228_io_deq_bits)
  );
  StreamMerger_229 last_merger_229 ( // @[Stab.scala 175:24]
    .clock(last_merger_229_clock),
    .reset(last_merger_229_reset),
    .io_stream1_ready(last_merger_229_io_stream1_ready),
    .io_stream1_valid(last_merger_229_io_stream1_valid),
    .io_stream1_bits(last_merger_229_io_stream1_bits),
    .io_stream2_ready(last_merger_229_io_stream2_ready),
    .io_stream2_valid(last_merger_229_io_stream2_valid),
    .io_stream2_bits(last_merger_229_io_stream2_bits),
    .io_result_ready(last_merger_229_io_result_ready),
    .io_result_valid(last_merger_229_io_result_valid),
    .io_result_bits(last_merger_229_io_result_bits)
  );
  Queue last_q_229 ( // @[Decoupled.scala 361:21]
    .clock(last_q_229_clock),
    .reset(last_q_229_reset),
    .io_enq_ready(last_q_229_io_enq_ready),
    .io_enq_valid(last_q_229_io_enq_valid),
    .io_enq_bits(last_q_229_io_enq_bits),
    .io_deq_ready(last_q_229_io_deq_ready),
    .io_deq_valid(last_q_229_io_deq_valid),
    .io_deq_bits(last_q_229_io_deq_bits)
  );
  StreamMerger_230 last_merger_230 ( // @[Stab.scala 175:24]
    .clock(last_merger_230_clock),
    .reset(last_merger_230_reset),
    .io_stream1_ready(last_merger_230_io_stream1_ready),
    .io_stream1_valid(last_merger_230_io_stream1_valid),
    .io_stream1_bits(last_merger_230_io_stream1_bits),
    .io_stream2_ready(last_merger_230_io_stream2_ready),
    .io_stream2_valid(last_merger_230_io_stream2_valid),
    .io_stream2_bits(last_merger_230_io_stream2_bits),
    .io_result_ready(last_merger_230_io_result_ready),
    .io_result_valid(last_merger_230_io_result_valid),
    .io_result_bits(last_merger_230_io_result_bits)
  );
  Queue last_q_230 ( // @[Decoupled.scala 361:21]
    .clock(last_q_230_clock),
    .reset(last_q_230_reset),
    .io_enq_ready(last_q_230_io_enq_ready),
    .io_enq_valid(last_q_230_io_enq_valid),
    .io_enq_bits(last_q_230_io_enq_bits),
    .io_deq_ready(last_q_230_io_deq_ready),
    .io_deq_valid(last_q_230_io_deq_valid),
    .io_deq_bits(last_q_230_io_deq_bits)
  );
  StreamMerger_231 last_merger_231 ( // @[Stab.scala 175:24]
    .clock(last_merger_231_clock),
    .reset(last_merger_231_reset),
    .io_stream1_ready(last_merger_231_io_stream1_ready),
    .io_stream1_valid(last_merger_231_io_stream1_valid),
    .io_stream1_bits(last_merger_231_io_stream1_bits),
    .io_stream2_ready(last_merger_231_io_stream2_ready),
    .io_stream2_valid(last_merger_231_io_stream2_valid),
    .io_stream2_bits(last_merger_231_io_stream2_bits),
    .io_result_ready(last_merger_231_io_result_ready),
    .io_result_valid(last_merger_231_io_result_valid),
    .io_result_bits(last_merger_231_io_result_bits)
  );
  Queue last_q_231 ( // @[Decoupled.scala 361:21]
    .clock(last_q_231_clock),
    .reset(last_q_231_reset),
    .io_enq_ready(last_q_231_io_enq_ready),
    .io_enq_valid(last_q_231_io_enq_valid),
    .io_enq_bits(last_q_231_io_enq_bits),
    .io_deq_ready(last_q_231_io_deq_ready),
    .io_deq_valid(last_q_231_io_deq_valid),
    .io_deq_bits(last_q_231_io_deq_bits)
  );
  StreamMerger_232 last_merger_232 ( // @[Stab.scala 175:24]
    .clock(last_merger_232_clock),
    .reset(last_merger_232_reset),
    .io_stream1_ready(last_merger_232_io_stream1_ready),
    .io_stream1_valid(last_merger_232_io_stream1_valid),
    .io_stream1_bits(last_merger_232_io_stream1_bits),
    .io_stream2_ready(last_merger_232_io_stream2_ready),
    .io_stream2_valid(last_merger_232_io_stream2_valid),
    .io_stream2_bits(last_merger_232_io_stream2_bits),
    .io_result_ready(last_merger_232_io_result_ready),
    .io_result_valid(last_merger_232_io_result_valid),
    .io_result_bits(last_merger_232_io_result_bits)
  );
  Queue last_q_232 ( // @[Decoupled.scala 361:21]
    .clock(last_q_232_clock),
    .reset(last_q_232_reset),
    .io_enq_ready(last_q_232_io_enq_ready),
    .io_enq_valid(last_q_232_io_enq_valid),
    .io_enq_bits(last_q_232_io_enq_bits),
    .io_deq_ready(last_q_232_io_deq_ready),
    .io_deq_valid(last_q_232_io_deq_valid),
    .io_deq_bits(last_q_232_io_deq_bits)
  );
  StreamMerger_233 last_merger_233 ( // @[Stab.scala 175:24]
    .clock(last_merger_233_clock),
    .reset(last_merger_233_reset),
    .io_stream1_ready(last_merger_233_io_stream1_ready),
    .io_stream1_valid(last_merger_233_io_stream1_valid),
    .io_stream1_bits(last_merger_233_io_stream1_bits),
    .io_stream2_ready(last_merger_233_io_stream2_ready),
    .io_stream2_valid(last_merger_233_io_stream2_valid),
    .io_stream2_bits(last_merger_233_io_stream2_bits),
    .io_result_ready(last_merger_233_io_result_ready),
    .io_result_valid(last_merger_233_io_result_valid),
    .io_result_bits(last_merger_233_io_result_bits)
  );
  Queue last_q_233 ( // @[Decoupled.scala 361:21]
    .clock(last_q_233_clock),
    .reset(last_q_233_reset),
    .io_enq_ready(last_q_233_io_enq_ready),
    .io_enq_valid(last_q_233_io_enq_valid),
    .io_enq_bits(last_q_233_io_enq_bits),
    .io_deq_ready(last_q_233_io_deq_ready),
    .io_deq_valid(last_q_233_io_deq_valid),
    .io_deq_bits(last_q_233_io_deq_bits)
  );
  StreamMerger_234 last_merger_234 ( // @[Stab.scala 175:24]
    .clock(last_merger_234_clock),
    .reset(last_merger_234_reset),
    .io_stream1_ready(last_merger_234_io_stream1_ready),
    .io_stream1_valid(last_merger_234_io_stream1_valid),
    .io_stream1_bits(last_merger_234_io_stream1_bits),
    .io_stream2_ready(last_merger_234_io_stream2_ready),
    .io_stream2_valid(last_merger_234_io_stream2_valid),
    .io_stream2_bits(last_merger_234_io_stream2_bits),
    .io_result_ready(last_merger_234_io_result_ready),
    .io_result_valid(last_merger_234_io_result_valid),
    .io_result_bits(last_merger_234_io_result_bits)
  );
  Queue last_q_234 ( // @[Decoupled.scala 361:21]
    .clock(last_q_234_clock),
    .reset(last_q_234_reset),
    .io_enq_ready(last_q_234_io_enq_ready),
    .io_enq_valid(last_q_234_io_enq_valid),
    .io_enq_bits(last_q_234_io_enq_bits),
    .io_deq_ready(last_q_234_io_deq_ready),
    .io_deq_valid(last_q_234_io_deq_valid),
    .io_deq_bits(last_q_234_io_deq_bits)
  );
  StreamMerger_235 last_merger_235 ( // @[Stab.scala 175:24]
    .clock(last_merger_235_clock),
    .reset(last_merger_235_reset),
    .io_stream1_ready(last_merger_235_io_stream1_ready),
    .io_stream1_valid(last_merger_235_io_stream1_valid),
    .io_stream1_bits(last_merger_235_io_stream1_bits),
    .io_stream2_ready(last_merger_235_io_stream2_ready),
    .io_stream2_valid(last_merger_235_io_stream2_valid),
    .io_stream2_bits(last_merger_235_io_stream2_bits),
    .io_result_ready(last_merger_235_io_result_ready),
    .io_result_valid(last_merger_235_io_result_valid),
    .io_result_bits(last_merger_235_io_result_bits)
  );
  Queue last_q_235 ( // @[Decoupled.scala 361:21]
    .clock(last_q_235_clock),
    .reset(last_q_235_reset),
    .io_enq_ready(last_q_235_io_enq_ready),
    .io_enq_valid(last_q_235_io_enq_valid),
    .io_enq_bits(last_q_235_io_enq_bits),
    .io_deq_ready(last_q_235_io_deq_ready),
    .io_deq_valid(last_q_235_io_deq_valid),
    .io_deq_bits(last_q_235_io_deq_bits)
  );
  StreamMerger_236 last_merger_236 ( // @[Stab.scala 175:24]
    .clock(last_merger_236_clock),
    .reset(last_merger_236_reset),
    .io_stream1_ready(last_merger_236_io_stream1_ready),
    .io_stream1_valid(last_merger_236_io_stream1_valid),
    .io_stream1_bits(last_merger_236_io_stream1_bits),
    .io_stream2_ready(last_merger_236_io_stream2_ready),
    .io_stream2_valid(last_merger_236_io_stream2_valid),
    .io_stream2_bits(last_merger_236_io_stream2_bits),
    .io_result_ready(last_merger_236_io_result_ready),
    .io_result_valid(last_merger_236_io_result_valid),
    .io_result_bits(last_merger_236_io_result_bits)
  );
  Queue last_q_236 ( // @[Decoupled.scala 361:21]
    .clock(last_q_236_clock),
    .reset(last_q_236_reset),
    .io_enq_ready(last_q_236_io_enq_ready),
    .io_enq_valid(last_q_236_io_enq_valid),
    .io_enq_bits(last_q_236_io_enq_bits),
    .io_deq_ready(last_q_236_io_deq_ready),
    .io_deq_valid(last_q_236_io_deq_valid),
    .io_deq_bits(last_q_236_io_deq_bits)
  );
  StreamMerger_237 last_merger_237 ( // @[Stab.scala 175:24]
    .clock(last_merger_237_clock),
    .reset(last_merger_237_reset),
    .io_stream1_ready(last_merger_237_io_stream1_ready),
    .io_stream1_valid(last_merger_237_io_stream1_valid),
    .io_stream1_bits(last_merger_237_io_stream1_bits),
    .io_stream2_ready(last_merger_237_io_stream2_ready),
    .io_stream2_valid(last_merger_237_io_stream2_valid),
    .io_stream2_bits(last_merger_237_io_stream2_bits),
    .io_result_ready(last_merger_237_io_result_ready),
    .io_result_valid(last_merger_237_io_result_valid),
    .io_result_bits(last_merger_237_io_result_bits)
  );
  Queue last_q_237 ( // @[Decoupled.scala 361:21]
    .clock(last_q_237_clock),
    .reset(last_q_237_reset),
    .io_enq_ready(last_q_237_io_enq_ready),
    .io_enq_valid(last_q_237_io_enq_valid),
    .io_enq_bits(last_q_237_io_enq_bits),
    .io_deq_ready(last_q_237_io_deq_ready),
    .io_deq_valid(last_q_237_io_deq_valid),
    .io_deq_bits(last_q_237_io_deq_bits)
  );
  StreamMerger_238 last_merger_238 ( // @[Stab.scala 175:24]
    .clock(last_merger_238_clock),
    .reset(last_merger_238_reset),
    .io_stream1_ready(last_merger_238_io_stream1_ready),
    .io_stream1_valid(last_merger_238_io_stream1_valid),
    .io_stream1_bits(last_merger_238_io_stream1_bits),
    .io_stream2_ready(last_merger_238_io_stream2_ready),
    .io_stream2_valid(last_merger_238_io_stream2_valid),
    .io_stream2_bits(last_merger_238_io_stream2_bits),
    .io_result_ready(last_merger_238_io_result_ready),
    .io_result_valid(last_merger_238_io_result_valid),
    .io_result_bits(last_merger_238_io_result_bits)
  );
  Queue last_q_238 ( // @[Decoupled.scala 361:21]
    .clock(last_q_238_clock),
    .reset(last_q_238_reset),
    .io_enq_ready(last_q_238_io_enq_ready),
    .io_enq_valid(last_q_238_io_enq_valid),
    .io_enq_bits(last_q_238_io_enq_bits),
    .io_deq_ready(last_q_238_io_deq_ready),
    .io_deq_valid(last_q_238_io_deq_valid),
    .io_deq_bits(last_q_238_io_deq_bits)
  );
  StreamMerger_239 last_merger_239 ( // @[Stab.scala 175:24]
    .clock(last_merger_239_clock),
    .reset(last_merger_239_reset),
    .io_stream1_ready(last_merger_239_io_stream1_ready),
    .io_stream1_valid(last_merger_239_io_stream1_valid),
    .io_stream1_bits(last_merger_239_io_stream1_bits),
    .io_stream2_ready(last_merger_239_io_stream2_ready),
    .io_stream2_valid(last_merger_239_io_stream2_valid),
    .io_stream2_bits(last_merger_239_io_stream2_bits),
    .io_result_ready(last_merger_239_io_result_ready),
    .io_result_valid(last_merger_239_io_result_valid),
    .io_result_bits(last_merger_239_io_result_bits)
  );
  Queue last_q_239 ( // @[Decoupled.scala 361:21]
    .clock(last_q_239_clock),
    .reset(last_q_239_reset),
    .io_enq_ready(last_q_239_io_enq_ready),
    .io_enq_valid(last_q_239_io_enq_valid),
    .io_enq_bits(last_q_239_io_enq_bits),
    .io_deq_ready(last_q_239_io_deq_ready),
    .io_deq_valid(last_q_239_io_deq_valid),
    .io_deq_bits(last_q_239_io_deq_bits)
  );
  StreamMerger_240 last_merger_240 ( // @[Stab.scala 175:24]
    .clock(last_merger_240_clock),
    .reset(last_merger_240_reset),
    .io_stream1_ready(last_merger_240_io_stream1_ready),
    .io_stream1_valid(last_merger_240_io_stream1_valid),
    .io_stream1_bits(last_merger_240_io_stream1_bits),
    .io_stream2_ready(last_merger_240_io_stream2_ready),
    .io_stream2_valid(last_merger_240_io_stream2_valid),
    .io_stream2_bits(last_merger_240_io_stream2_bits),
    .io_result_ready(last_merger_240_io_result_ready),
    .io_result_valid(last_merger_240_io_result_valid),
    .io_result_bits(last_merger_240_io_result_bits)
  );
  Queue last_q_240 ( // @[Decoupled.scala 361:21]
    .clock(last_q_240_clock),
    .reset(last_q_240_reset),
    .io_enq_ready(last_q_240_io_enq_ready),
    .io_enq_valid(last_q_240_io_enq_valid),
    .io_enq_bits(last_q_240_io_enq_bits),
    .io_deq_ready(last_q_240_io_deq_ready),
    .io_deq_valid(last_q_240_io_deq_valid),
    .io_deq_bits(last_q_240_io_deq_bits)
  );
  StreamMerger_241 last_merger_241 ( // @[Stab.scala 175:24]
    .clock(last_merger_241_clock),
    .reset(last_merger_241_reset),
    .io_stream1_ready(last_merger_241_io_stream1_ready),
    .io_stream1_valid(last_merger_241_io_stream1_valid),
    .io_stream1_bits(last_merger_241_io_stream1_bits),
    .io_stream2_ready(last_merger_241_io_stream2_ready),
    .io_stream2_valid(last_merger_241_io_stream2_valid),
    .io_stream2_bits(last_merger_241_io_stream2_bits),
    .io_result_ready(last_merger_241_io_result_ready),
    .io_result_valid(last_merger_241_io_result_valid),
    .io_result_bits(last_merger_241_io_result_bits)
  );
  Queue last_q_241 ( // @[Decoupled.scala 361:21]
    .clock(last_q_241_clock),
    .reset(last_q_241_reset),
    .io_enq_ready(last_q_241_io_enq_ready),
    .io_enq_valid(last_q_241_io_enq_valid),
    .io_enq_bits(last_q_241_io_enq_bits),
    .io_deq_ready(last_q_241_io_deq_ready),
    .io_deq_valid(last_q_241_io_deq_valid),
    .io_deq_bits(last_q_241_io_deq_bits)
  );
  StreamMerger_242 last_merger_242 ( // @[Stab.scala 175:24]
    .clock(last_merger_242_clock),
    .reset(last_merger_242_reset),
    .io_stream1_ready(last_merger_242_io_stream1_ready),
    .io_stream1_valid(last_merger_242_io_stream1_valid),
    .io_stream1_bits(last_merger_242_io_stream1_bits),
    .io_stream2_ready(last_merger_242_io_stream2_ready),
    .io_stream2_valid(last_merger_242_io_stream2_valid),
    .io_stream2_bits(last_merger_242_io_stream2_bits),
    .io_result_ready(last_merger_242_io_result_ready),
    .io_result_valid(last_merger_242_io_result_valid),
    .io_result_bits(last_merger_242_io_result_bits)
  );
  Queue last_q_242 ( // @[Decoupled.scala 361:21]
    .clock(last_q_242_clock),
    .reset(last_q_242_reset),
    .io_enq_ready(last_q_242_io_enq_ready),
    .io_enq_valid(last_q_242_io_enq_valid),
    .io_enq_bits(last_q_242_io_enq_bits),
    .io_deq_ready(last_q_242_io_deq_ready),
    .io_deq_valid(last_q_242_io_deq_valid),
    .io_deq_bits(last_q_242_io_deq_bits)
  );
  StreamMerger_243 last_merger_243 ( // @[Stab.scala 175:24]
    .clock(last_merger_243_clock),
    .reset(last_merger_243_reset),
    .io_stream1_ready(last_merger_243_io_stream1_ready),
    .io_stream1_valid(last_merger_243_io_stream1_valid),
    .io_stream1_bits(last_merger_243_io_stream1_bits),
    .io_stream2_ready(last_merger_243_io_stream2_ready),
    .io_stream2_valid(last_merger_243_io_stream2_valid),
    .io_stream2_bits(last_merger_243_io_stream2_bits),
    .io_result_ready(last_merger_243_io_result_ready),
    .io_result_valid(last_merger_243_io_result_valid),
    .io_result_bits(last_merger_243_io_result_bits)
  );
  Queue last_q_243 ( // @[Decoupled.scala 361:21]
    .clock(last_q_243_clock),
    .reset(last_q_243_reset),
    .io_enq_ready(last_q_243_io_enq_ready),
    .io_enq_valid(last_q_243_io_enq_valid),
    .io_enq_bits(last_q_243_io_enq_bits),
    .io_deq_ready(last_q_243_io_deq_ready),
    .io_deq_valid(last_q_243_io_deq_valid),
    .io_deq_bits(last_q_243_io_deq_bits)
  );
  StreamMerger_244 last_merger_244 ( // @[Stab.scala 175:24]
    .clock(last_merger_244_clock),
    .reset(last_merger_244_reset),
    .io_stream1_ready(last_merger_244_io_stream1_ready),
    .io_stream1_valid(last_merger_244_io_stream1_valid),
    .io_stream1_bits(last_merger_244_io_stream1_bits),
    .io_stream2_ready(last_merger_244_io_stream2_ready),
    .io_stream2_valid(last_merger_244_io_stream2_valid),
    .io_stream2_bits(last_merger_244_io_stream2_bits),
    .io_result_ready(last_merger_244_io_result_ready),
    .io_result_valid(last_merger_244_io_result_valid),
    .io_result_bits(last_merger_244_io_result_bits)
  );
  Queue last_q_244 ( // @[Decoupled.scala 361:21]
    .clock(last_q_244_clock),
    .reset(last_q_244_reset),
    .io_enq_ready(last_q_244_io_enq_ready),
    .io_enq_valid(last_q_244_io_enq_valid),
    .io_enq_bits(last_q_244_io_enq_bits),
    .io_deq_ready(last_q_244_io_deq_ready),
    .io_deq_valid(last_q_244_io_deq_valid),
    .io_deq_bits(last_q_244_io_deq_bits)
  );
  StreamMerger_245 last_merger_245 ( // @[Stab.scala 175:24]
    .clock(last_merger_245_clock),
    .reset(last_merger_245_reset),
    .io_stream1_ready(last_merger_245_io_stream1_ready),
    .io_stream1_valid(last_merger_245_io_stream1_valid),
    .io_stream1_bits(last_merger_245_io_stream1_bits),
    .io_stream2_ready(last_merger_245_io_stream2_ready),
    .io_stream2_valid(last_merger_245_io_stream2_valid),
    .io_stream2_bits(last_merger_245_io_stream2_bits),
    .io_result_ready(last_merger_245_io_result_ready),
    .io_result_valid(last_merger_245_io_result_valid),
    .io_result_bits(last_merger_245_io_result_bits)
  );
  Queue last_q_245 ( // @[Decoupled.scala 361:21]
    .clock(last_q_245_clock),
    .reset(last_q_245_reset),
    .io_enq_ready(last_q_245_io_enq_ready),
    .io_enq_valid(last_q_245_io_enq_valid),
    .io_enq_bits(last_q_245_io_enq_bits),
    .io_deq_ready(last_q_245_io_deq_ready),
    .io_deq_valid(last_q_245_io_deq_valid),
    .io_deq_bits(last_q_245_io_deq_bits)
  );
  StreamMerger_246 last_merger_246 ( // @[Stab.scala 175:24]
    .clock(last_merger_246_clock),
    .reset(last_merger_246_reset),
    .io_stream1_ready(last_merger_246_io_stream1_ready),
    .io_stream1_valid(last_merger_246_io_stream1_valid),
    .io_stream1_bits(last_merger_246_io_stream1_bits),
    .io_stream2_ready(last_merger_246_io_stream2_ready),
    .io_stream2_valid(last_merger_246_io_stream2_valid),
    .io_stream2_bits(last_merger_246_io_stream2_bits),
    .io_result_ready(last_merger_246_io_result_ready),
    .io_result_valid(last_merger_246_io_result_valid),
    .io_result_bits(last_merger_246_io_result_bits)
  );
  Queue last_q_246 ( // @[Decoupled.scala 361:21]
    .clock(last_q_246_clock),
    .reset(last_q_246_reset),
    .io_enq_ready(last_q_246_io_enq_ready),
    .io_enq_valid(last_q_246_io_enq_valid),
    .io_enq_bits(last_q_246_io_enq_bits),
    .io_deq_ready(last_q_246_io_deq_ready),
    .io_deq_valid(last_q_246_io_deq_valid),
    .io_deq_bits(last_q_246_io_deq_bits)
  );
  StreamMerger_247 last_merger_247 ( // @[Stab.scala 175:24]
    .clock(last_merger_247_clock),
    .reset(last_merger_247_reset),
    .io_stream1_ready(last_merger_247_io_stream1_ready),
    .io_stream1_valid(last_merger_247_io_stream1_valid),
    .io_stream1_bits(last_merger_247_io_stream1_bits),
    .io_stream2_ready(last_merger_247_io_stream2_ready),
    .io_stream2_valid(last_merger_247_io_stream2_valid),
    .io_stream2_bits(last_merger_247_io_stream2_bits),
    .io_result_ready(last_merger_247_io_result_ready),
    .io_result_valid(last_merger_247_io_result_valid),
    .io_result_bits(last_merger_247_io_result_bits)
  );
  Queue last_q_247 ( // @[Decoupled.scala 361:21]
    .clock(last_q_247_clock),
    .reset(last_q_247_reset),
    .io_enq_ready(last_q_247_io_enq_ready),
    .io_enq_valid(last_q_247_io_enq_valid),
    .io_enq_bits(last_q_247_io_enq_bits),
    .io_deq_ready(last_q_247_io_deq_ready),
    .io_deq_valid(last_q_247_io_deq_valid),
    .io_deq_bits(last_q_247_io_deq_bits)
  );
  StreamMerger_248 last_merger_248 ( // @[Stab.scala 175:24]
    .clock(last_merger_248_clock),
    .reset(last_merger_248_reset),
    .io_stream1_ready(last_merger_248_io_stream1_ready),
    .io_stream1_valid(last_merger_248_io_stream1_valid),
    .io_stream1_bits(last_merger_248_io_stream1_bits),
    .io_stream2_ready(last_merger_248_io_stream2_ready),
    .io_stream2_valid(last_merger_248_io_stream2_valid),
    .io_stream2_bits(last_merger_248_io_stream2_bits),
    .io_result_ready(last_merger_248_io_result_ready),
    .io_result_valid(last_merger_248_io_result_valid),
    .io_result_bits(last_merger_248_io_result_bits)
  );
  Queue last_q_248 ( // @[Decoupled.scala 361:21]
    .clock(last_q_248_clock),
    .reset(last_q_248_reset),
    .io_enq_ready(last_q_248_io_enq_ready),
    .io_enq_valid(last_q_248_io_enq_valid),
    .io_enq_bits(last_q_248_io_enq_bits),
    .io_deq_ready(last_q_248_io_deq_ready),
    .io_deq_valid(last_q_248_io_deq_valid),
    .io_deq_bits(last_q_248_io_deq_bits)
  );
  StreamMerger_249 last_merger_249 ( // @[Stab.scala 175:24]
    .clock(last_merger_249_clock),
    .reset(last_merger_249_reset),
    .io_stream1_ready(last_merger_249_io_stream1_ready),
    .io_stream1_valid(last_merger_249_io_stream1_valid),
    .io_stream1_bits(last_merger_249_io_stream1_bits),
    .io_stream2_ready(last_merger_249_io_stream2_ready),
    .io_stream2_valid(last_merger_249_io_stream2_valid),
    .io_stream2_bits(last_merger_249_io_stream2_bits),
    .io_result_ready(last_merger_249_io_result_ready),
    .io_result_valid(last_merger_249_io_result_valid),
    .io_result_bits(last_merger_249_io_result_bits)
  );
  Queue last_q_249 ( // @[Decoupled.scala 361:21]
    .clock(last_q_249_clock),
    .reset(last_q_249_reset),
    .io_enq_ready(last_q_249_io_enq_ready),
    .io_enq_valid(last_q_249_io_enq_valid),
    .io_enq_bits(last_q_249_io_enq_bits),
    .io_deq_ready(last_q_249_io_deq_ready),
    .io_deq_valid(last_q_249_io_deq_valid),
    .io_deq_bits(last_q_249_io_deq_bits)
  );
  StreamMerger_250 last_merger_250 ( // @[Stab.scala 175:24]
    .clock(last_merger_250_clock),
    .reset(last_merger_250_reset),
    .io_stream1_ready(last_merger_250_io_stream1_ready),
    .io_stream1_valid(last_merger_250_io_stream1_valid),
    .io_stream1_bits(last_merger_250_io_stream1_bits),
    .io_stream2_ready(last_merger_250_io_stream2_ready),
    .io_stream2_valid(last_merger_250_io_stream2_valid),
    .io_stream2_bits(last_merger_250_io_stream2_bits),
    .io_result_ready(last_merger_250_io_result_ready),
    .io_result_valid(last_merger_250_io_result_valid),
    .io_result_bits(last_merger_250_io_result_bits)
  );
  Queue last_q_250 ( // @[Decoupled.scala 361:21]
    .clock(last_q_250_clock),
    .reset(last_q_250_reset),
    .io_enq_ready(last_q_250_io_enq_ready),
    .io_enq_valid(last_q_250_io_enq_valid),
    .io_enq_bits(last_q_250_io_enq_bits),
    .io_deq_ready(last_q_250_io_deq_ready),
    .io_deq_valid(last_q_250_io_deq_valid),
    .io_deq_bits(last_q_250_io_deq_bits)
  );
  StreamMerger_251 last_merger_251 ( // @[Stab.scala 175:24]
    .clock(last_merger_251_clock),
    .reset(last_merger_251_reset),
    .io_stream1_ready(last_merger_251_io_stream1_ready),
    .io_stream1_valid(last_merger_251_io_stream1_valid),
    .io_stream1_bits(last_merger_251_io_stream1_bits),
    .io_stream2_ready(last_merger_251_io_stream2_ready),
    .io_stream2_valid(last_merger_251_io_stream2_valid),
    .io_stream2_bits(last_merger_251_io_stream2_bits),
    .io_result_ready(last_merger_251_io_result_ready),
    .io_result_valid(last_merger_251_io_result_valid),
    .io_result_bits(last_merger_251_io_result_bits)
  );
  Queue last_q_251 ( // @[Decoupled.scala 361:21]
    .clock(last_q_251_clock),
    .reset(last_q_251_reset),
    .io_enq_ready(last_q_251_io_enq_ready),
    .io_enq_valid(last_q_251_io_enq_valid),
    .io_enq_bits(last_q_251_io_enq_bits),
    .io_deq_ready(last_q_251_io_deq_ready),
    .io_deq_valid(last_q_251_io_deq_valid),
    .io_deq_bits(last_q_251_io_deq_bits)
  );
  StreamMerger_252 last_merger_252 ( // @[Stab.scala 175:24]
    .clock(last_merger_252_clock),
    .reset(last_merger_252_reset),
    .io_stream1_ready(last_merger_252_io_stream1_ready),
    .io_stream1_valid(last_merger_252_io_stream1_valid),
    .io_stream1_bits(last_merger_252_io_stream1_bits),
    .io_stream2_ready(last_merger_252_io_stream2_ready),
    .io_stream2_valid(last_merger_252_io_stream2_valid),
    .io_stream2_bits(last_merger_252_io_stream2_bits),
    .io_result_ready(last_merger_252_io_result_ready),
    .io_result_valid(last_merger_252_io_result_valid),
    .io_result_bits(last_merger_252_io_result_bits)
  );
  Queue last_q_252 ( // @[Decoupled.scala 361:21]
    .clock(last_q_252_clock),
    .reset(last_q_252_reset),
    .io_enq_ready(last_q_252_io_enq_ready),
    .io_enq_valid(last_q_252_io_enq_valid),
    .io_enq_bits(last_q_252_io_enq_bits),
    .io_deq_ready(last_q_252_io_deq_ready),
    .io_deq_valid(last_q_252_io_deq_valid),
    .io_deq_bits(last_q_252_io_deq_bits)
  );
  StreamMerger_253 last_merger_253 ( // @[Stab.scala 175:24]
    .clock(last_merger_253_clock),
    .reset(last_merger_253_reset),
    .io_stream1_ready(last_merger_253_io_stream1_ready),
    .io_stream1_valid(last_merger_253_io_stream1_valid),
    .io_stream1_bits(last_merger_253_io_stream1_bits),
    .io_stream2_ready(last_merger_253_io_stream2_ready),
    .io_stream2_valid(last_merger_253_io_stream2_valid),
    .io_stream2_bits(last_merger_253_io_stream2_bits),
    .io_result_ready(last_merger_253_io_result_ready),
    .io_result_valid(last_merger_253_io_result_valid),
    .io_result_bits(last_merger_253_io_result_bits)
  );
  Queue last_q_253 ( // @[Decoupled.scala 361:21]
    .clock(last_q_253_clock),
    .reset(last_q_253_reset),
    .io_enq_ready(last_q_253_io_enq_ready),
    .io_enq_valid(last_q_253_io_enq_valid),
    .io_enq_bits(last_q_253_io_enq_bits),
    .io_deq_ready(last_q_253_io_deq_ready),
    .io_deq_valid(last_q_253_io_deq_valid),
    .io_deq_bits(last_q_253_io_deq_bits)
  );
  StreamMerger_254 last_merger_254 ( // @[Stab.scala 175:24]
    .clock(last_merger_254_clock),
    .reset(last_merger_254_reset),
    .io_stream1_ready(last_merger_254_io_stream1_ready),
    .io_stream1_valid(last_merger_254_io_stream1_valid),
    .io_stream1_bits(last_merger_254_io_stream1_bits),
    .io_stream2_ready(last_merger_254_io_stream2_ready),
    .io_stream2_valid(last_merger_254_io_stream2_valid),
    .io_stream2_bits(last_merger_254_io_stream2_bits),
    .io_result_ready(last_merger_254_io_result_ready),
    .io_result_valid(last_merger_254_io_result_valid),
    .io_result_bits(last_merger_254_io_result_bits)
  );
  Queue last ( // @[Decoupled.scala 361:21]
    .clock(last_clock),
    .reset(last_reset),
    .io_enq_ready(last_io_enq_ready),
    .io_enq_valid(last_io_enq_valid),
    .io_enq_bits(last_io_enq_bits),
    .io_deq_ready(last_io_deq_ready),
    .io_deq_valid(last_io_deq_valid),
    .io_deq_bits(last_io_deq_bits)
  );
  assign io_stream_in_0_ready = last_merger_io_stream1_ready; // @[Stab.scala 176:23]
  assign io_stream_in_1_ready = last_merger_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_2_ready = last_merger_1_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_3_ready = last_merger_2_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_4_ready = last_merger_3_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_5_ready = last_merger_4_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_6_ready = last_merger_5_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_7_ready = last_merger_6_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_8_ready = last_merger_7_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_9_ready = last_merger_8_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_10_ready = last_merger_9_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_11_ready = last_merger_10_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_12_ready = last_merger_11_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_13_ready = last_merger_12_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_14_ready = last_merger_13_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_15_ready = last_merger_14_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_16_ready = last_merger_15_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_17_ready = last_merger_16_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_18_ready = last_merger_17_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_19_ready = last_merger_18_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_20_ready = last_merger_19_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_21_ready = last_merger_20_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_22_ready = last_merger_21_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_23_ready = last_merger_22_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_24_ready = last_merger_23_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_25_ready = last_merger_24_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_26_ready = last_merger_25_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_27_ready = last_merger_26_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_28_ready = last_merger_27_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_29_ready = last_merger_28_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_30_ready = last_merger_29_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_31_ready = last_merger_30_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_32_ready = last_merger_31_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_33_ready = last_merger_32_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_34_ready = last_merger_33_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_35_ready = last_merger_34_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_36_ready = last_merger_35_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_37_ready = last_merger_36_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_38_ready = last_merger_37_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_39_ready = last_merger_38_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_40_ready = last_merger_39_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_41_ready = last_merger_40_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_42_ready = last_merger_41_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_43_ready = last_merger_42_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_44_ready = last_merger_43_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_45_ready = last_merger_44_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_46_ready = last_merger_45_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_47_ready = last_merger_46_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_48_ready = last_merger_47_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_49_ready = last_merger_48_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_50_ready = last_merger_49_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_51_ready = last_merger_50_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_52_ready = last_merger_51_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_53_ready = last_merger_52_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_54_ready = last_merger_53_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_55_ready = last_merger_54_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_56_ready = last_merger_55_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_57_ready = last_merger_56_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_58_ready = last_merger_57_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_59_ready = last_merger_58_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_60_ready = last_merger_59_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_61_ready = last_merger_60_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_62_ready = last_merger_61_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_63_ready = last_merger_62_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_64_ready = last_merger_63_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_65_ready = last_merger_64_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_66_ready = last_merger_65_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_67_ready = last_merger_66_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_68_ready = last_merger_67_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_69_ready = last_merger_68_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_70_ready = last_merger_69_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_71_ready = last_merger_70_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_72_ready = last_merger_71_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_73_ready = last_merger_72_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_74_ready = last_merger_73_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_75_ready = last_merger_74_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_76_ready = last_merger_75_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_77_ready = last_merger_76_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_78_ready = last_merger_77_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_79_ready = last_merger_78_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_80_ready = last_merger_79_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_81_ready = last_merger_80_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_82_ready = last_merger_81_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_83_ready = last_merger_82_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_84_ready = last_merger_83_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_85_ready = last_merger_84_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_86_ready = last_merger_85_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_87_ready = last_merger_86_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_88_ready = last_merger_87_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_89_ready = last_merger_88_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_90_ready = last_merger_89_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_91_ready = last_merger_90_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_92_ready = last_merger_91_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_93_ready = last_merger_92_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_94_ready = last_merger_93_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_95_ready = last_merger_94_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_96_ready = last_merger_95_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_97_ready = last_merger_96_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_98_ready = last_merger_97_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_99_ready = last_merger_98_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_100_ready = last_merger_99_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_101_ready = last_merger_100_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_102_ready = last_merger_101_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_103_ready = last_merger_102_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_104_ready = last_merger_103_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_105_ready = last_merger_104_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_106_ready = last_merger_105_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_107_ready = last_merger_106_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_108_ready = last_merger_107_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_109_ready = last_merger_108_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_110_ready = last_merger_109_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_111_ready = last_merger_110_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_112_ready = last_merger_111_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_113_ready = last_merger_112_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_114_ready = last_merger_113_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_115_ready = last_merger_114_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_116_ready = last_merger_115_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_117_ready = last_merger_116_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_118_ready = last_merger_117_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_119_ready = last_merger_118_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_120_ready = last_merger_119_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_121_ready = last_merger_120_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_122_ready = last_merger_121_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_123_ready = last_merger_122_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_124_ready = last_merger_123_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_125_ready = last_merger_124_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_126_ready = last_merger_125_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_127_ready = last_merger_126_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_128_ready = last_merger_127_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_129_ready = last_merger_128_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_130_ready = last_merger_129_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_131_ready = last_merger_130_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_132_ready = last_merger_131_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_133_ready = last_merger_132_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_134_ready = last_merger_133_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_135_ready = last_merger_134_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_136_ready = last_merger_135_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_137_ready = last_merger_136_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_138_ready = last_merger_137_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_139_ready = last_merger_138_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_140_ready = last_merger_139_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_141_ready = last_merger_140_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_142_ready = last_merger_141_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_143_ready = last_merger_142_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_144_ready = last_merger_143_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_145_ready = last_merger_144_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_146_ready = last_merger_145_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_147_ready = last_merger_146_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_148_ready = last_merger_147_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_149_ready = last_merger_148_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_150_ready = last_merger_149_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_151_ready = last_merger_150_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_152_ready = last_merger_151_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_153_ready = last_merger_152_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_154_ready = last_merger_153_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_155_ready = last_merger_154_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_156_ready = last_merger_155_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_157_ready = last_merger_156_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_158_ready = last_merger_157_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_159_ready = last_merger_158_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_160_ready = last_merger_159_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_161_ready = last_merger_160_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_162_ready = last_merger_161_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_163_ready = last_merger_162_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_164_ready = last_merger_163_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_165_ready = last_merger_164_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_166_ready = last_merger_165_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_167_ready = last_merger_166_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_168_ready = last_merger_167_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_169_ready = last_merger_168_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_170_ready = last_merger_169_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_171_ready = last_merger_170_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_172_ready = last_merger_171_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_173_ready = last_merger_172_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_174_ready = last_merger_173_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_175_ready = last_merger_174_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_176_ready = last_merger_175_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_177_ready = last_merger_176_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_178_ready = last_merger_177_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_179_ready = last_merger_178_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_180_ready = last_merger_179_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_181_ready = last_merger_180_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_182_ready = last_merger_181_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_183_ready = last_merger_182_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_184_ready = last_merger_183_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_185_ready = last_merger_184_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_186_ready = last_merger_185_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_187_ready = last_merger_186_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_188_ready = last_merger_187_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_189_ready = last_merger_188_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_190_ready = last_merger_189_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_191_ready = last_merger_190_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_192_ready = last_merger_191_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_193_ready = last_merger_192_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_194_ready = last_merger_193_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_195_ready = last_merger_194_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_196_ready = last_merger_195_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_197_ready = last_merger_196_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_198_ready = last_merger_197_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_199_ready = last_merger_198_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_200_ready = last_merger_199_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_201_ready = last_merger_200_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_202_ready = last_merger_201_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_203_ready = last_merger_202_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_204_ready = last_merger_203_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_205_ready = last_merger_204_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_206_ready = last_merger_205_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_207_ready = last_merger_206_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_208_ready = last_merger_207_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_209_ready = last_merger_208_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_210_ready = last_merger_209_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_211_ready = last_merger_210_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_212_ready = last_merger_211_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_213_ready = last_merger_212_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_214_ready = last_merger_213_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_215_ready = last_merger_214_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_216_ready = last_merger_215_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_217_ready = last_merger_216_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_218_ready = last_merger_217_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_219_ready = last_merger_218_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_220_ready = last_merger_219_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_221_ready = last_merger_220_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_222_ready = last_merger_221_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_223_ready = last_merger_222_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_224_ready = last_merger_223_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_225_ready = last_merger_224_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_226_ready = last_merger_225_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_227_ready = last_merger_226_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_228_ready = last_merger_227_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_229_ready = last_merger_228_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_230_ready = last_merger_229_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_231_ready = last_merger_230_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_232_ready = last_merger_231_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_233_ready = last_merger_232_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_234_ready = last_merger_233_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_235_ready = last_merger_234_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_236_ready = last_merger_235_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_237_ready = last_merger_236_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_238_ready = last_merger_237_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_239_ready = last_merger_238_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_240_ready = last_merger_239_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_241_ready = last_merger_240_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_242_ready = last_merger_241_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_243_ready = last_merger_242_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_244_ready = last_merger_243_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_245_ready = last_merger_244_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_246_ready = last_merger_245_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_247_ready = last_merger_246_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_248_ready = last_merger_247_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_249_ready = last_merger_248_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_250_ready = last_merger_249_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_251_ready = last_merger_250_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_252_ready = last_merger_251_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_253_ready = last_merger_252_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_254_ready = last_merger_253_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_in_255_ready = last_merger_254_io_stream2_ready; // @[Stab.scala 177:23]
  assign io_stream_out_valid = last_io_deq_valid; // @[Stab.scala 180:17]
  assign io_stream_out_bits = last_io_deq_bits; // @[Stab.scala 180:17]
  assign last_merger_clock = clock;
  assign last_merger_reset = reset;
  assign last_merger_io_stream1_valid = io_stream_in_0_valid; // @[Stab.scala 176:23]
  assign last_merger_io_stream1_bits = io_stream_in_0_bits; // @[Stab.scala 176:23]
  assign last_merger_io_stream2_valid = io_stream_in_1_valid; // @[Stab.scala 177:23]
  assign last_merger_io_stream2_bits = io_stream_in_1_bits; // @[Stab.scala 177:23]
  assign last_merger_io_result_ready = last_q_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_clock = clock;
  assign last_q_reset = reset;
  assign last_q_io_enq_valid = last_merger_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_io_enq_bits = last_merger_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_io_deq_ready = last_merger_1_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_1_clock = clock;
  assign last_merger_1_reset = reset;
  assign last_merger_1_io_stream1_valid = last_q_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_1_io_stream1_bits = last_q_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_1_io_stream2_valid = io_stream_in_2_valid; // @[Stab.scala 177:23]
  assign last_merger_1_io_stream2_bits = io_stream_in_2_bits; // @[Stab.scala 177:23]
  assign last_merger_1_io_result_ready = last_q_1_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_1_clock = clock;
  assign last_q_1_reset = reset;
  assign last_q_1_io_enq_valid = last_merger_1_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_1_io_enq_bits = last_merger_1_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_1_io_deq_ready = last_merger_2_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_2_clock = clock;
  assign last_merger_2_reset = reset;
  assign last_merger_2_io_stream1_valid = last_q_1_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_2_io_stream1_bits = last_q_1_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_2_io_stream2_valid = io_stream_in_3_valid; // @[Stab.scala 177:23]
  assign last_merger_2_io_stream2_bits = io_stream_in_3_bits; // @[Stab.scala 177:23]
  assign last_merger_2_io_result_ready = last_q_2_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_2_clock = clock;
  assign last_q_2_reset = reset;
  assign last_q_2_io_enq_valid = last_merger_2_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_2_io_enq_bits = last_merger_2_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_2_io_deq_ready = last_merger_3_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_3_clock = clock;
  assign last_merger_3_reset = reset;
  assign last_merger_3_io_stream1_valid = last_q_2_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_3_io_stream1_bits = last_q_2_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_3_io_stream2_valid = io_stream_in_4_valid; // @[Stab.scala 177:23]
  assign last_merger_3_io_stream2_bits = io_stream_in_4_bits; // @[Stab.scala 177:23]
  assign last_merger_3_io_result_ready = last_q_3_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_3_clock = clock;
  assign last_q_3_reset = reset;
  assign last_q_3_io_enq_valid = last_merger_3_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_3_io_enq_bits = last_merger_3_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_3_io_deq_ready = last_merger_4_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_4_clock = clock;
  assign last_merger_4_reset = reset;
  assign last_merger_4_io_stream1_valid = last_q_3_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_4_io_stream1_bits = last_q_3_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_4_io_stream2_valid = io_stream_in_5_valid; // @[Stab.scala 177:23]
  assign last_merger_4_io_stream2_bits = io_stream_in_5_bits; // @[Stab.scala 177:23]
  assign last_merger_4_io_result_ready = last_q_4_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_4_clock = clock;
  assign last_q_4_reset = reset;
  assign last_q_4_io_enq_valid = last_merger_4_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_4_io_enq_bits = last_merger_4_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_4_io_deq_ready = last_merger_5_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_5_clock = clock;
  assign last_merger_5_reset = reset;
  assign last_merger_5_io_stream1_valid = last_q_4_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_5_io_stream1_bits = last_q_4_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_5_io_stream2_valid = io_stream_in_6_valid; // @[Stab.scala 177:23]
  assign last_merger_5_io_stream2_bits = io_stream_in_6_bits; // @[Stab.scala 177:23]
  assign last_merger_5_io_result_ready = last_q_5_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_5_clock = clock;
  assign last_q_5_reset = reset;
  assign last_q_5_io_enq_valid = last_merger_5_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_5_io_enq_bits = last_merger_5_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_5_io_deq_ready = last_merger_6_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_6_clock = clock;
  assign last_merger_6_reset = reset;
  assign last_merger_6_io_stream1_valid = last_q_5_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_6_io_stream1_bits = last_q_5_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_6_io_stream2_valid = io_stream_in_7_valid; // @[Stab.scala 177:23]
  assign last_merger_6_io_stream2_bits = io_stream_in_7_bits; // @[Stab.scala 177:23]
  assign last_merger_6_io_result_ready = last_q_6_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_6_clock = clock;
  assign last_q_6_reset = reset;
  assign last_q_6_io_enq_valid = last_merger_6_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_6_io_enq_bits = last_merger_6_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_6_io_deq_ready = last_merger_7_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_7_clock = clock;
  assign last_merger_7_reset = reset;
  assign last_merger_7_io_stream1_valid = last_q_6_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_7_io_stream1_bits = last_q_6_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_7_io_stream2_valid = io_stream_in_8_valid; // @[Stab.scala 177:23]
  assign last_merger_7_io_stream2_bits = io_stream_in_8_bits; // @[Stab.scala 177:23]
  assign last_merger_7_io_result_ready = last_q_7_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_7_clock = clock;
  assign last_q_7_reset = reset;
  assign last_q_7_io_enq_valid = last_merger_7_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_7_io_enq_bits = last_merger_7_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_7_io_deq_ready = last_merger_8_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_8_clock = clock;
  assign last_merger_8_reset = reset;
  assign last_merger_8_io_stream1_valid = last_q_7_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_8_io_stream1_bits = last_q_7_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_8_io_stream2_valid = io_stream_in_9_valid; // @[Stab.scala 177:23]
  assign last_merger_8_io_stream2_bits = io_stream_in_9_bits; // @[Stab.scala 177:23]
  assign last_merger_8_io_result_ready = last_q_8_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_8_clock = clock;
  assign last_q_8_reset = reset;
  assign last_q_8_io_enq_valid = last_merger_8_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_8_io_enq_bits = last_merger_8_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_8_io_deq_ready = last_merger_9_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_9_clock = clock;
  assign last_merger_9_reset = reset;
  assign last_merger_9_io_stream1_valid = last_q_8_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_9_io_stream1_bits = last_q_8_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_9_io_stream2_valid = io_stream_in_10_valid; // @[Stab.scala 177:23]
  assign last_merger_9_io_stream2_bits = io_stream_in_10_bits; // @[Stab.scala 177:23]
  assign last_merger_9_io_result_ready = last_q_9_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_9_clock = clock;
  assign last_q_9_reset = reset;
  assign last_q_9_io_enq_valid = last_merger_9_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_9_io_enq_bits = last_merger_9_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_9_io_deq_ready = last_merger_10_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_10_clock = clock;
  assign last_merger_10_reset = reset;
  assign last_merger_10_io_stream1_valid = last_q_9_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_10_io_stream1_bits = last_q_9_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_10_io_stream2_valid = io_stream_in_11_valid; // @[Stab.scala 177:23]
  assign last_merger_10_io_stream2_bits = io_stream_in_11_bits; // @[Stab.scala 177:23]
  assign last_merger_10_io_result_ready = last_q_10_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_10_clock = clock;
  assign last_q_10_reset = reset;
  assign last_q_10_io_enq_valid = last_merger_10_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_10_io_enq_bits = last_merger_10_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_10_io_deq_ready = last_merger_11_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_11_clock = clock;
  assign last_merger_11_reset = reset;
  assign last_merger_11_io_stream1_valid = last_q_10_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_11_io_stream1_bits = last_q_10_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_11_io_stream2_valid = io_stream_in_12_valid; // @[Stab.scala 177:23]
  assign last_merger_11_io_stream2_bits = io_stream_in_12_bits; // @[Stab.scala 177:23]
  assign last_merger_11_io_result_ready = last_q_11_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_11_clock = clock;
  assign last_q_11_reset = reset;
  assign last_q_11_io_enq_valid = last_merger_11_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_11_io_enq_bits = last_merger_11_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_11_io_deq_ready = last_merger_12_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_12_clock = clock;
  assign last_merger_12_reset = reset;
  assign last_merger_12_io_stream1_valid = last_q_11_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_12_io_stream1_bits = last_q_11_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_12_io_stream2_valid = io_stream_in_13_valid; // @[Stab.scala 177:23]
  assign last_merger_12_io_stream2_bits = io_stream_in_13_bits; // @[Stab.scala 177:23]
  assign last_merger_12_io_result_ready = last_q_12_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_12_clock = clock;
  assign last_q_12_reset = reset;
  assign last_q_12_io_enq_valid = last_merger_12_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_12_io_enq_bits = last_merger_12_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_12_io_deq_ready = last_merger_13_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_13_clock = clock;
  assign last_merger_13_reset = reset;
  assign last_merger_13_io_stream1_valid = last_q_12_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_13_io_stream1_bits = last_q_12_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_13_io_stream2_valid = io_stream_in_14_valid; // @[Stab.scala 177:23]
  assign last_merger_13_io_stream2_bits = io_stream_in_14_bits; // @[Stab.scala 177:23]
  assign last_merger_13_io_result_ready = last_q_13_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_13_clock = clock;
  assign last_q_13_reset = reset;
  assign last_q_13_io_enq_valid = last_merger_13_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_13_io_enq_bits = last_merger_13_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_13_io_deq_ready = last_merger_14_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_14_clock = clock;
  assign last_merger_14_reset = reset;
  assign last_merger_14_io_stream1_valid = last_q_13_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_14_io_stream1_bits = last_q_13_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_14_io_stream2_valid = io_stream_in_15_valid; // @[Stab.scala 177:23]
  assign last_merger_14_io_stream2_bits = io_stream_in_15_bits; // @[Stab.scala 177:23]
  assign last_merger_14_io_result_ready = last_q_14_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_14_clock = clock;
  assign last_q_14_reset = reset;
  assign last_q_14_io_enq_valid = last_merger_14_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_14_io_enq_bits = last_merger_14_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_14_io_deq_ready = last_merger_15_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_15_clock = clock;
  assign last_merger_15_reset = reset;
  assign last_merger_15_io_stream1_valid = last_q_14_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_15_io_stream1_bits = last_q_14_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_15_io_stream2_valid = io_stream_in_16_valid; // @[Stab.scala 177:23]
  assign last_merger_15_io_stream2_bits = io_stream_in_16_bits; // @[Stab.scala 177:23]
  assign last_merger_15_io_result_ready = last_q_15_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_15_clock = clock;
  assign last_q_15_reset = reset;
  assign last_q_15_io_enq_valid = last_merger_15_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_15_io_enq_bits = last_merger_15_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_15_io_deq_ready = last_merger_16_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_16_clock = clock;
  assign last_merger_16_reset = reset;
  assign last_merger_16_io_stream1_valid = last_q_15_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_16_io_stream1_bits = last_q_15_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_16_io_stream2_valid = io_stream_in_17_valid; // @[Stab.scala 177:23]
  assign last_merger_16_io_stream2_bits = io_stream_in_17_bits; // @[Stab.scala 177:23]
  assign last_merger_16_io_result_ready = last_q_16_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_16_clock = clock;
  assign last_q_16_reset = reset;
  assign last_q_16_io_enq_valid = last_merger_16_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_16_io_enq_bits = last_merger_16_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_16_io_deq_ready = last_merger_17_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_17_clock = clock;
  assign last_merger_17_reset = reset;
  assign last_merger_17_io_stream1_valid = last_q_16_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_17_io_stream1_bits = last_q_16_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_17_io_stream2_valid = io_stream_in_18_valid; // @[Stab.scala 177:23]
  assign last_merger_17_io_stream2_bits = io_stream_in_18_bits; // @[Stab.scala 177:23]
  assign last_merger_17_io_result_ready = last_q_17_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_17_clock = clock;
  assign last_q_17_reset = reset;
  assign last_q_17_io_enq_valid = last_merger_17_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_17_io_enq_bits = last_merger_17_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_17_io_deq_ready = last_merger_18_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_18_clock = clock;
  assign last_merger_18_reset = reset;
  assign last_merger_18_io_stream1_valid = last_q_17_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_18_io_stream1_bits = last_q_17_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_18_io_stream2_valid = io_stream_in_19_valid; // @[Stab.scala 177:23]
  assign last_merger_18_io_stream2_bits = io_stream_in_19_bits; // @[Stab.scala 177:23]
  assign last_merger_18_io_result_ready = last_q_18_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_18_clock = clock;
  assign last_q_18_reset = reset;
  assign last_q_18_io_enq_valid = last_merger_18_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_18_io_enq_bits = last_merger_18_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_18_io_deq_ready = last_merger_19_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_19_clock = clock;
  assign last_merger_19_reset = reset;
  assign last_merger_19_io_stream1_valid = last_q_18_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_19_io_stream1_bits = last_q_18_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_19_io_stream2_valid = io_stream_in_20_valid; // @[Stab.scala 177:23]
  assign last_merger_19_io_stream2_bits = io_stream_in_20_bits; // @[Stab.scala 177:23]
  assign last_merger_19_io_result_ready = last_q_19_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_19_clock = clock;
  assign last_q_19_reset = reset;
  assign last_q_19_io_enq_valid = last_merger_19_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_19_io_enq_bits = last_merger_19_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_19_io_deq_ready = last_merger_20_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_20_clock = clock;
  assign last_merger_20_reset = reset;
  assign last_merger_20_io_stream1_valid = last_q_19_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_20_io_stream1_bits = last_q_19_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_20_io_stream2_valid = io_stream_in_21_valid; // @[Stab.scala 177:23]
  assign last_merger_20_io_stream2_bits = io_stream_in_21_bits; // @[Stab.scala 177:23]
  assign last_merger_20_io_result_ready = last_q_20_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_20_clock = clock;
  assign last_q_20_reset = reset;
  assign last_q_20_io_enq_valid = last_merger_20_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_20_io_enq_bits = last_merger_20_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_20_io_deq_ready = last_merger_21_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_21_clock = clock;
  assign last_merger_21_reset = reset;
  assign last_merger_21_io_stream1_valid = last_q_20_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_21_io_stream1_bits = last_q_20_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_21_io_stream2_valid = io_stream_in_22_valid; // @[Stab.scala 177:23]
  assign last_merger_21_io_stream2_bits = io_stream_in_22_bits; // @[Stab.scala 177:23]
  assign last_merger_21_io_result_ready = last_q_21_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_21_clock = clock;
  assign last_q_21_reset = reset;
  assign last_q_21_io_enq_valid = last_merger_21_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_21_io_enq_bits = last_merger_21_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_21_io_deq_ready = last_merger_22_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_22_clock = clock;
  assign last_merger_22_reset = reset;
  assign last_merger_22_io_stream1_valid = last_q_21_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_22_io_stream1_bits = last_q_21_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_22_io_stream2_valid = io_stream_in_23_valid; // @[Stab.scala 177:23]
  assign last_merger_22_io_stream2_bits = io_stream_in_23_bits; // @[Stab.scala 177:23]
  assign last_merger_22_io_result_ready = last_q_22_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_22_clock = clock;
  assign last_q_22_reset = reset;
  assign last_q_22_io_enq_valid = last_merger_22_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_22_io_enq_bits = last_merger_22_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_22_io_deq_ready = last_merger_23_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_23_clock = clock;
  assign last_merger_23_reset = reset;
  assign last_merger_23_io_stream1_valid = last_q_22_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_23_io_stream1_bits = last_q_22_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_23_io_stream2_valid = io_stream_in_24_valid; // @[Stab.scala 177:23]
  assign last_merger_23_io_stream2_bits = io_stream_in_24_bits; // @[Stab.scala 177:23]
  assign last_merger_23_io_result_ready = last_q_23_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_23_clock = clock;
  assign last_q_23_reset = reset;
  assign last_q_23_io_enq_valid = last_merger_23_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_23_io_enq_bits = last_merger_23_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_23_io_deq_ready = last_merger_24_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_24_clock = clock;
  assign last_merger_24_reset = reset;
  assign last_merger_24_io_stream1_valid = last_q_23_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_24_io_stream1_bits = last_q_23_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_24_io_stream2_valid = io_stream_in_25_valid; // @[Stab.scala 177:23]
  assign last_merger_24_io_stream2_bits = io_stream_in_25_bits; // @[Stab.scala 177:23]
  assign last_merger_24_io_result_ready = last_q_24_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_24_clock = clock;
  assign last_q_24_reset = reset;
  assign last_q_24_io_enq_valid = last_merger_24_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_24_io_enq_bits = last_merger_24_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_24_io_deq_ready = last_merger_25_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_25_clock = clock;
  assign last_merger_25_reset = reset;
  assign last_merger_25_io_stream1_valid = last_q_24_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_25_io_stream1_bits = last_q_24_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_25_io_stream2_valid = io_stream_in_26_valid; // @[Stab.scala 177:23]
  assign last_merger_25_io_stream2_bits = io_stream_in_26_bits; // @[Stab.scala 177:23]
  assign last_merger_25_io_result_ready = last_q_25_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_25_clock = clock;
  assign last_q_25_reset = reset;
  assign last_q_25_io_enq_valid = last_merger_25_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_25_io_enq_bits = last_merger_25_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_25_io_deq_ready = last_merger_26_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_26_clock = clock;
  assign last_merger_26_reset = reset;
  assign last_merger_26_io_stream1_valid = last_q_25_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_26_io_stream1_bits = last_q_25_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_26_io_stream2_valid = io_stream_in_27_valid; // @[Stab.scala 177:23]
  assign last_merger_26_io_stream2_bits = io_stream_in_27_bits; // @[Stab.scala 177:23]
  assign last_merger_26_io_result_ready = last_q_26_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_26_clock = clock;
  assign last_q_26_reset = reset;
  assign last_q_26_io_enq_valid = last_merger_26_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_26_io_enq_bits = last_merger_26_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_26_io_deq_ready = last_merger_27_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_27_clock = clock;
  assign last_merger_27_reset = reset;
  assign last_merger_27_io_stream1_valid = last_q_26_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_27_io_stream1_bits = last_q_26_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_27_io_stream2_valid = io_stream_in_28_valid; // @[Stab.scala 177:23]
  assign last_merger_27_io_stream2_bits = io_stream_in_28_bits; // @[Stab.scala 177:23]
  assign last_merger_27_io_result_ready = last_q_27_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_27_clock = clock;
  assign last_q_27_reset = reset;
  assign last_q_27_io_enq_valid = last_merger_27_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_27_io_enq_bits = last_merger_27_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_27_io_deq_ready = last_merger_28_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_28_clock = clock;
  assign last_merger_28_reset = reset;
  assign last_merger_28_io_stream1_valid = last_q_27_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_28_io_stream1_bits = last_q_27_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_28_io_stream2_valid = io_stream_in_29_valid; // @[Stab.scala 177:23]
  assign last_merger_28_io_stream2_bits = io_stream_in_29_bits; // @[Stab.scala 177:23]
  assign last_merger_28_io_result_ready = last_q_28_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_28_clock = clock;
  assign last_q_28_reset = reset;
  assign last_q_28_io_enq_valid = last_merger_28_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_28_io_enq_bits = last_merger_28_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_28_io_deq_ready = last_merger_29_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_29_clock = clock;
  assign last_merger_29_reset = reset;
  assign last_merger_29_io_stream1_valid = last_q_28_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_29_io_stream1_bits = last_q_28_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_29_io_stream2_valid = io_stream_in_30_valid; // @[Stab.scala 177:23]
  assign last_merger_29_io_stream2_bits = io_stream_in_30_bits; // @[Stab.scala 177:23]
  assign last_merger_29_io_result_ready = last_q_29_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_29_clock = clock;
  assign last_q_29_reset = reset;
  assign last_q_29_io_enq_valid = last_merger_29_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_29_io_enq_bits = last_merger_29_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_29_io_deq_ready = last_merger_30_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_30_clock = clock;
  assign last_merger_30_reset = reset;
  assign last_merger_30_io_stream1_valid = last_q_29_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_30_io_stream1_bits = last_q_29_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_30_io_stream2_valid = io_stream_in_31_valid; // @[Stab.scala 177:23]
  assign last_merger_30_io_stream2_bits = io_stream_in_31_bits; // @[Stab.scala 177:23]
  assign last_merger_30_io_result_ready = last_q_30_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_30_clock = clock;
  assign last_q_30_reset = reset;
  assign last_q_30_io_enq_valid = last_merger_30_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_30_io_enq_bits = last_merger_30_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_30_io_deq_ready = last_merger_31_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_31_clock = clock;
  assign last_merger_31_reset = reset;
  assign last_merger_31_io_stream1_valid = last_q_30_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_31_io_stream1_bits = last_q_30_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_31_io_stream2_valid = io_stream_in_32_valid; // @[Stab.scala 177:23]
  assign last_merger_31_io_stream2_bits = io_stream_in_32_bits; // @[Stab.scala 177:23]
  assign last_merger_31_io_result_ready = last_q_31_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_31_clock = clock;
  assign last_q_31_reset = reset;
  assign last_q_31_io_enq_valid = last_merger_31_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_31_io_enq_bits = last_merger_31_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_31_io_deq_ready = last_merger_32_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_32_clock = clock;
  assign last_merger_32_reset = reset;
  assign last_merger_32_io_stream1_valid = last_q_31_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_32_io_stream1_bits = last_q_31_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_32_io_stream2_valid = io_stream_in_33_valid; // @[Stab.scala 177:23]
  assign last_merger_32_io_stream2_bits = io_stream_in_33_bits; // @[Stab.scala 177:23]
  assign last_merger_32_io_result_ready = last_q_32_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_32_clock = clock;
  assign last_q_32_reset = reset;
  assign last_q_32_io_enq_valid = last_merger_32_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_32_io_enq_bits = last_merger_32_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_32_io_deq_ready = last_merger_33_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_33_clock = clock;
  assign last_merger_33_reset = reset;
  assign last_merger_33_io_stream1_valid = last_q_32_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_33_io_stream1_bits = last_q_32_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_33_io_stream2_valid = io_stream_in_34_valid; // @[Stab.scala 177:23]
  assign last_merger_33_io_stream2_bits = io_stream_in_34_bits; // @[Stab.scala 177:23]
  assign last_merger_33_io_result_ready = last_q_33_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_33_clock = clock;
  assign last_q_33_reset = reset;
  assign last_q_33_io_enq_valid = last_merger_33_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_33_io_enq_bits = last_merger_33_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_33_io_deq_ready = last_merger_34_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_34_clock = clock;
  assign last_merger_34_reset = reset;
  assign last_merger_34_io_stream1_valid = last_q_33_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_34_io_stream1_bits = last_q_33_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_34_io_stream2_valid = io_stream_in_35_valid; // @[Stab.scala 177:23]
  assign last_merger_34_io_stream2_bits = io_stream_in_35_bits; // @[Stab.scala 177:23]
  assign last_merger_34_io_result_ready = last_q_34_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_34_clock = clock;
  assign last_q_34_reset = reset;
  assign last_q_34_io_enq_valid = last_merger_34_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_34_io_enq_bits = last_merger_34_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_34_io_deq_ready = last_merger_35_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_35_clock = clock;
  assign last_merger_35_reset = reset;
  assign last_merger_35_io_stream1_valid = last_q_34_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_35_io_stream1_bits = last_q_34_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_35_io_stream2_valid = io_stream_in_36_valid; // @[Stab.scala 177:23]
  assign last_merger_35_io_stream2_bits = io_stream_in_36_bits; // @[Stab.scala 177:23]
  assign last_merger_35_io_result_ready = last_q_35_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_35_clock = clock;
  assign last_q_35_reset = reset;
  assign last_q_35_io_enq_valid = last_merger_35_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_35_io_enq_bits = last_merger_35_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_35_io_deq_ready = last_merger_36_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_36_clock = clock;
  assign last_merger_36_reset = reset;
  assign last_merger_36_io_stream1_valid = last_q_35_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_36_io_stream1_bits = last_q_35_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_36_io_stream2_valid = io_stream_in_37_valid; // @[Stab.scala 177:23]
  assign last_merger_36_io_stream2_bits = io_stream_in_37_bits; // @[Stab.scala 177:23]
  assign last_merger_36_io_result_ready = last_q_36_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_36_clock = clock;
  assign last_q_36_reset = reset;
  assign last_q_36_io_enq_valid = last_merger_36_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_36_io_enq_bits = last_merger_36_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_36_io_deq_ready = last_merger_37_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_37_clock = clock;
  assign last_merger_37_reset = reset;
  assign last_merger_37_io_stream1_valid = last_q_36_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_37_io_stream1_bits = last_q_36_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_37_io_stream2_valid = io_stream_in_38_valid; // @[Stab.scala 177:23]
  assign last_merger_37_io_stream2_bits = io_stream_in_38_bits; // @[Stab.scala 177:23]
  assign last_merger_37_io_result_ready = last_q_37_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_37_clock = clock;
  assign last_q_37_reset = reset;
  assign last_q_37_io_enq_valid = last_merger_37_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_37_io_enq_bits = last_merger_37_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_37_io_deq_ready = last_merger_38_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_38_clock = clock;
  assign last_merger_38_reset = reset;
  assign last_merger_38_io_stream1_valid = last_q_37_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_38_io_stream1_bits = last_q_37_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_38_io_stream2_valid = io_stream_in_39_valid; // @[Stab.scala 177:23]
  assign last_merger_38_io_stream2_bits = io_stream_in_39_bits; // @[Stab.scala 177:23]
  assign last_merger_38_io_result_ready = last_q_38_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_38_clock = clock;
  assign last_q_38_reset = reset;
  assign last_q_38_io_enq_valid = last_merger_38_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_38_io_enq_bits = last_merger_38_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_38_io_deq_ready = last_merger_39_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_39_clock = clock;
  assign last_merger_39_reset = reset;
  assign last_merger_39_io_stream1_valid = last_q_38_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_39_io_stream1_bits = last_q_38_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_39_io_stream2_valid = io_stream_in_40_valid; // @[Stab.scala 177:23]
  assign last_merger_39_io_stream2_bits = io_stream_in_40_bits; // @[Stab.scala 177:23]
  assign last_merger_39_io_result_ready = last_q_39_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_39_clock = clock;
  assign last_q_39_reset = reset;
  assign last_q_39_io_enq_valid = last_merger_39_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_39_io_enq_bits = last_merger_39_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_39_io_deq_ready = last_merger_40_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_40_clock = clock;
  assign last_merger_40_reset = reset;
  assign last_merger_40_io_stream1_valid = last_q_39_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_40_io_stream1_bits = last_q_39_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_40_io_stream2_valid = io_stream_in_41_valid; // @[Stab.scala 177:23]
  assign last_merger_40_io_stream2_bits = io_stream_in_41_bits; // @[Stab.scala 177:23]
  assign last_merger_40_io_result_ready = last_q_40_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_40_clock = clock;
  assign last_q_40_reset = reset;
  assign last_q_40_io_enq_valid = last_merger_40_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_40_io_enq_bits = last_merger_40_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_40_io_deq_ready = last_merger_41_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_41_clock = clock;
  assign last_merger_41_reset = reset;
  assign last_merger_41_io_stream1_valid = last_q_40_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_41_io_stream1_bits = last_q_40_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_41_io_stream2_valid = io_stream_in_42_valid; // @[Stab.scala 177:23]
  assign last_merger_41_io_stream2_bits = io_stream_in_42_bits; // @[Stab.scala 177:23]
  assign last_merger_41_io_result_ready = last_q_41_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_41_clock = clock;
  assign last_q_41_reset = reset;
  assign last_q_41_io_enq_valid = last_merger_41_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_41_io_enq_bits = last_merger_41_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_41_io_deq_ready = last_merger_42_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_42_clock = clock;
  assign last_merger_42_reset = reset;
  assign last_merger_42_io_stream1_valid = last_q_41_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_42_io_stream1_bits = last_q_41_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_42_io_stream2_valid = io_stream_in_43_valid; // @[Stab.scala 177:23]
  assign last_merger_42_io_stream2_bits = io_stream_in_43_bits; // @[Stab.scala 177:23]
  assign last_merger_42_io_result_ready = last_q_42_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_42_clock = clock;
  assign last_q_42_reset = reset;
  assign last_q_42_io_enq_valid = last_merger_42_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_42_io_enq_bits = last_merger_42_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_42_io_deq_ready = last_merger_43_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_43_clock = clock;
  assign last_merger_43_reset = reset;
  assign last_merger_43_io_stream1_valid = last_q_42_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_43_io_stream1_bits = last_q_42_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_43_io_stream2_valid = io_stream_in_44_valid; // @[Stab.scala 177:23]
  assign last_merger_43_io_stream2_bits = io_stream_in_44_bits; // @[Stab.scala 177:23]
  assign last_merger_43_io_result_ready = last_q_43_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_43_clock = clock;
  assign last_q_43_reset = reset;
  assign last_q_43_io_enq_valid = last_merger_43_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_43_io_enq_bits = last_merger_43_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_43_io_deq_ready = last_merger_44_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_44_clock = clock;
  assign last_merger_44_reset = reset;
  assign last_merger_44_io_stream1_valid = last_q_43_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_44_io_stream1_bits = last_q_43_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_44_io_stream2_valid = io_stream_in_45_valid; // @[Stab.scala 177:23]
  assign last_merger_44_io_stream2_bits = io_stream_in_45_bits; // @[Stab.scala 177:23]
  assign last_merger_44_io_result_ready = last_q_44_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_44_clock = clock;
  assign last_q_44_reset = reset;
  assign last_q_44_io_enq_valid = last_merger_44_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_44_io_enq_bits = last_merger_44_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_44_io_deq_ready = last_merger_45_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_45_clock = clock;
  assign last_merger_45_reset = reset;
  assign last_merger_45_io_stream1_valid = last_q_44_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_45_io_stream1_bits = last_q_44_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_45_io_stream2_valid = io_stream_in_46_valid; // @[Stab.scala 177:23]
  assign last_merger_45_io_stream2_bits = io_stream_in_46_bits; // @[Stab.scala 177:23]
  assign last_merger_45_io_result_ready = last_q_45_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_45_clock = clock;
  assign last_q_45_reset = reset;
  assign last_q_45_io_enq_valid = last_merger_45_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_45_io_enq_bits = last_merger_45_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_45_io_deq_ready = last_merger_46_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_46_clock = clock;
  assign last_merger_46_reset = reset;
  assign last_merger_46_io_stream1_valid = last_q_45_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_46_io_stream1_bits = last_q_45_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_46_io_stream2_valid = io_stream_in_47_valid; // @[Stab.scala 177:23]
  assign last_merger_46_io_stream2_bits = io_stream_in_47_bits; // @[Stab.scala 177:23]
  assign last_merger_46_io_result_ready = last_q_46_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_46_clock = clock;
  assign last_q_46_reset = reset;
  assign last_q_46_io_enq_valid = last_merger_46_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_46_io_enq_bits = last_merger_46_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_46_io_deq_ready = last_merger_47_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_47_clock = clock;
  assign last_merger_47_reset = reset;
  assign last_merger_47_io_stream1_valid = last_q_46_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_47_io_stream1_bits = last_q_46_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_47_io_stream2_valid = io_stream_in_48_valid; // @[Stab.scala 177:23]
  assign last_merger_47_io_stream2_bits = io_stream_in_48_bits; // @[Stab.scala 177:23]
  assign last_merger_47_io_result_ready = last_q_47_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_47_clock = clock;
  assign last_q_47_reset = reset;
  assign last_q_47_io_enq_valid = last_merger_47_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_47_io_enq_bits = last_merger_47_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_47_io_deq_ready = last_merger_48_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_48_clock = clock;
  assign last_merger_48_reset = reset;
  assign last_merger_48_io_stream1_valid = last_q_47_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_48_io_stream1_bits = last_q_47_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_48_io_stream2_valid = io_stream_in_49_valid; // @[Stab.scala 177:23]
  assign last_merger_48_io_stream2_bits = io_stream_in_49_bits; // @[Stab.scala 177:23]
  assign last_merger_48_io_result_ready = last_q_48_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_48_clock = clock;
  assign last_q_48_reset = reset;
  assign last_q_48_io_enq_valid = last_merger_48_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_48_io_enq_bits = last_merger_48_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_48_io_deq_ready = last_merger_49_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_49_clock = clock;
  assign last_merger_49_reset = reset;
  assign last_merger_49_io_stream1_valid = last_q_48_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_49_io_stream1_bits = last_q_48_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_49_io_stream2_valid = io_stream_in_50_valid; // @[Stab.scala 177:23]
  assign last_merger_49_io_stream2_bits = io_stream_in_50_bits; // @[Stab.scala 177:23]
  assign last_merger_49_io_result_ready = last_q_49_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_49_clock = clock;
  assign last_q_49_reset = reset;
  assign last_q_49_io_enq_valid = last_merger_49_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_49_io_enq_bits = last_merger_49_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_49_io_deq_ready = last_merger_50_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_50_clock = clock;
  assign last_merger_50_reset = reset;
  assign last_merger_50_io_stream1_valid = last_q_49_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_50_io_stream1_bits = last_q_49_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_50_io_stream2_valid = io_stream_in_51_valid; // @[Stab.scala 177:23]
  assign last_merger_50_io_stream2_bits = io_stream_in_51_bits; // @[Stab.scala 177:23]
  assign last_merger_50_io_result_ready = last_q_50_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_50_clock = clock;
  assign last_q_50_reset = reset;
  assign last_q_50_io_enq_valid = last_merger_50_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_50_io_enq_bits = last_merger_50_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_50_io_deq_ready = last_merger_51_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_51_clock = clock;
  assign last_merger_51_reset = reset;
  assign last_merger_51_io_stream1_valid = last_q_50_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_51_io_stream1_bits = last_q_50_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_51_io_stream2_valid = io_stream_in_52_valid; // @[Stab.scala 177:23]
  assign last_merger_51_io_stream2_bits = io_stream_in_52_bits; // @[Stab.scala 177:23]
  assign last_merger_51_io_result_ready = last_q_51_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_51_clock = clock;
  assign last_q_51_reset = reset;
  assign last_q_51_io_enq_valid = last_merger_51_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_51_io_enq_bits = last_merger_51_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_51_io_deq_ready = last_merger_52_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_52_clock = clock;
  assign last_merger_52_reset = reset;
  assign last_merger_52_io_stream1_valid = last_q_51_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_52_io_stream1_bits = last_q_51_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_52_io_stream2_valid = io_stream_in_53_valid; // @[Stab.scala 177:23]
  assign last_merger_52_io_stream2_bits = io_stream_in_53_bits; // @[Stab.scala 177:23]
  assign last_merger_52_io_result_ready = last_q_52_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_52_clock = clock;
  assign last_q_52_reset = reset;
  assign last_q_52_io_enq_valid = last_merger_52_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_52_io_enq_bits = last_merger_52_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_52_io_deq_ready = last_merger_53_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_53_clock = clock;
  assign last_merger_53_reset = reset;
  assign last_merger_53_io_stream1_valid = last_q_52_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_53_io_stream1_bits = last_q_52_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_53_io_stream2_valid = io_stream_in_54_valid; // @[Stab.scala 177:23]
  assign last_merger_53_io_stream2_bits = io_stream_in_54_bits; // @[Stab.scala 177:23]
  assign last_merger_53_io_result_ready = last_q_53_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_53_clock = clock;
  assign last_q_53_reset = reset;
  assign last_q_53_io_enq_valid = last_merger_53_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_53_io_enq_bits = last_merger_53_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_53_io_deq_ready = last_merger_54_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_54_clock = clock;
  assign last_merger_54_reset = reset;
  assign last_merger_54_io_stream1_valid = last_q_53_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_54_io_stream1_bits = last_q_53_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_54_io_stream2_valid = io_stream_in_55_valid; // @[Stab.scala 177:23]
  assign last_merger_54_io_stream2_bits = io_stream_in_55_bits; // @[Stab.scala 177:23]
  assign last_merger_54_io_result_ready = last_q_54_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_54_clock = clock;
  assign last_q_54_reset = reset;
  assign last_q_54_io_enq_valid = last_merger_54_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_54_io_enq_bits = last_merger_54_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_54_io_deq_ready = last_merger_55_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_55_clock = clock;
  assign last_merger_55_reset = reset;
  assign last_merger_55_io_stream1_valid = last_q_54_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_55_io_stream1_bits = last_q_54_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_55_io_stream2_valid = io_stream_in_56_valid; // @[Stab.scala 177:23]
  assign last_merger_55_io_stream2_bits = io_stream_in_56_bits; // @[Stab.scala 177:23]
  assign last_merger_55_io_result_ready = last_q_55_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_55_clock = clock;
  assign last_q_55_reset = reset;
  assign last_q_55_io_enq_valid = last_merger_55_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_55_io_enq_bits = last_merger_55_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_55_io_deq_ready = last_merger_56_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_56_clock = clock;
  assign last_merger_56_reset = reset;
  assign last_merger_56_io_stream1_valid = last_q_55_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_56_io_stream1_bits = last_q_55_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_56_io_stream2_valid = io_stream_in_57_valid; // @[Stab.scala 177:23]
  assign last_merger_56_io_stream2_bits = io_stream_in_57_bits; // @[Stab.scala 177:23]
  assign last_merger_56_io_result_ready = last_q_56_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_56_clock = clock;
  assign last_q_56_reset = reset;
  assign last_q_56_io_enq_valid = last_merger_56_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_56_io_enq_bits = last_merger_56_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_56_io_deq_ready = last_merger_57_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_57_clock = clock;
  assign last_merger_57_reset = reset;
  assign last_merger_57_io_stream1_valid = last_q_56_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_57_io_stream1_bits = last_q_56_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_57_io_stream2_valid = io_stream_in_58_valid; // @[Stab.scala 177:23]
  assign last_merger_57_io_stream2_bits = io_stream_in_58_bits; // @[Stab.scala 177:23]
  assign last_merger_57_io_result_ready = last_q_57_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_57_clock = clock;
  assign last_q_57_reset = reset;
  assign last_q_57_io_enq_valid = last_merger_57_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_57_io_enq_bits = last_merger_57_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_57_io_deq_ready = last_merger_58_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_58_clock = clock;
  assign last_merger_58_reset = reset;
  assign last_merger_58_io_stream1_valid = last_q_57_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_58_io_stream1_bits = last_q_57_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_58_io_stream2_valid = io_stream_in_59_valid; // @[Stab.scala 177:23]
  assign last_merger_58_io_stream2_bits = io_stream_in_59_bits; // @[Stab.scala 177:23]
  assign last_merger_58_io_result_ready = last_q_58_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_58_clock = clock;
  assign last_q_58_reset = reset;
  assign last_q_58_io_enq_valid = last_merger_58_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_58_io_enq_bits = last_merger_58_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_58_io_deq_ready = last_merger_59_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_59_clock = clock;
  assign last_merger_59_reset = reset;
  assign last_merger_59_io_stream1_valid = last_q_58_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_59_io_stream1_bits = last_q_58_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_59_io_stream2_valid = io_stream_in_60_valid; // @[Stab.scala 177:23]
  assign last_merger_59_io_stream2_bits = io_stream_in_60_bits; // @[Stab.scala 177:23]
  assign last_merger_59_io_result_ready = last_q_59_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_59_clock = clock;
  assign last_q_59_reset = reset;
  assign last_q_59_io_enq_valid = last_merger_59_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_59_io_enq_bits = last_merger_59_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_59_io_deq_ready = last_merger_60_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_60_clock = clock;
  assign last_merger_60_reset = reset;
  assign last_merger_60_io_stream1_valid = last_q_59_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_60_io_stream1_bits = last_q_59_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_60_io_stream2_valid = io_stream_in_61_valid; // @[Stab.scala 177:23]
  assign last_merger_60_io_stream2_bits = io_stream_in_61_bits; // @[Stab.scala 177:23]
  assign last_merger_60_io_result_ready = last_q_60_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_60_clock = clock;
  assign last_q_60_reset = reset;
  assign last_q_60_io_enq_valid = last_merger_60_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_60_io_enq_bits = last_merger_60_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_60_io_deq_ready = last_merger_61_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_61_clock = clock;
  assign last_merger_61_reset = reset;
  assign last_merger_61_io_stream1_valid = last_q_60_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_61_io_stream1_bits = last_q_60_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_61_io_stream2_valid = io_stream_in_62_valid; // @[Stab.scala 177:23]
  assign last_merger_61_io_stream2_bits = io_stream_in_62_bits; // @[Stab.scala 177:23]
  assign last_merger_61_io_result_ready = last_q_61_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_61_clock = clock;
  assign last_q_61_reset = reset;
  assign last_q_61_io_enq_valid = last_merger_61_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_61_io_enq_bits = last_merger_61_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_61_io_deq_ready = last_merger_62_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_62_clock = clock;
  assign last_merger_62_reset = reset;
  assign last_merger_62_io_stream1_valid = last_q_61_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_62_io_stream1_bits = last_q_61_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_62_io_stream2_valid = io_stream_in_63_valid; // @[Stab.scala 177:23]
  assign last_merger_62_io_stream2_bits = io_stream_in_63_bits; // @[Stab.scala 177:23]
  assign last_merger_62_io_result_ready = last_q_62_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_62_clock = clock;
  assign last_q_62_reset = reset;
  assign last_q_62_io_enq_valid = last_merger_62_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_62_io_enq_bits = last_merger_62_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_62_io_deq_ready = last_merger_63_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_63_clock = clock;
  assign last_merger_63_reset = reset;
  assign last_merger_63_io_stream1_valid = last_q_62_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_63_io_stream1_bits = last_q_62_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_63_io_stream2_valid = io_stream_in_64_valid; // @[Stab.scala 177:23]
  assign last_merger_63_io_stream2_bits = io_stream_in_64_bits; // @[Stab.scala 177:23]
  assign last_merger_63_io_result_ready = last_q_63_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_63_clock = clock;
  assign last_q_63_reset = reset;
  assign last_q_63_io_enq_valid = last_merger_63_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_63_io_enq_bits = last_merger_63_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_63_io_deq_ready = last_merger_64_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_64_clock = clock;
  assign last_merger_64_reset = reset;
  assign last_merger_64_io_stream1_valid = last_q_63_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_64_io_stream1_bits = last_q_63_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_64_io_stream2_valid = io_stream_in_65_valid; // @[Stab.scala 177:23]
  assign last_merger_64_io_stream2_bits = io_stream_in_65_bits; // @[Stab.scala 177:23]
  assign last_merger_64_io_result_ready = last_q_64_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_64_clock = clock;
  assign last_q_64_reset = reset;
  assign last_q_64_io_enq_valid = last_merger_64_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_64_io_enq_bits = last_merger_64_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_64_io_deq_ready = last_merger_65_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_65_clock = clock;
  assign last_merger_65_reset = reset;
  assign last_merger_65_io_stream1_valid = last_q_64_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_65_io_stream1_bits = last_q_64_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_65_io_stream2_valid = io_stream_in_66_valid; // @[Stab.scala 177:23]
  assign last_merger_65_io_stream2_bits = io_stream_in_66_bits; // @[Stab.scala 177:23]
  assign last_merger_65_io_result_ready = last_q_65_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_65_clock = clock;
  assign last_q_65_reset = reset;
  assign last_q_65_io_enq_valid = last_merger_65_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_65_io_enq_bits = last_merger_65_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_65_io_deq_ready = last_merger_66_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_66_clock = clock;
  assign last_merger_66_reset = reset;
  assign last_merger_66_io_stream1_valid = last_q_65_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_66_io_stream1_bits = last_q_65_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_66_io_stream2_valid = io_stream_in_67_valid; // @[Stab.scala 177:23]
  assign last_merger_66_io_stream2_bits = io_stream_in_67_bits; // @[Stab.scala 177:23]
  assign last_merger_66_io_result_ready = last_q_66_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_66_clock = clock;
  assign last_q_66_reset = reset;
  assign last_q_66_io_enq_valid = last_merger_66_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_66_io_enq_bits = last_merger_66_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_66_io_deq_ready = last_merger_67_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_67_clock = clock;
  assign last_merger_67_reset = reset;
  assign last_merger_67_io_stream1_valid = last_q_66_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_67_io_stream1_bits = last_q_66_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_67_io_stream2_valid = io_stream_in_68_valid; // @[Stab.scala 177:23]
  assign last_merger_67_io_stream2_bits = io_stream_in_68_bits; // @[Stab.scala 177:23]
  assign last_merger_67_io_result_ready = last_q_67_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_67_clock = clock;
  assign last_q_67_reset = reset;
  assign last_q_67_io_enq_valid = last_merger_67_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_67_io_enq_bits = last_merger_67_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_67_io_deq_ready = last_merger_68_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_68_clock = clock;
  assign last_merger_68_reset = reset;
  assign last_merger_68_io_stream1_valid = last_q_67_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_68_io_stream1_bits = last_q_67_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_68_io_stream2_valid = io_stream_in_69_valid; // @[Stab.scala 177:23]
  assign last_merger_68_io_stream2_bits = io_stream_in_69_bits; // @[Stab.scala 177:23]
  assign last_merger_68_io_result_ready = last_q_68_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_68_clock = clock;
  assign last_q_68_reset = reset;
  assign last_q_68_io_enq_valid = last_merger_68_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_68_io_enq_bits = last_merger_68_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_68_io_deq_ready = last_merger_69_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_69_clock = clock;
  assign last_merger_69_reset = reset;
  assign last_merger_69_io_stream1_valid = last_q_68_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_69_io_stream1_bits = last_q_68_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_69_io_stream2_valid = io_stream_in_70_valid; // @[Stab.scala 177:23]
  assign last_merger_69_io_stream2_bits = io_stream_in_70_bits; // @[Stab.scala 177:23]
  assign last_merger_69_io_result_ready = last_q_69_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_69_clock = clock;
  assign last_q_69_reset = reset;
  assign last_q_69_io_enq_valid = last_merger_69_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_69_io_enq_bits = last_merger_69_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_69_io_deq_ready = last_merger_70_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_70_clock = clock;
  assign last_merger_70_reset = reset;
  assign last_merger_70_io_stream1_valid = last_q_69_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_70_io_stream1_bits = last_q_69_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_70_io_stream2_valid = io_stream_in_71_valid; // @[Stab.scala 177:23]
  assign last_merger_70_io_stream2_bits = io_stream_in_71_bits; // @[Stab.scala 177:23]
  assign last_merger_70_io_result_ready = last_q_70_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_70_clock = clock;
  assign last_q_70_reset = reset;
  assign last_q_70_io_enq_valid = last_merger_70_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_70_io_enq_bits = last_merger_70_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_70_io_deq_ready = last_merger_71_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_71_clock = clock;
  assign last_merger_71_reset = reset;
  assign last_merger_71_io_stream1_valid = last_q_70_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_71_io_stream1_bits = last_q_70_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_71_io_stream2_valid = io_stream_in_72_valid; // @[Stab.scala 177:23]
  assign last_merger_71_io_stream2_bits = io_stream_in_72_bits; // @[Stab.scala 177:23]
  assign last_merger_71_io_result_ready = last_q_71_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_71_clock = clock;
  assign last_q_71_reset = reset;
  assign last_q_71_io_enq_valid = last_merger_71_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_71_io_enq_bits = last_merger_71_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_71_io_deq_ready = last_merger_72_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_72_clock = clock;
  assign last_merger_72_reset = reset;
  assign last_merger_72_io_stream1_valid = last_q_71_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_72_io_stream1_bits = last_q_71_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_72_io_stream2_valid = io_stream_in_73_valid; // @[Stab.scala 177:23]
  assign last_merger_72_io_stream2_bits = io_stream_in_73_bits; // @[Stab.scala 177:23]
  assign last_merger_72_io_result_ready = last_q_72_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_72_clock = clock;
  assign last_q_72_reset = reset;
  assign last_q_72_io_enq_valid = last_merger_72_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_72_io_enq_bits = last_merger_72_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_72_io_deq_ready = last_merger_73_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_73_clock = clock;
  assign last_merger_73_reset = reset;
  assign last_merger_73_io_stream1_valid = last_q_72_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_73_io_stream1_bits = last_q_72_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_73_io_stream2_valid = io_stream_in_74_valid; // @[Stab.scala 177:23]
  assign last_merger_73_io_stream2_bits = io_stream_in_74_bits; // @[Stab.scala 177:23]
  assign last_merger_73_io_result_ready = last_q_73_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_73_clock = clock;
  assign last_q_73_reset = reset;
  assign last_q_73_io_enq_valid = last_merger_73_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_73_io_enq_bits = last_merger_73_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_73_io_deq_ready = last_merger_74_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_74_clock = clock;
  assign last_merger_74_reset = reset;
  assign last_merger_74_io_stream1_valid = last_q_73_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_74_io_stream1_bits = last_q_73_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_74_io_stream2_valid = io_stream_in_75_valid; // @[Stab.scala 177:23]
  assign last_merger_74_io_stream2_bits = io_stream_in_75_bits; // @[Stab.scala 177:23]
  assign last_merger_74_io_result_ready = last_q_74_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_74_clock = clock;
  assign last_q_74_reset = reset;
  assign last_q_74_io_enq_valid = last_merger_74_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_74_io_enq_bits = last_merger_74_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_74_io_deq_ready = last_merger_75_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_75_clock = clock;
  assign last_merger_75_reset = reset;
  assign last_merger_75_io_stream1_valid = last_q_74_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_75_io_stream1_bits = last_q_74_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_75_io_stream2_valid = io_stream_in_76_valid; // @[Stab.scala 177:23]
  assign last_merger_75_io_stream2_bits = io_stream_in_76_bits; // @[Stab.scala 177:23]
  assign last_merger_75_io_result_ready = last_q_75_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_75_clock = clock;
  assign last_q_75_reset = reset;
  assign last_q_75_io_enq_valid = last_merger_75_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_75_io_enq_bits = last_merger_75_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_75_io_deq_ready = last_merger_76_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_76_clock = clock;
  assign last_merger_76_reset = reset;
  assign last_merger_76_io_stream1_valid = last_q_75_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_76_io_stream1_bits = last_q_75_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_76_io_stream2_valid = io_stream_in_77_valid; // @[Stab.scala 177:23]
  assign last_merger_76_io_stream2_bits = io_stream_in_77_bits; // @[Stab.scala 177:23]
  assign last_merger_76_io_result_ready = last_q_76_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_76_clock = clock;
  assign last_q_76_reset = reset;
  assign last_q_76_io_enq_valid = last_merger_76_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_76_io_enq_bits = last_merger_76_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_76_io_deq_ready = last_merger_77_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_77_clock = clock;
  assign last_merger_77_reset = reset;
  assign last_merger_77_io_stream1_valid = last_q_76_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_77_io_stream1_bits = last_q_76_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_77_io_stream2_valid = io_stream_in_78_valid; // @[Stab.scala 177:23]
  assign last_merger_77_io_stream2_bits = io_stream_in_78_bits; // @[Stab.scala 177:23]
  assign last_merger_77_io_result_ready = last_q_77_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_77_clock = clock;
  assign last_q_77_reset = reset;
  assign last_q_77_io_enq_valid = last_merger_77_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_77_io_enq_bits = last_merger_77_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_77_io_deq_ready = last_merger_78_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_78_clock = clock;
  assign last_merger_78_reset = reset;
  assign last_merger_78_io_stream1_valid = last_q_77_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_78_io_stream1_bits = last_q_77_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_78_io_stream2_valid = io_stream_in_79_valid; // @[Stab.scala 177:23]
  assign last_merger_78_io_stream2_bits = io_stream_in_79_bits; // @[Stab.scala 177:23]
  assign last_merger_78_io_result_ready = last_q_78_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_78_clock = clock;
  assign last_q_78_reset = reset;
  assign last_q_78_io_enq_valid = last_merger_78_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_78_io_enq_bits = last_merger_78_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_78_io_deq_ready = last_merger_79_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_79_clock = clock;
  assign last_merger_79_reset = reset;
  assign last_merger_79_io_stream1_valid = last_q_78_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_79_io_stream1_bits = last_q_78_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_79_io_stream2_valid = io_stream_in_80_valid; // @[Stab.scala 177:23]
  assign last_merger_79_io_stream2_bits = io_stream_in_80_bits; // @[Stab.scala 177:23]
  assign last_merger_79_io_result_ready = last_q_79_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_79_clock = clock;
  assign last_q_79_reset = reset;
  assign last_q_79_io_enq_valid = last_merger_79_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_79_io_enq_bits = last_merger_79_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_79_io_deq_ready = last_merger_80_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_80_clock = clock;
  assign last_merger_80_reset = reset;
  assign last_merger_80_io_stream1_valid = last_q_79_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_80_io_stream1_bits = last_q_79_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_80_io_stream2_valid = io_stream_in_81_valid; // @[Stab.scala 177:23]
  assign last_merger_80_io_stream2_bits = io_stream_in_81_bits; // @[Stab.scala 177:23]
  assign last_merger_80_io_result_ready = last_q_80_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_80_clock = clock;
  assign last_q_80_reset = reset;
  assign last_q_80_io_enq_valid = last_merger_80_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_80_io_enq_bits = last_merger_80_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_80_io_deq_ready = last_merger_81_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_81_clock = clock;
  assign last_merger_81_reset = reset;
  assign last_merger_81_io_stream1_valid = last_q_80_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_81_io_stream1_bits = last_q_80_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_81_io_stream2_valid = io_stream_in_82_valid; // @[Stab.scala 177:23]
  assign last_merger_81_io_stream2_bits = io_stream_in_82_bits; // @[Stab.scala 177:23]
  assign last_merger_81_io_result_ready = last_q_81_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_81_clock = clock;
  assign last_q_81_reset = reset;
  assign last_q_81_io_enq_valid = last_merger_81_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_81_io_enq_bits = last_merger_81_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_81_io_deq_ready = last_merger_82_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_82_clock = clock;
  assign last_merger_82_reset = reset;
  assign last_merger_82_io_stream1_valid = last_q_81_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_82_io_stream1_bits = last_q_81_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_82_io_stream2_valid = io_stream_in_83_valid; // @[Stab.scala 177:23]
  assign last_merger_82_io_stream2_bits = io_stream_in_83_bits; // @[Stab.scala 177:23]
  assign last_merger_82_io_result_ready = last_q_82_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_82_clock = clock;
  assign last_q_82_reset = reset;
  assign last_q_82_io_enq_valid = last_merger_82_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_82_io_enq_bits = last_merger_82_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_82_io_deq_ready = last_merger_83_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_83_clock = clock;
  assign last_merger_83_reset = reset;
  assign last_merger_83_io_stream1_valid = last_q_82_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_83_io_stream1_bits = last_q_82_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_83_io_stream2_valid = io_stream_in_84_valid; // @[Stab.scala 177:23]
  assign last_merger_83_io_stream2_bits = io_stream_in_84_bits; // @[Stab.scala 177:23]
  assign last_merger_83_io_result_ready = last_q_83_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_83_clock = clock;
  assign last_q_83_reset = reset;
  assign last_q_83_io_enq_valid = last_merger_83_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_83_io_enq_bits = last_merger_83_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_83_io_deq_ready = last_merger_84_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_84_clock = clock;
  assign last_merger_84_reset = reset;
  assign last_merger_84_io_stream1_valid = last_q_83_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_84_io_stream1_bits = last_q_83_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_84_io_stream2_valid = io_stream_in_85_valid; // @[Stab.scala 177:23]
  assign last_merger_84_io_stream2_bits = io_stream_in_85_bits; // @[Stab.scala 177:23]
  assign last_merger_84_io_result_ready = last_q_84_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_84_clock = clock;
  assign last_q_84_reset = reset;
  assign last_q_84_io_enq_valid = last_merger_84_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_84_io_enq_bits = last_merger_84_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_84_io_deq_ready = last_merger_85_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_85_clock = clock;
  assign last_merger_85_reset = reset;
  assign last_merger_85_io_stream1_valid = last_q_84_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_85_io_stream1_bits = last_q_84_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_85_io_stream2_valid = io_stream_in_86_valid; // @[Stab.scala 177:23]
  assign last_merger_85_io_stream2_bits = io_stream_in_86_bits; // @[Stab.scala 177:23]
  assign last_merger_85_io_result_ready = last_q_85_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_85_clock = clock;
  assign last_q_85_reset = reset;
  assign last_q_85_io_enq_valid = last_merger_85_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_85_io_enq_bits = last_merger_85_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_85_io_deq_ready = last_merger_86_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_86_clock = clock;
  assign last_merger_86_reset = reset;
  assign last_merger_86_io_stream1_valid = last_q_85_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_86_io_stream1_bits = last_q_85_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_86_io_stream2_valid = io_stream_in_87_valid; // @[Stab.scala 177:23]
  assign last_merger_86_io_stream2_bits = io_stream_in_87_bits; // @[Stab.scala 177:23]
  assign last_merger_86_io_result_ready = last_q_86_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_86_clock = clock;
  assign last_q_86_reset = reset;
  assign last_q_86_io_enq_valid = last_merger_86_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_86_io_enq_bits = last_merger_86_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_86_io_deq_ready = last_merger_87_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_87_clock = clock;
  assign last_merger_87_reset = reset;
  assign last_merger_87_io_stream1_valid = last_q_86_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_87_io_stream1_bits = last_q_86_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_87_io_stream2_valid = io_stream_in_88_valid; // @[Stab.scala 177:23]
  assign last_merger_87_io_stream2_bits = io_stream_in_88_bits; // @[Stab.scala 177:23]
  assign last_merger_87_io_result_ready = last_q_87_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_87_clock = clock;
  assign last_q_87_reset = reset;
  assign last_q_87_io_enq_valid = last_merger_87_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_87_io_enq_bits = last_merger_87_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_87_io_deq_ready = last_merger_88_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_88_clock = clock;
  assign last_merger_88_reset = reset;
  assign last_merger_88_io_stream1_valid = last_q_87_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_88_io_stream1_bits = last_q_87_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_88_io_stream2_valid = io_stream_in_89_valid; // @[Stab.scala 177:23]
  assign last_merger_88_io_stream2_bits = io_stream_in_89_bits; // @[Stab.scala 177:23]
  assign last_merger_88_io_result_ready = last_q_88_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_88_clock = clock;
  assign last_q_88_reset = reset;
  assign last_q_88_io_enq_valid = last_merger_88_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_88_io_enq_bits = last_merger_88_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_88_io_deq_ready = last_merger_89_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_89_clock = clock;
  assign last_merger_89_reset = reset;
  assign last_merger_89_io_stream1_valid = last_q_88_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_89_io_stream1_bits = last_q_88_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_89_io_stream2_valid = io_stream_in_90_valid; // @[Stab.scala 177:23]
  assign last_merger_89_io_stream2_bits = io_stream_in_90_bits; // @[Stab.scala 177:23]
  assign last_merger_89_io_result_ready = last_q_89_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_89_clock = clock;
  assign last_q_89_reset = reset;
  assign last_q_89_io_enq_valid = last_merger_89_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_89_io_enq_bits = last_merger_89_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_89_io_deq_ready = last_merger_90_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_90_clock = clock;
  assign last_merger_90_reset = reset;
  assign last_merger_90_io_stream1_valid = last_q_89_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_90_io_stream1_bits = last_q_89_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_90_io_stream2_valid = io_stream_in_91_valid; // @[Stab.scala 177:23]
  assign last_merger_90_io_stream2_bits = io_stream_in_91_bits; // @[Stab.scala 177:23]
  assign last_merger_90_io_result_ready = last_q_90_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_90_clock = clock;
  assign last_q_90_reset = reset;
  assign last_q_90_io_enq_valid = last_merger_90_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_90_io_enq_bits = last_merger_90_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_90_io_deq_ready = last_merger_91_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_91_clock = clock;
  assign last_merger_91_reset = reset;
  assign last_merger_91_io_stream1_valid = last_q_90_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_91_io_stream1_bits = last_q_90_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_91_io_stream2_valid = io_stream_in_92_valid; // @[Stab.scala 177:23]
  assign last_merger_91_io_stream2_bits = io_stream_in_92_bits; // @[Stab.scala 177:23]
  assign last_merger_91_io_result_ready = last_q_91_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_91_clock = clock;
  assign last_q_91_reset = reset;
  assign last_q_91_io_enq_valid = last_merger_91_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_91_io_enq_bits = last_merger_91_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_91_io_deq_ready = last_merger_92_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_92_clock = clock;
  assign last_merger_92_reset = reset;
  assign last_merger_92_io_stream1_valid = last_q_91_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_92_io_stream1_bits = last_q_91_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_92_io_stream2_valid = io_stream_in_93_valid; // @[Stab.scala 177:23]
  assign last_merger_92_io_stream2_bits = io_stream_in_93_bits; // @[Stab.scala 177:23]
  assign last_merger_92_io_result_ready = last_q_92_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_92_clock = clock;
  assign last_q_92_reset = reset;
  assign last_q_92_io_enq_valid = last_merger_92_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_92_io_enq_bits = last_merger_92_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_92_io_deq_ready = last_merger_93_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_93_clock = clock;
  assign last_merger_93_reset = reset;
  assign last_merger_93_io_stream1_valid = last_q_92_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_93_io_stream1_bits = last_q_92_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_93_io_stream2_valid = io_stream_in_94_valid; // @[Stab.scala 177:23]
  assign last_merger_93_io_stream2_bits = io_stream_in_94_bits; // @[Stab.scala 177:23]
  assign last_merger_93_io_result_ready = last_q_93_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_93_clock = clock;
  assign last_q_93_reset = reset;
  assign last_q_93_io_enq_valid = last_merger_93_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_93_io_enq_bits = last_merger_93_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_93_io_deq_ready = last_merger_94_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_94_clock = clock;
  assign last_merger_94_reset = reset;
  assign last_merger_94_io_stream1_valid = last_q_93_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_94_io_stream1_bits = last_q_93_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_94_io_stream2_valid = io_stream_in_95_valid; // @[Stab.scala 177:23]
  assign last_merger_94_io_stream2_bits = io_stream_in_95_bits; // @[Stab.scala 177:23]
  assign last_merger_94_io_result_ready = last_q_94_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_94_clock = clock;
  assign last_q_94_reset = reset;
  assign last_q_94_io_enq_valid = last_merger_94_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_94_io_enq_bits = last_merger_94_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_94_io_deq_ready = last_merger_95_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_95_clock = clock;
  assign last_merger_95_reset = reset;
  assign last_merger_95_io_stream1_valid = last_q_94_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_95_io_stream1_bits = last_q_94_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_95_io_stream2_valid = io_stream_in_96_valid; // @[Stab.scala 177:23]
  assign last_merger_95_io_stream2_bits = io_stream_in_96_bits; // @[Stab.scala 177:23]
  assign last_merger_95_io_result_ready = last_q_95_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_95_clock = clock;
  assign last_q_95_reset = reset;
  assign last_q_95_io_enq_valid = last_merger_95_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_95_io_enq_bits = last_merger_95_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_95_io_deq_ready = last_merger_96_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_96_clock = clock;
  assign last_merger_96_reset = reset;
  assign last_merger_96_io_stream1_valid = last_q_95_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_96_io_stream1_bits = last_q_95_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_96_io_stream2_valid = io_stream_in_97_valid; // @[Stab.scala 177:23]
  assign last_merger_96_io_stream2_bits = io_stream_in_97_bits; // @[Stab.scala 177:23]
  assign last_merger_96_io_result_ready = last_q_96_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_96_clock = clock;
  assign last_q_96_reset = reset;
  assign last_q_96_io_enq_valid = last_merger_96_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_96_io_enq_bits = last_merger_96_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_96_io_deq_ready = last_merger_97_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_97_clock = clock;
  assign last_merger_97_reset = reset;
  assign last_merger_97_io_stream1_valid = last_q_96_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_97_io_stream1_bits = last_q_96_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_97_io_stream2_valid = io_stream_in_98_valid; // @[Stab.scala 177:23]
  assign last_merger_97_io_stream2_bits = io_stream_in_98_bits; // @[Stab.scala 177:23]
  assign last_merger_97_io_result_ready = last_q_97_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_97_clock = clock;
  assign last_q_97_reset = reset;
  assign last_q_97_io_enq_valid = last_merger_97_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_97_io_enq_bits = last_merger_97_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_97_io_deq_ready = last_merger_98_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_98_clock = clock;
  assign last_merger_98_reset = reset;
  assign last_merger_98_io_stream1_valid = last_q_97_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_98_io_stream1_bits = last_q_97_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_98_io_stream2_valid = io_stream_in_99_valid; // @[Stab.scala 177:23]
  assign last_merger_98_io_stream2_bits = io_stream_in_99_bits; // @[Stab.scala 177:23]
  assign last_merger_98_io_result_ready = last_q_98_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_98_clock = clock;
  assign last_q_98_reset = reset;
  assign last_q_98_io_enq_valid = last_merger_98_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_98_io_enq_bits = last_merger_98_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_98_io_deq_ready = last_merger_99_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_99_clock = clock;
  assign last_merger_99_reset = reset;
  assign last_merger_99_io_stream1_valid = last_q_98_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_99_io_stream1_bits = last_q_98_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_99_io_stream2_valid = io_stream_in_100_valid; // @[Stab.scala 177:23]
  assign last_merger_99_io_stream2_bits = io_stream_in_100_bits; // @[Stab.scala 177:23]
  assign last_merger_99_io_result_ready = last_q_99_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_99_clock = clock;
  assign last_q_99_reset = reset;
  assign last_q_99_io_enq_valid = last_merger_99_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_99_io_enq_bits = last_merger_99_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_99_io_deq_ready = last_merger_100_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_100_clock = clock;
  assign last_merger_100_reset = reset;
  assign last_merger_100_io_stream1_valid = last_q_99_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_100_io_stream1_bits = last_q_99_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_100_io_stream2_valid = io_stream_in_101_valid; // @[Stab.scala 177:23]
  assign last_merger_100_io_stream2_bits = io_stream_in_101_bits; // @[Stab.scala 177:23]
  assign last_merger_100_io_result_ready = last_q_100_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_100_clock = clock;
  assign last_q_100_reset = reset;
  assign last_q_100_io_enq_valid = last_merger_100_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_100_io_enq_bits = last_merger_100_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_100_io_deq_ready = last_merger_101_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_101_clock = clock;
  assign last_merger_101_reset = reset;
  assign last_merger_101_io_stream1_valid = last_q_100_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_101_io_stream1_bits = last_q_100_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_101_io_stream2_valid = io_stream_in_102_valid; // @[Stab.scala 177:23]
  assign last_merger_101_io_stream2_bits = io_stream_in_102_bits; // @[Stab.scala 177:23]
  assign last_merger_101_io_result_ready = last_q_101_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_101_clock = clock;
  assign last_q_101_reset = reset;
  assign last_q_101_io_enq_valid = last_merger_101_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_101_io_enq_bits = last_merger_101_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_101_io_deq_ready = last_merger_102_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_102_clock = clock;
  assign last_merger_102_reset = reset;
  assign last_merger_102_io_stream1_valid = last_q_101_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_102_io_stream1_bits = last_q_101_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_102_io_stream2_valid = io_stream_in_103_valid; // @[Stab.scala 177:23]
  assign last_merger_102_io_stream2_bits = io_stream_in_103_bits; // @[Stab.scala 177:23]
  assign last_merger_102_io_result_ready = last_q_102_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_102_clock = clock;
  assign last_q_102_reset = reset;
  assign last_q_102_io_enq_valid = last_merger_102_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_102_io_enq_bits = last_merger_102_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_102_io_deq_ready = last_merger_103_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_103_clock = clock;
  assign last_merger_103_reset = reset;
  assign last_merger_103_io_stream1_valid = last_q_102_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_103_io_stream1_bits = last_q_102_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_103_io_stream2_valid = io_stream_in_104_valid; // @[Stab.scala 177:23]
  assign last_merger_103_io_stream2_bits = io_stream_in_104_bits; // @[Stab.scala 177:23]
  assign last_merger_103_io_result_ready = last_q_103_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_103_clock = clock;
  assign last_q_103_reset = reset;
  assign last_q_103_io_enq_valid = last_merger_103_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_103_io_enq_bits = last_merger_103_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_103_io_deq_ready = last_merger_104_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_104_clock = clock;
  assign last_merger_104_reset = reset;
  assign last_merger_104_io_stream1_valid = last_q_103_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_104_io_stream1_bits = last_q_103_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_104_io_stream2_valid = io_stream_in_105_valid; // @[Stab.scala 177:23]
  assign last_merger_104_io_stream2_bits = io_stream_in_105_bits; // @[Stab.scala 177:23]
  assign last_merger_104_io_result_ready = last_q_104_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_104_clock = clock;
  assign last_q_104_reset = reset;
  assign last_q_104_io_enq_valid = last_merger_104_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_104_io_enq_bits = last_merger_104_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_104_io_deq_ready = last_merger_105_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_105_clock = clock;
  assign last_merger_105_reset = reset;
  assign last_merger_105_io_stream1_valid = last_q_104_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_105_io_stream1_bits = last_q_104_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_105_io_stream2_valid = io_stream_in_106_valid; // @[Stab.scala 177:23]
  assign last_merger_105_io_stream2_bits = io_stream_in_106_bits; // @[Stab.scala 177:23]
  assign last_merger_105_io_result_ready = last_q_105_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_105_clock = clock;
  assign last_q_105_reset = reset;
  assign last_q_105_io_enq_valid = last_merger_105_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_105_io_enq_bits = last_merger_105_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_105_io_deq_ready = last_merger_106_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_106_clock = clock;
  assign last_merger_106_reset = reset;
  assign last_merger_106_io_stream1_valid = last_q_105_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_106_io_stream1_bits = last_q_105_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_106_io_stream2_valid = io_stream_in_107_valid; // @[Stab.scala 177:23]
  assign last_merger_106_io_stream2_bits = io_stream_in_107_bits; // @[Stab.scala 177:23]
  assign last_merger_106_io_result_ready = last_q_106_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_106_clock = clock;
  assign last_q_106_reset = reset;
  assign last_q_106_io_enq_valid = last_merger_106_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_106_io_enq_bits = last_merger_106_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_106_io_deq_ready = last_merger_107_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_107_clock = clock;
  assign last_merger_107_reset = reset;
  assign last_merger_107_io_stream1_valid = last_q_106_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_107_io_stream1_bits = last_q_106_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_107_io_stream2_valid = io_stream_in_108_valid; // @[Stab.scala 177:23]
  assign last_merger_107_io_stream2_bits = io_stream_in_108_bits; // @[Stab.scala 177:23]
  assign last_merger_107_io_result_ready = last_q_107_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_107_clock = clock;
  assign last_q_107_reset = reset;
  assign last_q_107_io_enq_valid = last_merger_107_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_107_io_enq_bits = last_merger_107_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_107_io_deq_ready = last_merger_108_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_108_clock = clock;
  assign last_merger_108_reset = reset;
  assign last_merger_108_io_stream1_valid = last_q_107_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_108_io_stream1_bits = last_q_107_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_108_io_stream2_valid = io_stream_in_109_valid; // @[Stab.scala 177:23]
  assign last_merger_108_io_stream2_bits = io_stream_in_109_bits; // @[Stab.scala 177:23]
  assign last_merger_108_io_result_ready = last_q_108_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_108_clock = clock;
  assign last_q_108_reset = reset;
  assign last_q_108_io_enq_valid = last_merger_108_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_108_io_enq_bits = last_merger_108_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_108_io_deq_ready = last_merger_109_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_109_clock = clock;
  assign last_merger_109_reset = reset;
  assign last_merger_109_io_stream1_valid = last_q_108_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_109_io_stream1_bits = last_q_108_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_109_io_stream2_valid = io_stream_in_110_valid; // @[Stab.scala 177:23]
  assign last_merger_109_io_stream2_bits = io_stream_in_110_bits; // @[Stab.scala 177:23]
  assign last_merger_109_io_result_ready = last_q_109_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_109_clock = clock;
  assign last_q_109_reset = reset;
  assign last_q_109_io_enq_valid = last_merger_109_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_109_io_enq_bits = last_merger_109_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_109_io_deq_ready = last_merger_110_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_110_clock = clock;
  assign last_merger_110_reset = reset;
  assign last_merger_110_io_stream1_valid = last_q_109_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_110_io_stream1_bits = last_q_109_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_110_io_stream2_valid = io_stream_in_111_valid; // @[Stab.scala 177:23]
  assign last_merger_110_io_stream2_bits = io_stream_in_111_bits; // @[Stab.scala 177:23]
  assign last_merger_110_io_result_ready = last_q_110_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_110_clock = clock;
  assign last_q_110_reset = reset;
  assign last_q_110_io_enq_valid = last_merger_110_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_110_io_enq_bits = last_merger_110_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_110_io_deq_ready = last_merger_111_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_111_clock = clock;
  assign last_merger_111_reset = reset;
  assign last_merger_111_io_stream1_valid = last_q_110_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_111_io_stream1_bits = last_q_110_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_111_io_stream2_valid = io_stream_in_112_valid; // @[Stab.scala 177:23]
  assign last_merger_111_io_stream2_bits = io_stream_in_112_bits; // @[Stab.scala 177:23]
  assign last_merger_111_io_result_ready = last_q_111_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_111_clock = clock;
  assign last_q_111_reset = reset;
  assign last_q_111_io_enq_valid = last_merger_111_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_111_io_enq_bits = last_merger_111_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_111_io_deq_ready = last_merger_112_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_112_clock = clock;
  assign last_merger_112_reset = reset;
  assign last_merger_112_io_stream1_valid = last_q_111_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_112_io_stream1_bits = last_q_111_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_112_io_stream2_valid = io_stream_in_113_valid; // @[Stab.scala 177:23]
  assign last_merger_112_io_stream2_bits = io_stream_in_113_bits; // @[Stab.scala 177:23]
  assign last_merger_112_io_result_ready = last_q_112_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_112_clock = clock;
  assign last_q_112_reset = reset;
  assign last_q_112_io_enq_valid = last_merger_112_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_112_io_enq_bits = last_merger_112_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_112_io_deq_ready = last_merger_113_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_113_clock = clock;
  assign last_merger_113_reset = reset;
  assign last_merger_113_io_stream1_valid = last_q_112_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_113_io_stream1_bits = last_q_112_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_113_io_stream2_valid = io_stream_in_114_valid; // @[Stab.scala 177:23]
  assign last_merger_113_io_stream2_bits = io_stream_in_114_bits; // @[Stab.scala 177:23]
  assign last_merger_113_io_result_ready = last_q_113_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_113_clock = clock;
  assign last_q_113_reset = reset;
  assign last_q_113_io_enq_valid = last_merger_113_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_113_io_enq_bits = last_merger_113_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_113_io_deq_ready = last_merger_114_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_114_clock = clock;
  assign last_merger_114_reset = reset;
  assign last_merger_114_io_stream1_valid = last_q_113_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_114_io_stream1_bits = last_q_113_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_114_io_stream2_valid = io_stream_in_115_valid; // @[Stab.scala 177:23]
  assign last_merger_114_io_stream2_bits = io_stream_in_115_bits; // @[Stab.scala 177:23]
  assign last_merger_114_io_result_ready = last_q_114_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_114_clock = clock;
  assign last_q_114_reset = reset;
  assign last_q_114_io_enq_valid = last_merger_114_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_114_io_enq_bits = last_merger_114_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_114_io_deq_ready = last_merger_115_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_115_clock = clock;
  assign last_merger_115_reset = reset;
  assign last_merger_115_io_stream1_valid = last_q_114_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_115_io_stream1_bits = last_q_114_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_115_io_stream2_valid = io_stream_in_116_valid; // @[Stab.scala 177:23]
  assign last_merger_115_io_stream2_bits = io_stream_in_116_bits; // @[Stab.scala 177:23]
  assign last_merger_115_io_result_ready = last_q_115_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_115_clock = clock;
  assign last_q_115_reset = reset;
  assign last_q_115_io_enq_valid = last_merger_115_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_115_io_enq_bits = last_merger_115_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_115_io_deq_ready = last_merger_116_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_116_clock = clock;
  assign last_merger_116_reset = reset;
  assign last_merger_116_io_stream1_valid = last_q_115_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_116_io_stream1_bits = last_q_115_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_116_io_stream2_valid = io_stream_in_117_valid; // @[Stab.scala 177:23]
  assign last_merger_116_io_stream2_bits = io_stream_in_117_bits; // @[Stab.scala 177:23]
  assign last_merger_116_io_result_ready = last_q_116_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_116_clock = clock;
  assign last_q_116_reset = reset;
  assign last_q_116_io_enq_valid = last_merger_116_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_116_io_enq_bits = last_merger_116_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_116_io_deq_ready = last_merger_117_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_117_clock = clock;
  assign last_merger_117_reset = reset;
  assign last_merger_117_io_stream1_valid = last_q_116_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_117_io_stream1_bits = last_q_116_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_117_io_stream2_valid = io_stream_in_118_valid; // @[Stab.scala 177:23]
  assign last_merger_117_io_stream2_bits = io_stream_in_118_bits; // @[Stab.scala 177:23]
  assign last_merger_117_io_result_ready = last_q_117_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_117_clock = clock;
  assign last_q_117_reset = reset;
  assign last_q_117_io_enq_valid = last_merger_117_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_117_io_enq_bits = last_merger_117_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_117_io_deq_ready = last_merger_118_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_118_clock = clock;
  assign last_merger_118_reset = reset;
  assign last_merger_118_io_stream1_valid = last_q_117_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_118_io_stream1_bits = last_q_117_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_118_io_stream2_valid = io_stream_in_119_valid; // @[Stab.scala 177:23]
  assign last_merger_118_io_stream2_bits = io_stream_in_119_bits; // @[Stab.scala 177:23]
  assign last_merger_118_io_result_ready = last_q_118_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_118_clock = clock;
  assign last_q_118_reset = reset;
  assign last_q_118_io_enq_valid = last_merger_118_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_118_io_enq_bits = last_merger_118_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_118_io_deq_ready = last_merger_119_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_119_clock = clock;
  assign last_merger_119_reset = reset;
  assign last_merger_119_io_stream1_valid = last_q_118_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_119_io_stream1_bits = last_q_118_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_119_io_stream2_valid = io_stream_in_120_valid; // @[Stab.scala 177:23]
  assign last_merger_119_io_stream2_bits = io_stream_in_120_bits; // @[Stab.scala 177:23]
  assign last_merger_119_io_result_ready = last_q_119_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_119_clock = clock;
  assign last_q_119_reset = reset;
  assign last_q_119_io_enq_valid = last_merger_119_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_119_io_enq_bits = last_merger_119_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_119_io_deq_ready = last_merger_120_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_120_clock = clock;
  assign last_merger_120_reset = reset;
  assign last_merger_120_io_stream1_valid = last_q_119_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_120_io_stream1_bits = last_q_119_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_120_io_stream2_valid = io_stream_in_121_valid; // @[Stab.scala 177:23]
  assign last_merger_120_io_stream2_bits = io_stream_in_121_bits; // @[Stab.scala 177:23]
  assign last_merger_120_io_result_ready = last_q_120_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_120_clock = clock;
  assign last_q_120_reset = reset;
  assign last_q_120_io_enq_valid = last_merger_120_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_120_io_enq_bits = last_merger_120_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_120_io_deq_ready = last_merger_121_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_121_clock = clock;
  assign last_merger_121_reset = reset;
  assign last_merger_121_io_stream1_valid = last_q_120_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_121_io_stream1_bits = last_q_120_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_121_io_stream2_valid = io_stream_in_122_valid; // @[Stab.scala 177:23]
  assign last_merger_121_io_stream2_bits = io_stream_in_122_bits; // @[Stab.scala 177:23]
  assign last_merger_121_io_result_ready = last_q_121_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_121_clock = clock;
  assign last_q_121_reset = reset;
  assign last_q_121_io_enq_valid = last_merger_121_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_121_io_enq_bits = last_merger_121_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_121_io_deq_ready = last_merger_122_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_122_clock = clock;
  assign last_merger_122_reset = reset;
  assign last_merger_122_io_stream1_valid = last_q_121_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_122_io_stream1_bits = last_q_121_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_122_io_stream2_valid = io_stream_in_123_valid; // @[Stab.scala 177:23]
  assign last_merger_122_io_stream2_bits = io_stream_in_123_bits; // @[Stab.scala 177:23]
  assign last_merger_122_io_result_ready = last_q_122_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_122_clock = clock;
  assign last_q_122_reset = reset;
  assign last_q_122_io_enq_valid = last_merger_122_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_122_io_enq_bits = last_merger_122_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_122_io_deq_ready = last_merger_123_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_123_clock = clock;
  assign last_merger_123_reset = reset;
  assign last_merger_123_io_stream1_valid = last_q_122_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_123_io_stream1_bits = last_q_122_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_123_io_stream2_valid = io_stream_in_124_valid; // @[Stab.scala 177:23]
  assign last_merger_123_io_stream2_bits = io_stream_in_124_bits; // @[Stab.scala 177:23]
  assign last_merger_123_io_result_ready = last_q_123_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_123_clock = clock;
  assign last_q_123_reset = reset;
  assign last_q_123_io_enq_valid = last_merger_123_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_123_io_enq_bits = last_merger_123_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_123_io_deq_ready = last_merger_124_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_124_clock = clock;
  assign last_merger_124_reset = reset;
  assign last_merger_124_io_stream1_valid = last_q_123_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_124_io_stream1_bits = last_q_123_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_124_io_stream2_valid = io_stream_in_125_valid; // @[Stab.scala 177:23]
  assign last_merger_124_io_stream2_bits = io_stream_in_125_bits; // @[Stab.scala 177:23]
  assign last_merger_124_io_result_ready = last_q_124_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_124_clock = clock;
  assign last_q_124_reset = reset;
  assign last_q_124_io_enq_valid = last_merger_124_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_124_io_enq_bits = last_merger_124_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_124_io_deq_ready = last_merger_125_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_125_clock = clock;
  assign last_merger_125_reset = reset;
  assign last_merger_125_io_stream1_valid = last_q_124_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_125_io_stream1_bits = last_q_124_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_125_io_stream2_valid = io_stream_in_126_valid; // @[Stab.scala 177:23]
  assign last_merger_125_io_stream2_bits = io_stream_in_126_bits; // @[Stab.scala 177:23]
  assign last_merger_125_io_result_ready = last_q_125_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_125_clock = clock;
  assign last_q_125_reset = reset;
  assign last_q_125_io_enq_valid = last_merger_125_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_125_io_enq_bits = last_merger_125_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_125_io_deq_ready = last_merger_126_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_126_clock = clock;
  assign last_merger_126_reset = reset;
  assign last_merger_126_io_stream1_valid = last_q_125_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_126_io_stream1_bits = last_q_125_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_126_io_stream2_valid = io_stream_in_127_valid; // @[Stab.scala 177:23]
  assign last_merger_126_io_stream2_bits = io_stream_in_127_bits; // @[Stab.scala 177:23]
  assign last_merger_126_io_result_ready = last_q_126_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_126_clock = clock;
  assign last_q_126_reset = reset;
  assign last_q_126_io_enq_valid = last_merger_126_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_126_io_enq_bits = last_merger_126_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_126_io_deq_ready = last_merger_127_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_127_clock = clock;
  assign last_merger_127_reset = reset;
  assign last_merger_127_io_stream1_valid = last_q_126_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_127_io_stream1_bits = last_q_126_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_127_io_stream2_valid = io_stream_in_128_valid; // @[Stab.scala 177:23]
  assign last_merger_127_io_stream2_bits = io_stream_in_128_bits; // @[Stab.scala 177:23]
  assign last_merger_127_io_result_ready = last_q_127_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_127_clock = clock;
  assign last_q_127_reset = reset;
  assign last_q_127_io_enq_valid = last_merger_127_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_127_io_enq_bits = last_merger_127_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_127_io_deq_ready = last_merger_128_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_128_clock = clock;
  assign last_merger_128_reset = reset;
  assign last_merger_128_io_stream1_valid = last_q_127_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_128_io_stream1_bits = last_q_127_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_128_io_stream2_valid = io_stream_in_129_valid; // @[Stab.scala 177:23]
  assign last_merger_128_io_stream2_bits = io_stream_in_129_bits; // @[Stab.scala 177:23]
  assign last_merger_128_io_result_ready = last_q_128_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_128_clock = clock;
  assign last_q_128_reset = reset;
  assign last_q_128_io_enq_valid = last_merger_128_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_128_io_enq_bits = last_merger_128_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_128_io_deq_ready = last_merger_129_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_129_clock = clock;
  assign last_merger_129_reset = reset;
  assign last_merger_129_io_stream1_valid = last_q_128_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_129_io_stream1_bits = last_q_128_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_129_io_stream2_valid = io_stream_in_130_valid; // @[Stab.scala 177:23]
  assign last_merger_129_io_stream2_bits = io_stream_in_130_bits; // @[Stab.scala 177:23]
  assign last_merger_129_io_result_ready = last_q_129_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_129_clock = clock;
  assign last_q_129_reset = reset;
  assign last_q_129_io_enq_valid = last_merger_129_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_129_io_enq_bits = last_merger_129_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_129_io_deq_ready = last_merger_130_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_130_clock = clock;
  assign last_merger_130_reset = reset;
  assign last_merger_130_io_stream1_valid = last_q_129_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_130_io_stream1_bits = last_q_129_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_130_io_stream2_valid = io_stream_in_131_valid; // @[Stab.scala 177:23]
  assign last_merger_130_io_stream2_bits = io_stream_in_131_bits; // @[Stab.scala 177:23]
  assign last_merger_130_io_result_ready = last_q_130_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_130_clock = clock;
  assign last_q_130_reset = reset;
  assign last_q_130_io_enq_valid = last_merger_130_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_130_io_enq_bits = last_merger_130_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_130_io_deq_ready = last_merger_131_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_131_clock = clock;
  assign last_merger_131_reset = reset;
  assign last_merger_131_io_stream1_valid = last_q_130_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_131_io_stream1_bits = last_q_130_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_131_io_stream2_valid = io_stream_in_132_valid; // @[Stab.scala 177:23]
  assign last_merger_131_io_stream2_bits = io_stream_in_132_bits; // @[Stab.scala 177:23]
  assign last_merger_131_io_result_ready = last_q_131_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_131_clock = clock;
  assign last_q_131_reset = reset;
  assign last_q_131_io_enq_valid = last_merger_131_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_131_io_enq_bits = last_merger_131_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_131_io_deq_ready = last_merger_132_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_132_clock = clock;
  assign last_merger_132_reset = reset;
  assign last_merger_132_io_stream1_valid = last_q_131_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_132_io_stream1_bits = last_q_131_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_132_io_stream2_valid = io_stream_in_133_valid; // @[Stab.scala 177:23]
  assign last_merger_132_io_stream2_bits = io_stream_in_133_bits; // @[Stab.scala 177:23]
  assign last_merger_132_io_result_ready = last_q_132_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_132_clock = clock;
  assign last_q_132_reset = reset;
  assign last_q_132_io_enq_valid = last_merger_132_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_132_io_enq_bits = last_merger_132_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_132_io_deq_ready = last_merger_133_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_133_clock = clock;
  assign last_merger_133_reset = reset;
  assign last_merger_133_io_stream1_valid = last_q_132_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_133_io_stream1_bits = last_q_132_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_133_io_stream2_valid = io_stream_in_134_valid; // @[Stab.scala 177:23]
  assign last_merger_133_io_stream2_bits = io_stream_in_134_bits; // @[Stab.scala 177:23]
  assign last_merger_133_io_result_ready = last_q_133_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_133_clock = clock;
  assign last_q_133_reset = reset;
  assign last_q_133_io_enq_valid = last_merger_133_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_133_io_enq_bits = last_merger_133_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_133_io_deq_ready = last_merger_134_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_134_clock = clock;
  assign last_merger_134_reset = reset;
  assign last_merger_134_io_stream1_valid = last_q_133_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_134_io_stream1_bits = last_q_133_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_134_io_stream2_valid = io_stream_in_135_valid; // @[Stab.scala 177:23]
  assign last_merger_134_io_stream2_bits = io_stream_in_135_bits; // @[Stab.scala 177:23]
  assign last_merger_134_io_result_ready = last_q_134_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_134_clock = clock;
  assign last_q_134_reset = reset;
  assign last_q_134_io_enq_valid = last_merger_134_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_134_io_enq_bits = last_merger_134_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_134_io_deq_ready = last_merger_135_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_135_clock = clock;
  assign last_merger_135_reset = reset;
  assign last_merger_135_io_stream1_valid = last_q_134_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_135_io_stream1_bits = last_q_134_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_135_io_stream2_valid = io_stream_in_136_valid; // @[Stab.scala 177:23]
  assign last_merger_135_io_stream2_bits = io_stream_in_136_bits; // @[Stab.scala 177:23]
  assign last_merger_135_io_result_ready = last_q_135_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_135_clock = clock;
  assign last_q_135_reset = reset;
  assign last_q_135_io_enq_valid = last_merger_135_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_135_io_enq_bits = last_merger_135_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_135_io_deq_ready = last_merger_136_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_136_clock = clock;
  assign last_merger_136_reset = reset;
  assign last_merger_136_io_stream1_valid = last_q_135_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_136_io_stream1_bits = last_q_135_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_136_io_stream2_valid = io_stream_in_137_valid; // @[Stab.scala 177:23]
  assign last_merger_136_io_stream2_bits = io_stream_in_137_bits; // @[Stab.scala 177:23]
  assign last_merger_136_io_result_ready = last_q_136_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_136_clock = clock;
  assign last_q_136_reset = reset;
  assign last_q_136_io_enq_valid = last_merger_136_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_136_io_enq_bits = last_merger_136_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_136_io_deq_ready = last_merger_137_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_137_clock = clock;
  assign last_merger_137_reset = reset;
  assign last_merger_137_io_stream1_valid = last_q_136_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_137_io_stream1_bits = last_q_136_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_137_io_stream2_valid = io_stream_in_138_valid; // @[Stab.scala 177:23]
  assign last_merger_137_io_stream2_bits = io_stream_in_138_bits; // @[Stab.scala 177:23]
  assign last_merger_137_io_result_ready = last_q_137_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_137_clock = clock;
  assign last_q_137_reset = reset;
  assign last_q_137_io_enq_valid = last_merger_137_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_137_io_enq_bits = last_merger_137_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_137_io_deq_ready = last_merger_138_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_138_clock = clock;
  assign last_merger_138_reset = reset;
  assign last_merger_138_io_stream1_valid = last_q_137_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_138_io_stream1_bits = last_q_137_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_138_io_stream2_valid = io_stream_in_139_valid; // @[Stab.scala 177:23]
  assign last_merger_138_io_stream2_bits = io_stream_in_139_bits; // @[Stab.scala 177:23]
  assign last_merger_138_io_result_ready = last_q_138_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_138_clock = clock;
  assign last_q_138_reset = reset;
  assign last_q_138_io_enq_valid = last_merger_138_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_138_io_enq_bits = last_merger_138_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_138_io_deq_ready = last_merger_139_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_139_clock = clock;
  assign last_merger_139_reset = reset;
  assign last_merger_139_io_stream1_valid = last_q_138_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_139_io_stream1_bits = last_q_138_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_139_io_stream2_valid = io_stream_in_140_valid; // @[Stab.scala 177:23]
  assign last_merger_139_io_stream2_bits = io_stream_in_140_bits; // @[Stab.scala 177:23]
  assign last_merger_139_io_result_ready = last_q_139_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_139_clock = clock;
  assign last_q_139_reset = reset;
  assign last_q_139_io_enq_valid = last_merger_139_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_139_io_enq_bits = last_merger_139_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_139_io_deq_ready = last_merger_140_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_140_clock = clock;
  assign last_merger_140_reset = reset;
  assign last_merger_140_io_stream1_valid = last_q_139_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_140_io_stream1_bits = last_q_139_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_140_io_stream2_valid = io_stream_in_141_valid; // @[Stab.scala 177:23]
  assign last_merger_140_io_stream2_bits = io_stream_in_141_bits; // @[Stab.scala 177:23]
  assign last_merger_140_io_result_ready = last_q_140_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_140_clock = clock;
  assign last_q_140_reset = reset;
  assign last_q_140_io_enq_valid = last_merger_140_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_140_io_enq_bits = last_merger_140_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_140_io_deq_ready = last_merger_141_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_141_clock = clock;
  assign last_merger_141_reset = reset;
  assign last_merger_141_io_stream1_valid = last_q_140_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_141_io_stream1_bits = last_q_140_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_141_io_stream2_valid = io_stream_in_142_valid; // @[Stab.scala 177:23]
  assign last_merger_141_io_stream2_bits = io_stream_in_142_bits; // @[Stab.scala 177:23]
  assign last_merger_141_io_result_ready = last_q_141_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_141_clock = clock;
  assign last_q_141_reset = reset;
  assign last_q_141_io_enq_valid = last_merger_141_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_141_io_enq_bits = last_merger_141_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_141_io_deq_ready = last_merger_142_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_142_clock = clock;
  assign last_merger_142_reset = reset;
  assign last_merger_142_io_stream1_valid = last_q_141_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_142_io_stream1_bits = last_q_141_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_142_io_stream2_valid = io_stream_in_143_valid; // @[Stab.scala 177:23]
  assign last_merger_142_io_stream2_bits = io_stream_in_143_bits; // @[Stab.scala 177:23]
  assign last_merger_142_io_result_ready = last_q_142_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_142_clock = clock;
  assign last_q_142_reset = reset;
  assign last_q_142_io_enq_valid = last_merger_142_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_142_io_enq_bits = last_merger_142_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_142_io_deq_ready = last_merger_143_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_143_clock = clock;
  assign last_merger_143_reset = reset;
  assign last_merger_143_io_stream1_valid = last_q_142_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_143_io_stream1_bits = last_q_142_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_143_io_stream2_valid = io_stream_in_144_valid; // @[Stab.scala 177:23]
  assign last_merger_143_io_stream2_bits = io_stream_in_144_bits; // @[Stab.scala 177:23]
  assign last_merger_143_io_result_ready = last_q_143_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_143_clock = clock;
  assign last_q_143_reset = reset;
  assign last_q_143_io_enq_valid = last_merger_143_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_143_io_enq_bits = last_merger_143_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_143_io_deq_ready = last_merger_144_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_144_clock = clock;
  assign last_merger_144_reset = reset;
  assign last_merger_144_io_stream1_valid = last_q_143_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_144_io_stream1_bits = last_q_143_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_144_io_stream2_valid = io_stream_in_145_valid; // @[Stab.scala 177:23]
  assign last_merger_144_io_stream2_bits = io_stream_in_145_bits; // @[Stab.scala 177:23]
  assign last_merger_144_io_result_ready = last_q_144_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_144_clock = clock;
  assign last_q_144_reset = reset;
  assign last_q_144_io_enq_valid = last_merger_144_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_144_io_enq_bits = last_merger_144_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_144_io_deq_ready = last_merger_145_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_145_clock = clock;
  assign last_merger_145_reset = reset;
  assign last_merger_145_io_stream1_valid = last_q_144_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_145_io_stream1_bits = last_q_144_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_145_io_stream2_valid = io_stream_in_146_valid; // @[Stab.scala 177:23]
  assign last_merger_145_io_stream2_bits = io_stream_in_146_bits; // @[Stab.scala 177:23]
  assign last_merger_145_io_result_ready = last_q_145_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_145_clock = clock;
  assign last_q_145_reset = reset;
  assign last_q_145_io_enq_valid = last_merger_145_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_145_io_enq_bits = last_merger_145_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_145_io_deq_ready = last_merger_146_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_146_clock = clock;
  assign last_merger_146_reset = reset;
  assign last_merger_146_io_stream1_valid = last_q_145_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_146_io_stream1_bits = last_q_145_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_146_io_stream2_valid = io_stream_in_147_valid; // @[Stab.scala 177:23]
  assign last_merger_146_io_stream2_bits = io_stream_in_147_bits; // @[Stab.scala 177:23]
  assign last_merger_146_io_result_ready = last_q_146_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_146_clock = clock;
  assign last_q_146_reset = reset;
  assign last_q_146_io_enq_valid = last_merger_146_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_146_io_enq_bits = last_merger_146_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_146_io_deq_ready = last_merger_147_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_147_clock = clock;
  assign last_merger_147_reset = reset;
  assign last_merger_147_io_stream1_valid = last_q_146_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_147_io_stream1_bits = last_q_146_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_147_io_stream2_valid = io_stream_in_148_valid; // @[Stab.scala 177:23]
  assign last_merger_147_io_stream2_bits = io_stream_in_148_bits; // @[Stab.scala 177:23]
  assign last_merger_147_io_result_ready = last_q_147_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_147_clock = clock;
  assign last_q_147_reset = reset;
  assign last_q_147_io_enq_valid = last_merger_147_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_147_io_enq_bits = last_merger_147_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_147_io_deq_ready = last_merger_148_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_148_clock = clock;
  assign last_merger_148_reset = reset;
  assign last_merger_148_io_stream1_valid = last_q_147_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_148_io_stream1_bits = last_q_147_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_148_io_stream2_valid = io_stream_in_149_valid; // @[Stab.scala 177:23]
  assign last_merger_148_io_stream2_bits = io_stream_in_149_bits; // @[Stab.scala 177:23]
  assign last_merger_148_io_result_ready = last_q_148_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_148_clock = clock;
  assign last_q_148_reset = reset;
  assign last_q_148_io_enq_valid = last_merger_148_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_148_io_enq_bits = last_merger_148_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_148_io_deq_ready = last_merger_149_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_149_clock = clock;
  assign last_merger_149_reset = reset;
  assign last_merger_149_io_stream1_valid = last_q_148_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_149_io_stream1_bits = last_q_148_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_149_io_stream2_valid = io_stream_in_150_valid; // @[Stab.scala 177:23]
  assign last_merger_149_io_stream2_bits = io_stream_in_150_bits; // @[Stab.scala 177:23]
  assign last_merger_149_io_result_ready = last_q_149_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_149_clock = clock;
  assign last_q_149_reset = reset;
  assign last_q_149_io_enq_valid = last_merger_149_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_149_io_enq_bits = last_merger_149_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_149_io_deq_ready = last_merger_150_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_150_clock = clock;
  assign last_merger_150_reset = reset;
  assign last_merger_150_io_stream1_valid = last_q_149_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_150_io_stream1_bits = last_q_149_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_150_io_stream2_valid = io_stream_in_151_valid; // @[Stab.scala 177:23]
  assign last_merger_150_io_stream2_bits = io_stream_in_151_bits; // @[Stab.scala 177:23]
  assign last_merger_150_io_result_ready = last_q_150_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_150_clock = clock;
  assign last_q_150_reset = reset;
  assign last_q_150_io_enq_valid = last_merger_150_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_150_io_enq_bits = last_merger_150_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_150_io_deq_ready = last_merger_151_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_151_clock = clock;
  assign last_merger_151_reset = reset;
  assign last_merger_151_io_stream1_valid = last_q_150_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_151_io_stream1_bits = last_q_150_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_151_io_stream2_valid = io_stream_in_152_valid; // @[Stab.scala 177:23]
  assign last_merger_151_io_stream2_bits = io_stream_in_152_bits; // @[Stab.scala 177:23]
  assign last_merger_151_io_result_ready = last_q_151_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_151_clock = clock;
  assign last_q_151_reset = reset;
  assign last_q_151_io_enq_valid = last_merger_151_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_151_io_enq_bits = last_merger_151_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_151_io_deq_ready = last_merger_152_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_152_clock = clock;
  assign last_merger_152_reset = reset;
  assign last_merger_152_io_stream1_valid = last_q_151_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_152_io_stream1_bits = last_q_151_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_152_io_stream2_valid = io_stream_in_153_valid; // @[Stab.scala 177:23]
  assign last_merger_152_io_stream2_bits = io_stream_in_153_bits; // @[Stab.scala 177:23]
  assign last_merger_152_io_result_ready = last_q_152_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_152_clock = clock;
  assign last_q_152_reset = reset;
  assign last_q_152_io_enq_valid = last_merger_152_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_152_io_enq_bits = last_merger_152_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_152_io_deq_ready = last_merger_153_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_153_clock = clock;
  assign last_merger_153_reset = reset;
  assign last_merger_153_io_stream1_valid = last_q_152_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_153_io_stream1_bits = last_q_152_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_153_io_stream2_valid = io_stream_in_154_valid; // @[Stab.scala 177:23]
  assign last_merger_153_io_stream2_bits = io_stream_in_154_bits; // @[Stab.scala 177:23]
  assign last_merger_153_io_result_ready = last_q_153_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_153_clock = clock;
  assign last_q_153_reset = reset;
  assign last_q_153_io_enq_valid = last_merger_153_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_153_io_enq_bits = last_merger_153_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_153_io_deq_ready = last_merger_154_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_154_clock = clock;
  assign last_merger_154_reset = reset;
  assign last_merger_154_io_stream1_valid = last_q_153_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_154_io_stream1_bits = last_q_153_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_154_io_stream2_valid = io_stream_in_155_valid; // @[Stab.scala 177:23]
  assign last_merger_154_io_stream2_bits = io_stream_in_155_bits; // @[Stab.scala 177:23]
  assign last_merger_154_io_result_ready = last_q_154_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_154_clock = clock;
  assign last_q_154_reset = reset;
  assign last_q_154_io_enq_valid = last_merger_154_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_154_io_enq_bits = last_merger_154_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_154_io_deq_ready = last_merger_155_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_155_clock = clock;
  assign last_merger_155_reset = reset;
  assign last_merger_155_io_stream1_valid = last_q_154_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_155_io_stream1_bits = last_q_154_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_155_io_stream2_valid = io_stream_in_156_valid; // @[Stab.scala 177:23]
  assign last_merger_155_io_stream2_bits = io_stream_in_156_bits; // @[Stab.scala 177:23]
  assign last_merger_155_io_result_ready = last_q_155_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_155_clock = clock;
  assign last_q_155_reset = reset;
  assign last_q_155_io_enq_valid = last_merger_155_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_155_io_enq_bits = last_merger_155_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_155_io_deq_ready = last_merger_156_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_156_clock = clock;
  assign last_merger_156_reset = reset;
  assign last_merger_156_io_stream1_valid = last_q_155_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_156_io_stream1_bits = last_q_155_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_156_io_stream2_valid = io_stream_in_157_valid; // @[Stab.scala 177:23]
  assign last_merger_156_io_stream2_bits = io_stream_in_157_bits; // @[Stab.scala 177:23]
  assign last_merger_156_io_result_ready = last_q_156_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_156_clock = clock;
  assign last_q_156_reset = reset;
  assign last_q_156_io_enq_valid = last_merger_156_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_156_io_enq_bits = last_merger_156_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_156_io_deq_ready = last_merger_157_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_157_clock = clock;
  assign last_merger_157_reset = reset;
  assign last_merger_157_io_stream1_valid = last_q_156_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_157_io_stream1_bits = last_q_156_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_157_io_stream2_valid = io_stream_in_158_valid; // @[Stab.scala 177:23]
  assign last_merger_157_io_stream2_bits = io_stream_in_158_bits; // @[Stab.scala 177:23]
  assign last_merger_157_io_result_ready = last_q_157_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_157_clock = clock;
  assign last_q_157_reset = reset;
  assign last_q_157_io_enq_valid = last_merger_157_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_157_io_enq_bits = last_merger_157_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_157_io_deq_ready = last_merger_158_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_158_clock = clock;
  assign last_merger_158_reset = reset;
  assign last_merger_158_io_stream1_valid = last_q_157_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_158_io_stream1_bits = last_q_157_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_158_io_stream2_valid = io_stream_in_159_valid; // @[Stab.scala 177:23]
  assign last_merger_158_io_stream2_bits = io_stream_in_159_bits; // @[Stab.scala 177:23]
  assign last_merger_158_io_result_ready = last_q_158_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_158_clock = clock;
  assign last_q_158_reset = reset;
  assign last_q_158_io_enq_valid = last_merger_158_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_158_io_enq_bits = last_merger_158_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_158_io_deq_ready = last_merger_159_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_159_clock = clock;
  assign last_merger_159_reset = reset;
  assign last_merger_159_io_stream1_valid = last_q_158_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_159_io_stream1_bits = last_q_158_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_159_io_stream2_valid = io_stream_in_160_valid; // @[Stab.scala 177:23]
  assign last_merger_159_io_stream2_bits = io_stream_in_160_bits; // @[Stab.scala 177:23]
  assign last_merger_159_io_result_ready = last_q_159_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_159_clock = clock;
  assign last_q_159_reset = reset;
  assign last_q_159_io_enq_valid = last_merger_159_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_159_io_enq_bits = last_merger_159_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_159_io_deq_ready = last_merger_160_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_160_clock = clock;
  assign last_merger_160_reset = reset;
  assign last_merger_160_io_stream1_valid = last_q_159_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_160_io_stream1_bits = last_q_159_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_160_io_stream2_valid = io_stream_in_161_valid; // @[Stab.scala 177:23]
  assign last_merger_160_io_stream2_bits = io_stream_in_161_bits; // @[Stab.scala 177:23]
  assign last_merger_160_io_result_ready = last_q_160_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_160_clock = clock;
  assign last_q_160_reset = reset;
  assign last_q_160_io_enq_valid = last_merger_160_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_160_io_enq_bits = last_merger_160_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_160_io_deq_ready = last_merger_161_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_161_clock = clock;
  assign last_merger_161_reset = reset;
  assign last_merger_161_io_stream1_valid = last_q_160_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_161_io_stream1_bits = last_q_160_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_161_io_stream2_valid = io_stream_in_162_valid; // @[Stab.scala 177:23]
  assign last_merger_161_io_stream2_bits = io_stream_in_162_bits; // @[Stab.scala 177:23]
  assign last_merger_161_io_result_ready = last_q_161_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_161_clock = clock;
  assign last_q_161_reset = reset;
  assign last_q_161_io_enq_valid = last_merger_161_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_161_io_enq_bits = last_merger_161_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_161_io_deq_ready = last_merger_162_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_162_clock = clock;
  assign last_merger_162_reset = reset;
  assign last_merger_162_io_stream1_valid = last_q_161_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_162_io_stream1_bits = last_q_161_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_162_io_stream2_valid = io_stream_in_163_valid; // @[Stab.scala 177:23]
  assign last_merger_162_io_stream2_bits = io_stream_in_163_bits; // @[Stab.scala 177:23]
  assign last_merger_162_io_result_ready = last_q_162_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_162_clock = clock;
  assign last_q_162_reset = reset;
  assign last_q_162_io_enq_valid = last_merger_162_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_162_io_enq_bits = last_merger_162_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_162_io_deq_ready = last_merger_163_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_163_clock = clock;
  assign last_merger_163_reset = reset;
  assign last_merger_163_io_stream1_valid = last_q_162_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_163_io_stream1_bits = last_q_162_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_163_io_stream2_valid = io_stream_in_164_valid; // @[Stab.scala 177:23]
  assign last_merger_163_io_stream2_bits = io_stream_in_164_bits; // @[Stab.scala 177:23]
  assign last_merger_163_io_result_ready = last_q_163_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_163_clock = clock;
  assign last_q_163_reset = reset;
  assign last_q_163_io_enq_valid = last_merger_163_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_163_io_enq_bits = last_merger_163_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_163_io_deq_ready = last_merger_164_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_164_clock = clock;
  assign last_merger_164_reset = reset;
  assign last_merger_164_io_stream1_valid = last_q_163_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_164_io_stream1_bits = last_q_163_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_164_io_stream2_valid = io_stream_in_165_valid; // @[Stab.scala 177:23]
  assign last_merger_164_io_stream2_bits = io_stream_in_165_bits; // @[Stab.scala 177:23]
  assign last_merger_164_io_result_ready = last_q_164_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_164_clock = clock;
  assign last_q_164_reset = reset;
  assign last_q_164_io_enq_valid = last_merger_164_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_164_io_enq_bits = last_merger_164_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_164_io_deq_ready = last_merger_165_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_165_clock = clock;
  assign last_merger_165_reset = reset;
  assign last_merger_165_io_stream1_valid = last_q_164_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_165_io_stream1_bits = last_q_164_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_165_io_stream2_valid = io_stream_in_166_valid; // @[Stab.scala 177:23]
  assign last_merger_165_io_stream2_bits = io_stream_in_166_bits; // @[Stab.scala 177:23]
  assign last_merger_165_io_result_ready = last_q_165_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_165_clock = clock;
  assign last_q_165_reset = reset;
  assign last_q_165_io_enq_valid = last_merger_165_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_165_io_enq_bits = last_merger_165_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_165_io_deq_ready = last_merger_166_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_166_clock = clock;
  assign last_merger_166_reset = reset;
  assign last_merger_166_io_stream1_valid = last_q_165_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_166_io_stream1_bits = last_q_165_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_166_io_stream2_valid = io_stream_in_167_valid; // @[Stab.scala 177:23]
  assign last_merger_166_io_stream2_bits = io_stream_in_167_bits; // @[Stab.scala 177:23]
  assign last_merger_166_io_result_ready = last_q_166_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_166_clock = clock;
  assign last_q_166_reset = reset;
  assign last_q_166_io_enq_valid = last_merger_166_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_166_io_enq_bits = last_merger_166_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_166_io_deq_ready = last_merger_167_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_167_clock = clock;
  assign last_merger_167_reset = reset;
  assign last_merger_167_io_stream1_valid = last_q_166_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_167_io_stream1_bits = last_q_166_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_167_io_stream2_valid = io_stream_in_168_valid; // @[Stab.scala 177:23]
  assign last_merger_167_io_stream2_bits = io_stream_in_168_bits; // @[Stab.scala 177:23]
  assign last_merger_167_io_result_ready = last_q_167_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_167_clock = clock;
  assign last_q_167_reset = reset;
  assign last_q_167_io_enq_valid = last_merger_167_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_167_io_enq_bits = last_merger_167_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_167_io_deq_ready = last_merger_168_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_168_clock = clock;
  assign last_merger_168_reset = reset;
  assign last_merger_168_io_stream1_valid = last_q_167_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_168_io_stream1_bits = last_q_167_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_168_io_stream2_valid = io_stream_in_169_valid; // @[Stab.scala 177:23]
  assign last_merger_168_io_stream2_bits = io_stream_in_169_bits; // @[Stab.scala 177:23]
  assign last_merger_168_io_result_ready = last_q_168_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_168_clock = clock;
  assign last_q_168_reset = reset;
  assign last_q_168_io_enq_valid = last_merger_168_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_168_io_enq_bits = last_merger_168_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_168_io_deq_ready = last_merger_169_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_169_clock = clock;
  assign last_merger_169_reset = reset;
  assign last_merger_169_io_stream1_valid = last_q_168_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_169_io_stream1_bits = last_q_168_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_169_io_stream2_valid = io_stream_in_170_valid; // @[Stab.scala 177:23]
  assign last_merger_169_io_stream2_bits = io_stream_in_170_bits; // @[Stab.scala 177:23]
  assign last_merger_169_io_result_ready = last_q_169_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_169_clock = clock;
  assign last_q_169_reset = reset;
  assign last_q_169_io_enq_valid = last_merger_169_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_169_io_enq_bits = last_merger_169_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_169_io_deq_ready = last_merger_170_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_170_clock = clock;
  assign last_merger_170_reset = reset;
  assign last_merger_170_io_stream1_valid = last_q_169_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_170_io_stream1_bits = last_q_169_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_170_io_stream2_valid = io_stream_in_171_valid; // @[Stab.scala 177:23]
  assign last_merger_170_io_stream2_bits = io_stream_in_171_bits; // @[Stab.scala 177:23]
  assign last_merger_170_io_result_ready = last_q_170_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_170_clock = clock;
  assign last_q_170_reset = reset;
  assign last_q_170_io_enq_valid = last_merger_170_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_170_io_enq_bits = last_merger_170_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_170_io_deq_ready = last_merger_171_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_171_clock = clock;
  assign last_merger_171_reset = reset;
  assign last_merger_171_io_stream1_valid = last_q_170_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_171_io_stream1_bits = last_q_170_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_171_io_stream2_valid = io_stream_in_172_valid; // @[Stab.scala 177:23]
  assign last_merger_171_io_stream2_bits = io_stream_in_172_bits; // @[Stab.scala 177:23]
  assign last_merger_171_io_result_ready = last_q_171_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_171_clock = clock;
  assign last_q_171_reset = reset;
  assign last_q_171_io_enq_valid = last_merger_171_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_171_io_enq_bits = last_merger_171_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_171_io_deq_ready = last_merger_172_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_172_clock = clock;
  assign last_merger_172_reset = reset;
  assign last_merger_172_io_stream1_valid = last_q_171_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_172_io_stream1_bits = last_q_171_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_172_io_stream2_valid = io_stream_in_173_valid; // @[Stab.scala 177:23]
  assign last_merger_172_io_stream2_bits = io_stream_in_173_bits; // @[Stab.scala 177:23]
  assign last_merger_172_io_result_ready = last_q_172_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_172_clock = clock;
  assign last_q_172_reset = reset;
  assign last_q_172_io_enq_valid = last_merger_172_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_172_io_enq_bits = last_merger_172_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_172_io_deq_ready = last_merger_173_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_173_clock = clock;
  assign last_merger_173_reset = reset;
  assign last_merger_173_io_stream1_valid = last_q_172_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_173_io_stream1_bits = last_q_172_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_173_io_stream2_valid = io_stream_in_174_valid; // @[Stab.scala 177:23]
  assign last_merger_173_io_stream2_bits = io_stream_in_174_bits; // @[Stab.scala 177:23]
  assign last_merger_173_io_result_ready = last_q_173_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_173_clock = clock;
  assign last_q_173_reset = reset;
  assign last_q_173_io_enq_valid = last_merger_173_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_173_io_enq_bits = last_merger_173_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_173_io_deq_ready = last_merger_174_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_174_clock = clock;
  assign last_merger_174_reset = reset;
  assign last_merger_174_io_stream1_valid = last_q_173_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_174_io_stream1_bits = last_q_173_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_174_io_stream2_valid = io_stream_in_175_valid; // @[Stab.scala 177:23]
  assign last_merger_174_io_stream2_bits = io_stream_in_175_bits; // @[Stab.scala 177:23]
  assign last_merger_174_io_result_ready = last_q_174_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_174_clock = clock;
  assign last_q_174_reset = reset;
  assign last_q_174_io_enq_valid = last_merger_174_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_174_io_enq_bits = last_merger_174_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_174_io_deq_ready = last_merger_175_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_175_clock = clock;
  assign last_merger_175_reset = reset;
  assign last_merger_175_io_stream1_valid = last_q_174_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_175_io_stream1_bits = last_q_174_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_175_io_stream2_valid = io_stream_in_176_valid; // @[Stab.scala 177:23]
  assign last_merger_175_io_stream2_bits = io_stream_in_176_bits; // @[Stab.scala 177:23]
  assign last_merger_175_io_result_ready = last_q_175_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_175_clock = clock;
  assign last_q_175_reset = reset;
  assign last_q_175_io_enq_valid = last_merger_175_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_175_io_enq_bits = last_merger_175_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_175_io_deq_ready = last_merger_176_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_176_clock = clock;
  assign last_merger_176_reset = reset;
  assign last_merger_176_io_stream1_valid = last_q_175_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_176_io_stream1_bits = last_q_175_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_176_io_stream2_valid = io_stream_in_177_valid; // @[Stab.scala 177:23]
  assign last_merger_176_io_stream2_bits = io_stream_in_177_bits; // @[Stab.scala 177:23]
  assign last_merger_176_io_result_ready = last_q_176_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_176_clock = clock;
  assign last_q_176_reset = reset;
  assign last_q_176_io_enq_valid = last_merger_176_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_176_io_enq_bits = last_merger_176_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_176_io_deq_ready = last_merger_177_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_177_clock = clock;
  assign last_merger_177_reset = reset;
  assign last_merger_177_io_stream1_valid = last_q_176_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_177_io_stream1_bits = last_q_176_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_177_io_stream2_valid = io_stream_in_178_valid; // @[Stab.scala 177:23]
  assign last_merger_177_io_stream2_bits = io_stream_in_178_bits; // @[Stab.scala 177:23]
  assign last_merger_177_io_result_ready = last_q_177_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_177_clock = clock;
  assign last_q_177_reset = reset;
  assign last_q_177_io_enq_valid = last_merger_177_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_177_io_enq_bits = last_merger_177_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_177_io_deq_ready = last_merger_178_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_178_clock = clock;
  assign last_merger_178_reset = reset;
  assign last_merger_178_io_stream1_valid = last_q_177_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_178_io_stream1_bits = last_q_177_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_178_io_stream2_valid = io_stream_in_179_valid; // @[Stab.scala 177:23]
  assign last_merger_178_io_stream2_bits = io_stream_in_179_bits; // @[Stab.scala 177:23]
  assign last_merger_178_io_result_ready = last_q_178_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_178_clock = clock;
  assign last_q_178_reset = reset;
  assign last_q_178_io_enq_valid = last_merger_178_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_178_io_enq_bits = last_merger_178_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_178_io_deq_ready = last_merger_179_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_179_clock = clock;
  assign last_merger_179_reset = reset;
  assign last_merger_179_io_stream1_valid = last_q_178_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_179_io_stream1_bits = last_q_178_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_179_io_stream2_valid = io_stream_in_180_valid; // @[Stab.scala 177:23]
  assign last_merger_179_io_stream2_bits = io_stream_in_180_bits; // @[Stab.scala 177:23]
  assign last_merger_179_io_result_ready = last_q_179_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_179_clock = clock;
  assign last_q_179_reset = reset;
  assign last_q_179_io_enq_valid = last_merger_179_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_179_io_enq_bits = last_merger_179_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_179_io_deq_ready = last_merger_180_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_180_clock = clock;
  assign last_merger_180_reset = reset;
  assign last_merger_180_io_stream1_valid = last_q_179_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_180_io_stream1_bits = last_q_179_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_180_io_stream2_valid = io_stream_in_181_valid; // @[Stab.scala 177:23]
  assign last_merger_180_io_stream2_bits = io_stream_in_181_bits; // @[Stab.scala 177:23]
  assign last_merger_180_io_result_ready = last_q_180_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_180_clock = clock;
  assign last_q_180_reset = reset;
  assign last_q_180_io_enq_valid = last_merger_180_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_180_io_enq_bits = last_merger_180_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_180_io_deq_ready = last_merger_181_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_181_clock = clock;
  assign last_merger_181_reset = reset;
  assign last_merger_181_io_stream1_valid = last_q_180_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_181_io_stream1_bits = last_q_180_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_181_io_stream2_valid = io_stream_in_182_valid; // @[Stab.scala 177:23]
  assign last_merger_181_io_stream2_bits = io_stream_in_182_bits; // @[Stab.scala 177:23]
  assign last_merger_181_io_result_ready = last_q_181_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_181_clock = clock;
  assign last_q_181_reset = reset;
  assign last_q_181_io_enq_valid = last_merger_181_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_181_io_enq_bits = last_merger_181_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_181_io_deq_ready = last_merger_182_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_182_clock = clock;
  assign last_merger_182_reset = reset;
  assign last_merger_182_io_stream1_valid = last_q_181_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_182_io_stream1_bits = last_q_181_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_182_io_stream2_valid = io_stream_in_183_valid; // @[Stab.scala 177:23]
  assign last_merger_182_io_stream2_bits = io_stream_in_183_bits; // @[Stab.scala 177:23]
  assign last_merger_182_io_result_ready = last_q_182_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_182_clock = clock;
  assign last_q_182_reset = reset;
  assign last_q_182_io_enq_valid = last_merger_182_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_182_io_enq_bits = last_merger_182_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_182_io_deq_ready = last_merger_183_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_183_clock = clock;
  assign last_merger_183_reset = reset;
  assign last_merger_183_io_stream1_valid = last_q_182_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_183_io_stream1_bits = last_q_182_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_183_io_stream2_valid = io_stream_in_184_valid; // @[Stab.scala 177:23]
  assign last_merger_183_io_stream2_bits = io_stream_in_184_bits; // @[Stab.scala 177:23]
  assign last_merger_183_io_result_ready = last_q_183_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_183_clock = clock;
  assign last_q_183_reset = reset;
  assign last_q_183_io_enq_valid = last_merger_183_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_183_io_enq_bits = last_merger_183_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_183_io_deq_ready = last_merger_184_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_184_clock = clock;
  assign last_merger_184_reset = reset;
  assign last_merger_184_io_stream1_valid = last_q_183_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_184_io_stream1_bits = last_q_183_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_184_io_stream2_valid = io_stream_in_185_valid; // @[Stab.scala 177:23]
  assign last_merger_184_io_stream2_bits = io_stream_in_185_bits; // @[Stab.scala 177:23]
  assign last_merger_184_io_result_ready = last_q_184_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_184_clock = clock;
  assign last_q_184_reset = reset;
  assign last_q_184_io_enq_valid = last_merger_184_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_184_io_enq_bits = last_merger_184_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_184_io_deq_ready = last_merger_185_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_185_clock = clock;
  assign last_merger_185_reset = reset;
  assign last_merger_185_io_stream1_valid = last_q_184_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_185_io_stream1_bits = last_q_184_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_185_io_stream2_valid = io_stream_in_186_valid; // @[Stab.scala 177:23]
  assign last_merger_185_io_stream2_bits = io_stream_in_186_bits; // @[Stab.scala 177:23]
  assign last_merger_185_io_result_ready = last_q_185_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_185_clock = clock;
  assign last_q_185_reset = reset;
  assign last_q_185_io_enq_valid = last_merger_185_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_185_io_enq_bits = last_merger_185_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_185_io_deq_ready = last_merger_186_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_186_clock = clock;
  assign last_merger_186_reset = reset;
  assign last_merger_186_io_stream1_valid = last_q_185_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_186_io_stream1_bits = last_q_185_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_186_io_stream2_valid = io_stream_in_187_valid; // @[Stab.scala 177:23]
  assign last_merger_186_io_stream2_bits = io_stream_in_187_bits; // @[Stab.scala 177:23]
  assign last_merger_186_io_result_ready = last_q_186_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_186_clock = clock;
  assign last_q_186_reset = reset;
  assign last_q_186_io_enq_valid = last_merger_186_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_186_io_enq_bits = last_merger_186_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_186_io_deq_ready = last_merger_187_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_187_clock = clock;
  assign last_merger_187_reset = reset;
  assign last_merger_187_io_stream1_valid = last_q_186_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_187_io_stream1_bits = last_q_186_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_187_io_stream2_valid = io_stream_in_188_valid; // @[Stab.scala 177:23]
  assign last_merger_187_io_stream2_bits = io_stream_in_188_bits; // @[Stab.scala 177:23]
  assign last_merger_187_io_result_ready = last_q_187_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_187_clock = clock;
  assign last_q_187_reset = reset;
  assign last_q_187_io_enq_valid = last_merger_187_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_187_io_enq_bits = last_merger_187_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_187_io_deq_ready = last_merger_188_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_188_clock = clock;
  assign last_merger_188_reset = reset;
  assign last_merger_188_io_stream1_valid = last_q_187_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_188_io_stream1_bits = last_q_187_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_188_io_stream2_valid = io_stream_in_189_valid; // @[Stab.scala 177:23]
  assign last_merger_188_io_stream2_bits = io_stream_in_189_bits; // @[Stab.scala 177:23]
  assign last_merger_188_io_result_ready = last_q_188_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_188_clock = clock;
  assign last_q_188_reset = reset;
  assign last_q_188_io_enq_valid = last_merger_188_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_188_io_enq_bits = last_merger_188_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_188_io_deq_ready = last_merger_189_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_189_clock = clock;
  assign last_merger_189_reset = reset;
  assign last_merger_189_io_stream1_valid = last_q_188_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_189_io_stream1_bits = last_q_188_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_189_io_stream2_valid = io_stream_in_190_valid; // @[Stab.scala 177:23]
  assign last_merger_189_io_stream2_bits = io_stream_in_190_bits; // @[Stab.scala 177:23]
  assign last_merger_189_io_result_ready = last_q_189_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_189_clock = clock;
  assign last_q_189_reset = reset;
  assign last_q_189_io_enq_valid = last_merger_189_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_189_io_enq_bits = last_merger_189_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_189_io_deq_ready = last_merger_190_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_190_clock = clock;
  assign last_merger_190_reset = reset;
  assign last_merger_190_io_stream1_valid = last_q_189_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_190_io_stream1_bits = last_q_189_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_190_io_stream2_valid = io_stream_in_191_valid; // @[Stab.scala 177:23]
  assign last_merger_190_io_stream2_bits = io_stream_in_191_bits; // @[Stab.scala 177:23]
  assign last_merger_190_io_result_ready = last_q_190_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_190_clock = clock;
  assign last_q_190_reset = reset;
  assign last_q_190_io_enq_valid = last_merger_190_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_190_io_enq_bits = last_merger_190_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_190_io_deq_ready = last_merger_191_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_191_clock = clock;
  assign last_merger_191_reset = reset;
  assign last_merger_191_io_stream1_valid = last_q_190_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_191_io_stream1_bits = last_q_190_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_191_io_stream2_valid = io_stream_in_192_valid; // @[Stab.scala 177:23]
  assign last_merger_191_io_stream2_bits = io_stream_in_192_bits; // @[Stab.scala 177:23]
  assign last_merger_191_io_result_ready = last_q_191_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_191_clock = clock;
  assign last_q_191_reset = reset;
  assign last_q_191_io_enq_valid = last_merger_191_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_191_io_enq_bits = last_merger_191_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_191_io_deq_ready = last_merger_192_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_192_clock = clock;
  assign last_merger_192_reset = reset;
  assign last_merger_192_io_stream1_valid = last_q_191_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_192_io_stream1_bits = last_q_191_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_192_io_stream2_valid = io_stream_in_193_valid; // @[Stab.scala 177:23]
  assign last_merger_192_io_stream2_bits = io_stream_in_193_bits; // @[Stab.scala 177:23]
  assign last_merger_192_io_result_ready = last_q_192_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_192_clock = clock;
  assign last_q_192_reset = reset;
  assign last_q_192_io_enq_valid = last_merger_192_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_192_io_enq_bits = last_merger_192_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_192_io_deq_ready = last_merger_193_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_193_clock = clock;
  assign last_merger_193_reset = reset;
  assign last_merger_193_io_stream1_valid = last_q_192_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_193_io_stream1_bits = last_q_192_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_193_io_stream2_valid = io_stream_in_194_valid; // @[Stab.scala 177:23]
  assign last_merger_193_io_stream2_bits = io_stream_in_194_bits; // @[Stab.scala 177:23]
  assign last_merger_193_io_result_ready = last_q_193_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_193_clock = clock;
  assign last_q_193_reset = reset;
  assign last_q_193_io_enq_valid = last_merger_193_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_193_io_enq_bits = last_merger_193_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_193_io_deq_ready = last_merger_194_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_194_clock = clock;
  assign last_merger_194_reset = reset;
  assign last_merger_194_io_stream1_valid = last_q_193_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_194_io_stream1_bits = last_q_193_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_194_io_stream2_valid = io_stream_in_195_valid; // @[Stab.scala 177:23]
  assign last_merger_194_io_stream2_bits = io_stream_in_195_bits; // @[Stab.scala 177:23]
  assign last_merger_194_io_result_ready = last_q_194_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_194_clock = clock;
  assign last_q_194_reset = reset;
  assign last_q_194_io_enq_valid = last_merger_194_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_194_io_enq_bits = last_merger_194_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_194_io_deq_ready = last_merger_195_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_195_clock = clock;
  assign last_merger_195_reset = reset;
  assign last_merger_195_io_stream1_valid = last_q_194_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_195_io_stream1_bits = last_q_194_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_195_io_stream2_valid = io_stream_in_196_valid; // @[Stab.scala 177:23]
  assign last_merger_195_io_stream2_bits = io_stream_in_196_bits; // @[Stab.scala 177:23]
  assign last_merger_195_io_result_ready = last_q_195_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_195_clock = clock;
  assign last_q_195_reset = reset;
  assign last_q_195_io_enq_valid = last_merger_195_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_195_io_enq_bits = last_merger_195_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_195_io_deq_ready = last_merger_196_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_196_clock = clock;
  assign last_merger_196_reset = reset;
  assign last_merger_196_io_stream1_valid = last_q_195_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_196_io_stream1_bits = last_q_195_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_196_io_stream2_valid = io_stream_in_197_valid; // @[Stab.scala 177:23]
  assign last_merger_196_io_stream2_bits = io_stream_in_197_bits; // @[Stab.scala 177:23]
  assign last_merger_196_io_result_ready = last_q_196_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_196_clock = clock;
  assign last_q_196_reset = reset;
  assign last_q_196_io_enq_valid = last_merger_196_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_196_io_enq_bits = last_merger_196_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_196_io_deq_ready = last_merger_197_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_197_clock = clock;
  assign last_merger_197_reset = reset;
  assign last_merger_197_io_stream1_valid = last_q_196_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_197_io_stream1_bits = last_q_196_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_197_io_stream2_valid = io_stream_in_198_valid; // @[Stab.scala 177:23]
  assign last_merger_197_io_stream2_bits = io_stream_in_198_bits; // @[Stab.scala 177:23]
  assign last_merger_197_io_result_ready = last_q_197_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_197_clock = clock;
  assign last_q_197_reset = reset;
  assign last_q_197_io_enq_valid = last_merger_197_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_197_io_enq_bits = last_merger_197_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_197_io_deq_ready = last_merger_198_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_198_clock = clock;
  assign last_merger_198_reset = reset;
  assign last_merger_198_io_stream1_valid = last_q_197_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_198_io_stream1_bits = last_q_197_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_198_io_stream2_valid = io_stream_in_199_valid; // @[Stab.scala 177:23]
  assign last_merger_198_io_stream2_bits = io_stream_in_199_bits; // @[Stab.scala 177:23]
  assign last_merger_198_io_result_ready = last_q_198_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_198_clock = clock;
  assign last_q_198_reset = reset;
  assign last_q_198_io_enq_valid = last_merger_198_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_198_io_enq_bits = last_merger_198_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_198_io_deq_ready = last_merger_199_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_199_clock = clock;
  assign last_merger_199_reset = reset;
  assign last_merger_199_io_stream1_valid = last_q_198_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_199_io_stream1_bits = last_q_198_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_199_io_stream2_valid = io_stream_in_200_valid; // @[Stab.scala 177:23]
  assign last_merger_199_io_stream2_bits = io_stream_in_200_bits; // @[Stab.scala 177:23]
  assign last_merger_199_io_result_ready = last_q_199_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_199_clock = clock;
  assign last_q_199_reset = reset;
  assign last_q_199_io_enq_valid = last_merger_199_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_199_io_enq_bits = last_merger_199_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_199_io_deq_ready = last_merger_200_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_200_clock = clock;
  assign last_merger_200_reset = reset;
  assign last_merger_200_io_stream1_valid = last_q_199_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_200_io_stream1_bits = last_q_199_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_200_io_stream2_valid = io_stream_in_201_valid; // @[Stab.scala 177:23]
  assign last_merger_200_io_stream2_bits = io_stream_in_201_bits; // @[Stab.scala 177:23]
  assign last_merger_200_io_result_ready = last_q_200_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_200_clock = clock;
  assign last_q_200_reset = reset;
  assign last_q_200_io_enq_valid = last_merger_200_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_200_io_enq_bits = last_merger_200_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_200_io_deq_ready = last_merger_201_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_201_clock = clock;
  assign last_merger_201_reset = reset;
  assign last_merger_201_io_stream1_valid = last_q_200_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_201_io_stream1_bits = last_q_200_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_201_io_stream2_valid = io_stream_in_202_valid; // @[Stab.scala 177:23]
  assign last_merger_201_io_stream2_bits = io_stream_in_202_bits; // @[Stab.scala 177:23]
  assign last_merger_201_io_result_ready = last_q_201_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_201_clock = clock;
  assign last_q_201_reset = reset;
  assign last_q_201_io_enq_valid = last_merger_201_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_201_io_enq_bits = last_merger_201_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_201_io_deq_ready = last_merger_202_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_202_clock = clock;
  assign last_merger_202_reset = reset;
  assign last_merger_202_io_stream1_valid = last_q_201_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_202_io_stream1_bits = last_q_201_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_202_io_stream2_valid = io_stream_in_203_valid; // @[Stab.scala 177:23]
  assign last_merger_202_io_stream2_bits = io_stream_in_203_bits; // @[Stab.scala 177:23]
  assign last_merger_202_io_result_ready = last_q_202_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_202_clock = clock;
  assign last_q_202_reset = reset;
  assign last_q_202_io_enq_valid = last_merger_202_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_202_io_enq_bits = last_merger_202_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_202_io_deq_ready = last_merger_203_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_203_clock = clock;
  assign last_merger_203_reset = reset;
  assign last_merger_203_io_stream1_valid = last_q_202_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_203_io_stream1_bits = last_q_202_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_203_io_stream2_valid = io_stream_in_204_valid; // @[Stab.scala 177:23]
  assign last_merger_203_io_stream2_bits = io_stream_in_204_bits; // @[Stab.scala 177:23]
  assign last_merger_203_io_result_ready = last_q_203_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_203_clock = clock;
  assign last_q_203_reset = reset;
  assign last_q_203_io_enq_valid = last_merger_203_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_203_io_enq_bits = last_merger_203_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_203_io_deq_ready = last_merger_204_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_204_clock = clock;
  assign last_merger_204_reset = reset;
  assign last_merger_204_io_stream1_valid = last_q_203_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_204_io_stream1_bits = last_q_203_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_204_io_stream2_valid = io_stream_in_205_valid; // @[Stab.scala 177:23]
  assign last_merger_204_io_stream2_bits = io_stream_in_205_bits; // @[Stab.scala 177:23]
  assign last_merger_204_io_result_ready = last_q_204_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_204_clock = clock;
  assign last_q_204_reset = reset;
  assign last_q_204_io_enq_valid = last_merger_204_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_204_io_enq_bits = last_merger_204_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_204_io_deq_ready = last_merger_205_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_205_clock = clock;
  assign last_merger_205_reset = reset;
  assign last_merger_205_io_stream1_valid = last_q_204_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_205_io_stream1_bits = last_q_204_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_205_io_stream2_valid = io_stream_in_206_valid; // @[Stab.scala 177:23]
  assign last_merger_205_io_stream2_bits = io_stream_in_206_bits; // @[Stab.scala 177:23]
  assign last_merger_205_io_result_ready = last_q_205_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_205_clock = clock;
  assign last_q_205_reset = reset;
  assign last_q_205_io_enq_valid = last_merger_205_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_205_io_enq_bits = last_merger_205_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_205_io_deq_ready = last_merger_206_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_206_clock = clock;
  assign last_merger_206_reset = reset;
  assign last_merger_206_io_stream1_valid = last_q_205_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_206_io_stream1_bits = last_q_205_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_206_io_stream2_valid = io_stream_in_207_valid; // @[Stab.scala 177:23]
  assign last_merger_206_io_stream2_bits = io_stream_in_207_bits; // @[Stab.scala 177:23]
  assign last_merger_206_io_result_ready = last_q_206_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_206_clock = clock;
  assign last_q_206_reset = reset;
  assign last_q_206_io_enq_valid = last_merger_206_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_206_io_enq_bits = last_merger_206_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_206_io_deq_ready = last_merger_207_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_207_clock = clock;
  assign last_merger_207_reset = reset;
  assign last_merger_207_io_stream1_valid = last_q_206_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_207_io_stream1_bits = last_q_206_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_207_io_stream2_valid = io_stream_in_208_valid; // @[Stab.scala 177:23]
  assign last_merger_207_io_stream2_bits = io_stream_in_208_bits; // @[Stab.scala 177:23]
  assign last_merger_207_io_result_ready = last_q_207_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_207_clock = clock;
  assign last_q_207_reset = reset;
  assign last_q_207_io_enq_valid = last_merger_207_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_207_io_enq_bits = last_merger_207_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_207_io_deq_ready = last_merger_208_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_208_clock = clock;
  assign last_merger_208_reset = reset;
  assign last_merger_208_io_stream1_valid = last_q_207_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_208_io_stream1_bits = last_q_207_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_208_io_stream2_valid = io_stream_in_209_valid; // @[Stab.scala 177:23]
  assign last_merger_208_io_stream2_bits = io_stream_in_209_bits; // @[Stab.scala 177:23]
  assign last_merger_208_io_result_ready = last_q_208_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_208_clock = clock;
  assign last_q_208_reset = reset;
  assign last_q_208_io_enq_valid = last_merger_208_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_208_io_enq_bits = last_merger_208_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_208_io_deq_ready = last_merger_209_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_209_clock = clock;
  assign last_merger_209_reset = reset;
  assign last_merger_209_io_stream1_valid = last_q_208_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_209_io_stream1_bits = last_q_208_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_209_io_stream2_valid = io_stream_in_210_valid; // @[Stab.scala 177:23]
  assign last_merger_209_io_stream2_bits = io_stream_in_210_bits; // @[Stab.scala 177:23]
  assign last_merger_209_io_result_ready = last_q_209_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_209_clock = clock;
  assign last_q_209_reset = reset;
  assign last_q_209_io_enq_valid = last_merger_209_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_209_io_enq_bits = last_merger_209_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_209_io_deq_ready = last_merger_210_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_210_clock = clock;
  assign last_merger_210_reset = reset;
  assign last_merger_210_io_stream1_valid = last_q_209_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_210_io_stream1_bits = last_q_209_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_210_io_stream2_valid = io_stream_in_211_valid; // @[Stab.scala 177:23]
  assign last_merger_210_io_stream2_bits = io_stream_in_211_bits; // @[Stab.scala 177:23]
  assign last_merger_210_io_result_ready = last_q_210_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_210_clock = clock;
  assign last_q_210_reset = reset;
  assign last_q_210_io_enq_valid = last_merger_210_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_210_io_enq_bits = last_merger_210_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_210_io_deq_ready = last_merger_211_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_211_clock = clock;
  assign last_merger_211_reset = reset;
  assign last_merger_211_io_stream1_valid = last_q_210_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_211_io_stream1_bits = last_q_210_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_211_io_stream2_valid = io_stream_in_212_valid; // @[Stab.scala 177:23]
  assign last_merger_211_io_stream2_bits = io_stream_in_212_bits; // @[Stab.scala 177:23]
  assign last_merger_211_io_result_ready = last_q_211_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_211_clock = clock;
  assign last_q_211_reset = reset;
  assign last_q_211_io_enq_valid = last_merger_211_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_211_io_enq_bits = last_merger_211_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_211_io_deq_ready = last_merger_212_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_212_clock = clock;
  assign last_merger_212_reset = reset;
  assign last_merger_212_io_stream1_valid = last_q_211_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_212_io_stream1_bits = last_q_211_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_212_io_stream2_valid = io_stream_in_213_valid; // @[Stab.scala 177:23]
  assign last_merger_212_io_stream2_bits = io_stream_in_213_bits; // @[Stab.scala 177:23]
  assign last_merger_212_io_result_ready = last_q_212_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_212_clock = clock;
  assign last_q_212_reset = reset;
  assign last_q_212_io_enq_valid = last_merger_212_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_212_io_enq_bits = last_merger_212_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_212_io_deq_ready = last_merger_213_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_213_clock = clock;
  assign last_merger_213_reset = reset;
  assign last_merger_213_io_stream1_valid = last_q_212_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_213_io_stream1_bits = last_q_212_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_213_io_stream2_valid = io_stream_in_214_valid; // @[Stab.scala 177:23]
  assign last_merger_213_io_stream2_bits = io_stream_in_214_bits; // @[Stab.scala 177:23]
  assign last_merger_213_io_result_ready = last_q_213_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_213_clock = clock;
  assign last_q_213_reset = reset;
  assign last_q_213_io_enq_valid = last_merger_213_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_213_io_enq_bits = last_merger_213_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_213_io_deq_ready = last_merger_214_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_214_clock = clock;
  assign last_merger_214_reset = reset;
  assign last_merger_214_io_stream1_valid = last_q_213_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_214_io_stream1_bits = last_q_213_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_214_io_stream2_valid = io_stream_in_215_valid; // @[Stab.scala 177:23]
  assign last_merger_214_io_stream2_bits = io_stream_in_215_bits; // @[Stab.scala 177:23]
  assign last_merger_214_io_result_ready = last_q_214_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_214_clock = clock;
  assign last_q_214_reset = reset;
  assign last_q_214_io_enq_valid = last_merger_214_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_214_io_enq_bits = last_merger_214_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_214_io_deq_ready = last_merger_215_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_215_clock = clock;
  assign last_merger_215_reset = reset;
  assign last_merger_215_io_stream1_valid = last_q_214_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_215_io_stream1_bits = last_q_214_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_215_io_stream2_valid = io_stream_in_216_valid; // @[Stab.scala 177:23]
  assign last_merger_215_io_stream2_bits = io_stream_in_216_bits; // @[Stab.scala 177:23]
  assign last_merger_215_io_result_ready = last_q_215_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_215_clock = clock;
  assign last_q_215_reset = reset;
  assign last_q_215_io_enq_valid = last_merger_215_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_215_io_enq_bits = last_merger_215_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_215_io_deq_ready = last_merger_216_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_216_clock = clock;
  assign last_merger_216_reset = reset;
  assign last_merger_216_io_stream1_valid = last_q_215_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_216_io_stream1_bits = last_q_215_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_216_io_stream2_valid = io_stream_in_217_valid; // @[Stab.scala 177:23]
  assign last_merger_216_io_stream2_bits = io_stream_in_217_bits; // @[Stab.scala 177:23]
  assign last_merger_216_io_result_ready = last_q_216_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_216_clock = clock;
  assign last_q_216_reset = reset;
  assign last_q_216_io_enq_valid = last_merger_216_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_216_io_enq_bits = last_merger_216_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_216_io_deq_ready = last_merger_217_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_217_clock = clock;
  assign last_merger_217_reset = reset;
  assign last_merger_217_io_stream1_valid = last_q_216_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_217_io_stream1_bits = last_q_216_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_217_io_stream2_valid = io_stream_in_218_valid; // @[Stab.scala 177:23]
  assign last_merger_217_io_stream2_bits = io_stream_in_218_bits; // @[Stab.scala 177:23]
  assign last_merger_217_io_result_ready = last_q_217_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_217_clock = clock;
  assign last_q_217_reset = reset;
  assign last_q_217_io_enq_valid = last_merger_217_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_217_io_enq_bits = last_merger_217_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_217_io_deq_ready = last_merger_218_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_218_clock = clock;
  assign last_merger_218_reset = reset;
  assign last_merger_218_io_stream1_valid = last_q_217_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_218_io_stream1_bits = last_q_217_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_218_io_stream2_valid = io_stream_in_219_valid; // @[Stab.scala 177:23]
  assign last_merger_218_io_stream2_bits = io_stream_in_219_bits; // @[Stab.scala 177:23]
  assign last_merger_218_io_result_ready = last_q_218_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_218_clock = clock;
  assign last_q_218_reset = reset;
  assign last_q_218_io_enq_valid = last_merger_218_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_218_io_enq_bits = last_merger_218_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_218_io_deq_ready = last_merger_219_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_219_clock = clock;
  assign last_merger_219_reset = reset;
  assign last_merger_219_io_stream1_valid = last_q_218_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_219_io_stream1_bits = last_q_218_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_219_io_stream2_valid = io_stream_in_220_valid; // @[Stab.scala 177:23]
  assign last_merger_219_io_stream2_bits = io_stream_in_220_bits; // @[Stab.scala 177:23]
  assign last_merger_219_io_result_ready = last_q_219_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_219_clock = clock;
  assign last_q_219_reset = reset;
  assign last_q_219_io_enq_valid = last_merger_219_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_219_io_enq_bits = last_merger_219_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_219_io_deq_ready = last_merger_220_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_220_clock = clock;
  assign last_merger_220_reset = reset;
  assign last_merger_220_io_stream1_valid = last_q_219_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_220_io_stream1_bits = last_q_219_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_220_io_stream2_valid = io_stream_in_221_valid; // @[Stab.scala 177:23]
  assign last_merger_220_io_stream2_bits = io_stream_in_221_bits; // @[Stab.scala 177:23]
  assign last_merger_220_io_result_ready = last_q_220_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_220_clock = clock;
  assign last_q_220_reset = reset;
  assign last_q_220_io_enq_valid = last_merger_220_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_220_io_enq_bits = last_merger_220_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_220_io_deq_ready = last_merger_221_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_221_clock = clock;
  assign last_merger_221_reset = reset;
  assign last_merger_221_io_stream1_valid = last_q_220_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_221_io_stream1_bits = last_q_220_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_221_io_stream2_valid = io_stream_in_222_valid; // @[Stab.scala 177:23]
  assign last_merger_221_io_stream2_bits = io_stream_in_222_bits; // @[Stab.scala 177:23]
  assign last_merger_221_io_result_ready = last_q_221_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_221_clock = clock;
  assign last_q_221_reset = reset;
  assign last_q_221_io_enq_valid = last_merger_221_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_221_io_enq_bits = last_merger_221_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_221_io_deq_ready = last_merger_222_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_222_clock = clock;
  assign last_merger_222_reset = reset;
  assign last_merger_222_io_stream1_valid = last_q_221_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_222_io_stream1_bits = last_q_221_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_222_io_stream2_valid = io_stream_in_223_valid; // @[Stab.scala 177:23]
  assign last_merger_222_io_stream2_bits = io_stream_in_223_bits; // @[Stab.scala 177:23]
  assign last_merger_222_io_result_ready = last_q_222_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_222_clock = clock;
  assign last_q_222_reset = reset;
  assign last_q_222_io_enq_valid = last_merger_222_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_222_io_enq_bits = last_merger_222_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_222_io_deq_ready = last_merger_223_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_223_clock = clock;
  assign last_merger_223_reset = reset;
  assign last_merger_223_io_stream1_valid = last_q_222_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_223_io_stream1_bits = last_q_222_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_223_io_stream2_valid = io_stream_in_224_valid; // @[Stab.scala 177:23]
  assign last_merger_223_io_stream2_bits = io_stream_in_224_bits; // @[Stab.scala 177:23]
  assign last_merger_223_io_result_ready = last_q_223_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_223_clock = clock;
  assign last_q_223_reset = reset;
  assign last_q_223_io_enq_valid = last_merger_223_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_223_io_enq_bits = last_merger_223_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_223_io_deq_ready = last_merger_224_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_224_clock = clock;
  assign last_merger_224_reset = reset;
  assign last_merger_224_io_stream1_valid = last_q_223_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_224_io_stream1_bits = last_q_223_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_224_io_stream2_valid = io_stream_in_225_valid; // @[Stab.scala 177:23]
  assign last_merger_224_io_stream2_bits = io_stream_in_225_bits; // @[Stab.scala 177:23]
  assign last_merger_224_io_result_ready = last_q_224_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_224_clock = clock;
  assign last_q_224_reset = reset;
  assign last_q_224_io_enq_valid = last_merger_224_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_224_io_enq_bits = last_merger_224_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_224_io_deq_ready = last_merger_225_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_225_clock = clock;
  assign last_merger_225_reset = reset;
  assign last_merger_225_io_stream1_valid = last_q_224_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_225_io_stream1_bits = last_q_224_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_225_io_stream2_valid = io_stream_in_226_valid; // @[Stab.scala 177:23]
  assign last_merger_225_io_stream2_bits = io_stream_in_226_bits; // @[Stab.scala 177:23]
  assign last_merger_225_io_result_ready = last_q_225_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_225_clock = clock;
  assign last_q_225_reset = reset;
  assign last_q_225_io_enq_valid = last_merger_225_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_225_io_enq_bits = last_merger_225_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_225_io_deq_ready = last_merger_226_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_226_clock = clock;
  assign last_merger_226_reset = reset;
  assign last_merger_226_io_stream1_valid = last_q_225_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_226_io_stream1_bits = last_q_225_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_226_io_stream2_valid = io_stream_in_227_valid; // @[Stab.scala 177:23]
  assign last_merger_226_io_stream2_bits = io_stream_in_227_bits; // @[Stab.scala 177:23]
  assign last_merger_226_io_result_ready = last_q_226_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_226_clock = clock;
  assign last_q_226_reset = reset;
  assign last_q_226_io_enq_valid = last_merger_226_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_226_io_enq_bits = last_merger_226_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_226_io_deq_ready = last_merger_227_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_227_clock = clock;
  assign last_merger_227_reset = reset;
  assign last_merger_227_io_stream1_valid = last_q_226_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_227_io_stream1_bits = last_q_226_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_227_io_stream2_valid = io_stream_in_228_valid; // @[Stab.scala 177:23]
  assign last_merger_227_io_stream2_bits = io_stream_in_228_bits; // @[Stab.scala 177:23]
  assign last_merger_227_io_result_ready = last_q_227_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_227_clock = clock;
  assign last_q_227_reset = reset;
  assign last_q_227_io_enq_valid = last_merger_227_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_227_io_enq_bits = last_merger_227_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_227_io_deq_ready = last_merger_228_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_228_clock = clock;
  assign last_merger_228_reset = reset;
  assign last_merger_228_io_stream1_valid = last_q_227_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_228_io_stream1_bits = last_q_227_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_228_io_stream2_valid = io_stream_in_229_valid; // @[Stab.scala 177:23]
  assign last_merger_228_io_stream2_bits = io_stream_in_229_bits; // @[Stab.scala 177:23]
  assign last_merger_228_io_result_ready = last_q_228_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_228_clock = clock;
  assign last_q_228_reset = reset;
  assign last_q_228_io_enq_valid = last_merger_228_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_228_io_enq_bits = last_merger_228_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_228_io_deq_ready = last_merger_229_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_229_clock = clock;
  assign last_merger_229_reset = reset;
  assign last_merger_229_io_stream1_valid = last_q_228_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_229_io_stream1_bits = last_q_228_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_229_io_stream2_valid = io_stream_in_230_valid; // @[Stab.scala 177:23]
  assign last_merger_229_io_stream2_bits = io_stream_in_230_bits; // @[Stab.scala 177:23]
  assign last_merger_229_io_result_ready = last_q_229_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_229_clock = clock;
  assign last_q_229_reset = reset;
  assign last_q_229_io_enq_valid = last_merger_229_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_229_io_enq_bits = last_merger_229_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_229_io_deq_ready = last_merger_230_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_230_clock = clock;
  assign last_merger_230_reset = reset;
  assign last_merger_230_io_stream1_valid = last_q_229_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_230_io_stream1_bits = last_q_229_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_230_io_stream2_valid = io_stream_in_231_valid; // @[Stab.scala 177:23]
  assign last_merger_230_io_stream2_bits = io_stream_in_231_bits; // @[Stab.scala 177:23]
  assign last_merger_230_io_result_ready = last_q_230_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_230_clock = clock;
  assign last_q_230_reset = reset;
  assign last_q_230_io_enq_valid = last_merger_230_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_230_io_enq_bits = last_merger_230_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_230_io_deq_ready = last_merger_231_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_231_clock = clock;
  assign last_merger_231_reset = reset;
  assign last_merger_231_io_stream1_valid = last_q_230_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_231_io_stream1_bits = last_q_230_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_231_io_stream2_valid = io_stream_in_232_valid; // @[Stab.scala 177:23]
  assign last_merger_231_io_stream2_bits = io_stream_in_232_bits; // @[Stab.scala 177:23]
  assign last_merger_231_io_result_ready = last_q_231_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_231_clock = clock;
  assign last_q_231_reset = reset;
  assign last_q_231_io_enq_valid = last_merger_231_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_231_io_enq_bits = last_merger_231_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_231_io_deq_ready = last_merger_232_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_232_clock = clock;
  assign last_merger_232_reset = reset;
  assign last_merger_232_io_stream1_valid = last_q_231_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_232_io_stream1_bits = last_q_231_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_232_io_stream2_valid = io_stream_in_233_valid; // @[Stab.scala 177:23]
  assign last_merger_232_io_stream2_bits = io_stream_in_233_bits; // @[Stab.scala 177:23]
  assign last_merger_232_io_result_ready = last_q_232_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_232_clock = clock;
  assign last_q_232_reset = reset;
  assign last_q_232_io_enq_valid = last_merger_232_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_232_io_enq_bits = last_merger_232_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_232_io_deq_ready = last_merger_233_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_233_clock = clock;
  assign last_merger_233_reset = reset;
  assign last_merger_233_io_stream1_valid = last_q_232_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_233_io_stream1_bits = last_q_232_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_233_io_stream2_valid = io_stream_in_234_valid; // @[Stab.scala 177:23]
  assign last_merger_233_io_stream2_bits = io_stream_in_234_bits; // @[Stab.scala 177:23]
  assign last_merger_233_io_result_ready = last_q_233_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_233_clock = clock;
  assign last_q_233_reset = reset;
  assign last_q_233_io_enq_valid = last_merger_233_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_233_io_enq_bits = last_merger_233_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_233_io_deq_ready = last_merger_234_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_234_clock = clock;
  assign last_merger_234_reset = reset;
  assign last_merger_234_io_stream1_valid = last_q_233_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_234_io_stream1_bits = last_q_233_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_234_io_stream2_valid = io_stream_in_235_valid; // @[Stab.scala 177:23]
  assign last_merger_234_io_stream2_bits = io_stream_in_235_bits; // @[Stab.scala 177:23]
  assign last_merger_234_io_result_ready = last_q_234_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_234_clock = clock;
  assign last_q_234_reset = reset;
  assign last_q_234_io_enq_valid = last_merger_234_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_234_io_enq_bits = last_merger_234_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_234_io_deq_ready = last_merger_235_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_235_clock = clock;
  assign last_merger_235_reset = reset;
  assign last_merger_235_io_stream1_valid = last_q_234_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_235_io_stream1_bits = last_q_234_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_235_io_stream2_valid = io_stream_in_236_valid; // @[Stab.scala 177:23]
  assign last_merger_235_io_stream2_bits = io_stream_in_236_bits; // @[Stab.scala 177:23]
  assign last_merger_235_io_result_ready = last_q_235_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_235_clock = clock;
  assign last_q_235_reset = reset;
  assign last_q_235_io_enq_valid = last_merger_235_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_235_io_enq_bits = last_merger_235_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_235_io_deq_ready = last_merger_236_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_236_clock = clock;
  assign last_merger_236_reset = reset;
  assign last_merger_236_io_stream1_valid = last_q_235_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_236_io_stream1_bits = last_q_235_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_236_io_stream2_valid = io_stream_in_237_valid; // @[Stab.scala 177:23]
  assign last_merger_236_io_stream2_bits = io_stream_in_237_bits; // @[Stab.scala 177:23]
  assign last_merger_236_io_result_ready = last_q_236_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_236_clock = clock;
  assign last_q_236_reset = reset;
  assign last_q_236_io_enq_valid = last_merger_236_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_236_io_enq_bits = last_merger_236_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_236_io_deq_ready = last_merger_237_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_237_clock = clock;
  assign last_merger_237_reset = reset;
  assign last_merger_237_io_stream1_valid = last_q_236_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_237_io_stream1_bits = last_q_236_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_237_io_stream2_valid = io_stream_in_238_valid; // @[Stab.scala 177:23]
  assign last_merger_237_io_stream2_bits = io_stream_in_238_bits; // @[Stab.scala 177:23]
  assign last_merger_237_io_result_ready = last_q_237_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_237_clock = clock;
  assign last_q_237_reset = reset;
  assign last_q_237_io_enq_valid = last_merger_237_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_237_io_enq_bits = last_merger_237_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_237_io_deq_ready = last_merger_238_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_238_clock = clock;
  assign last_merger_238_reset = reset;
  assign last_merger_238_io_stream1_valid = last_q_237_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_238_io_stream1_bits = last_q_237_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_238_io_stream2_valid = io_stream_in_239_valid; // @[Stab.scala 177:23]
  assign last_merger_238_io_stream2_bits = io_stream_in_239_bits; // @[Stab.scala 177:23]
  assign last_merger_238_io_result_ready = last_q_238_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_238_clock = clock;
  assign last_q_238_reset = reset;
  assign last_q_238_io_enq_valid = last_merger_238_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_238_io_enq_bits = last_merger_238_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_238_io_deq_ready = last_merger_239_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_239_clock = clock;
  assign last_merger_239_reset = reset;
  assign last_merger_239_io_stream1_valid = last_q_238_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_239_io_stream1_bits = last_q_238_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_239_io_stream2_valid = io_stream_in_240_valid; // @[Stab.scala 177:23]
  assign last_merger_239_io_stream2_bits = io_stream_in_240_bits; // @[Stab.scala 177:23]
  assign last_merger_239_io_result_ready = last_q_239_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_239_clock = clock;
  assign last_q_239_reset = reset;
  assign last_q_239_io_enq_valid = last_merger_239_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_239_io_enq_bits = last_merger_239_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_239_io_deq_ready = last_merger_240_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_240_clock = clock;
  assign last_merger_240_reset = reset;
  assign last_merger_240_io_stream1_valid = last_q_239_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_240_io_stream1_bits = last_q_239_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_240_io_stream2_valid = io_stream_in_241_valid; // @[Stab.scala 177:23]
  assign last_merger_240_io_stream2_bits = io_stream_in_241_bits; // @[Stab.scala 177:23]
  assign last_merger_240_io_result_ready = last_q_240_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_240_clock = clock;
  assign last_q_240_reset = reset;
  assign last_q_240_io_enq_valid = last_merger_240_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_240_io_enq_bits = last_merger_240_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_240_io_deq_ready = last_merger_241_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_241_clock = clock;
  assign last_merger_241_reset = reset;
  assign last_merger_241_io_stream1_valid = last_q_240_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_241_io_stream1_bits = last_q_240_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_241_io_stream2_valid = io_stream_in_242_valid; // @[Stab.scala 177:23]
  assign last_merger_241_io_stream2_bits = io_stream_in_242_bits; // @[Stab.scala 177:23]
  assign last_merger_241_io_result_ready = last_q_241_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_241_clock = clock;
  assign last_q_241_reset = reset;
  assign last_q_241_io_enq_valid = last_merger_241_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_241_io_enq_bits = last_merger_241_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_241_io_deq_ready = last_merger_242_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_242_clock = clock;
  assign last_merger_242_reset = reset;
  assign last_merger_242_io_stream1_valid = last_q_241_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_242_io_stream1_bits = last_q_241_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_242_io_stream2_valid = io_stream_in_243_valid; // @[Stab.scala 177:23]
  assign last_merger_242_io_stream2_bits = io_stream_in_243_bits; // @[Stab.scala 177:23]
  assign last_merger_242_io_result_ready = last_q_242_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_242_clock = clock;
  assign last_q_242_reset = reset;
  assign last_q_242_io_enq_valid = last_merger_242_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_242_io_enq_bits = last_merger_242_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_242_io_deq_ready = last_merger_243_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_243_clock = clock;
  assign last_merger_243_reset = reset;
  assign last_merger_243_io_stream1_valid = last_q_242_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_243_io_stream1_bits = last_q_242_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_243_io_stream2_valid = io_stream_in_244_valid; // @[Stab.scala 177:23]
  assign last_merger_243_io_stream2_bits = io_stream_in_244_bits; // @[Stab.scala 177:23]
  assign last_merger_243_io_result_ready = last_q_243_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_243_clock = clock;
  assign last_q_243_reset = reset;
  assign last_q_243_io_enq_valid = last_merger_243_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_243_io_enq_bits = last_merger_243_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_243_io_deq_ready = last_merger_244_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_244_clock = clock;
  assign last_merger_244_reset = reset;
  assign last_merger_244_io_stream1_valid = last_q_243_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_244_io_stream1_bits = last_q_243_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_244_io_stream2_valid = io_stream_in_245_valid; // @[Stab.scala 177:23]
  assign last_merger_244_io_stream2_bits = io_stream_in_245_bits; // @[Stab.scala 177:23]
  assign last_merger_244_io_result_ready = last_q_244_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_244_clock = clock;
  assign last_q_244_reset = reset;
  assign last_q_244_io_enq_valid = last_merger_244_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_244_io_enq_bits = last_merger_244_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_244_io_deq_ready = last_merger_245_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_245_clock = clock;
  assign last_merger_245_reset = reset;
  assign last_merger_245_io_stream1_valid = last_q_244_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_245_io_stream1_bits = last_q_244_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_245_io_stream2_valid = io_stream_in_246_valid; // @[Stab.scala 177:23]
  assign last_merger_245_io_stream2_bits = io_stream_in_246_bits; // @[Stab.scala 177:23]
  assign last_merger_245_io_result_ready = last_q_245_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_245_clock = clock;
  assign last_q_245_reset = reset;
  assign last_q_245_io_enq_valid = last_merger_245_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_245_io_enq_bits = last_merger_245_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_245_io_deq_ready = last_merger_246_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_246_clock = clock;
  assign last_merger_246_reset = reset;
  assign last_merger_246_io_stream1_valid = last_q_245_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_246_io_stream1_bits = last_q_245_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_246_io_stream2_valid = io_stream_in_247_valid; // @[Stab.scala 177:23]
  assign last_merger_246_io_stream2_bits = io_stream_in_247_bits; // @[Stab.scala 177:23]
  assign last_merger_246_io_result_ready = last_q_246_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_246_clock = clock;
  assign last_q_246_reset = reset;
  assign last_q_246_io_enq_valid = last_merger_246_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_246_io_enq_bits = last_merger_246_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_246_io_deq_ready = last_merger_247_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_247_clock = clock;
  assign last_merger_247_reset = reset;
  assign last_merger_247_io_stream1_valid = last_q_246_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_247_io_stream1_bits = last_q_246_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_247_io_stream2_valid = io_stream_in_248_valid; // @[Stab.scala 177:23]
  assign last_merger_247_io_stream2_bits = io_stream_in_248_bits; // @[Stab.scala 177:23]
  assign last_merger_247_io_result_ready = last_q_247_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_247_clock = clock;
  assign last_q_247_reset = reset;
  assign last_q_247_io_enq_valid = last_merger_247_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_247_io_enq_bits = last_merger_247_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_247_io_deq_ready = last_merger_248_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_248_clock = clock;
  assign last_merger_248_reset = reset;
  assign last_merger_248_io_stream1_valid = last_q_247_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_248_io_stream1_bits = last_q_247_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_248_io_stream2_valid = io_stream_in_249_valid; // @[Stab.scala 177:23]
  assign last_merger_248_io_stream2_bits = io_stream_in_249_bits; // @[Stab.scala 177:23]
  assign last_merger_248_io_result_ready = last_q_248_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_248_clock = clock;
  assign last_q_248_reset = reset;
  assign last_q_248_io_enq_valid = last_merger_248_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_248_io_enq_bits = last_merger_248_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_248_io_deq_ready = last_merger_249_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_249_clock = clock;
  assign last_merger_249_reset = reset;
  assign last_merger_249_io_stream1_valid = last_q_248_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_249_io_stream1_bits = last_q_248_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_249_io_stream2_valid = io_stream_in_250_valid; // @[Stab.scala 177:23]
  assign last_merger_249_io_stream2_bits = io_stream_in_250_bits; // @[Stab.scala 177:23]
  assign last_merger_249_io_result_ready = last_q_249_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_249_clock = clock;
  assign last_q_249_reset = reset;
  assign last_q_249_io_enq_valid = last_merger_249_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_249_io_enq_bits = last_merger_249_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_249_io_deq_ready = last_merger_250_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_250_clock = clock;
  assign last_merger_250_reset = reset;
  assign last_merger_250_io_stream1_valid = last_q_249_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_250_io_stream1_bits = last_q_249_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_250_io_stream2_valid = io_stream_in_251_valid; // @[Stab.scala 177:23]
  assign last_merger_250_io_stream2_bits = io_stream_in_251_bits; // @[Stab.scala 177:23]
  assign last_merger_250_io_result_ready = last_q_250_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_250_clock = clock;
  assign last_q_250_reset = reset;
  assign last_q_250_io_enq_valid = last_merger_250_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_250_io_enq_bits = last_merger_250_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_250_io_deq_ready = last_merger_251_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_251_clock = clock;
  assign last_merger_251_reset = reset;
  assign last_merger_251_io_stream1_valid = last_q_250_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_251_io_stream1_bits = last_q_250_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_251_io_stream2_valid = io_stream_in_252_valid; // @[Stab.scala 177:23]
  assign last_merger_251_io_stream2_bits = io_stream_in_252_bits; // @[Stab.scala 177:23]
  assign last_merger_251_io_result_ready = last_q_251_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_251_clock = clock;
  assign last_q_251_reset = reset;
  assign last_q_251_io_enq_valid = last_merger_251_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_251_io_enq_bits = last_merger_251_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_251_io_deq_ready = last_merger_252_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_252_clock = clock;
  assign last_merger_252_reset = reset;
  assign last_merger_252_io_stream1_valid = last_q_251_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_252_io_stream1_bits = last_q_251_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_252_io_stream2_valid = io_stream_in_253_valid; // @[Stab.scala 177:23]
  assign last_merger_252_io_stream2_bits = io_stream_in_253_bits; // @[Stab.scala 177:23]
  assign last_merger_252_io_result_ready = last_q_252_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_252_clock = clock;
  assign last_q_252_reset = reset;
  assign last_q_252_io_enq_valid = last_merger_252_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_252_io_enq_bits = last_merger_252_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_252_io_deq_ready = last_merger_253_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_253_clock = clock;
  assign last_merger_253_reset = reset;
  assign last_merger_253_io_stream1_valid = last_q_252_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_253_io_stream1_bits = last_q_252_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_253_io_stream2_valid = io_stream_in_254_valid; // @[Stab.scala 177:23]
  assign last_merger_253_io_stream2_bits = io_stream_in_254_bits; // @[Stab.scala 177:23]
  assign last_merger_253_io_result_ready = last_q_253_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_q_253_clock = clock;
  assign last_q_253_reset = reset;
  assign last_q_253_io_enq_valid = last_merger_253_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_q_253_io_enq_bits = last_merger_253_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_q_253_io_deq_ready = last_merger_254_io_stream1_ready; // @[Stab.scala 176:23]
  assign last_merger_254_clock = clock;
  assign last_merger_254_reset = reset;
  assign last_merger_254_io_stream1_valid = last_q_253_io_deq_valid; // @[Stab.scala 176:23]
  assign last_merger_254_io_stream1_bits = last_q_253_io_deq_bits; // @[Stab.scala 176:23]
  assign last_merger_254_io_stream2_valid = io_stream_in_255_valid; // @[Stab.scala 177:23]
  assign last_merger_254_io_stream2_bits = io_stream_in_255_bits; // @[Stab.scala 177:23]
  assign last_merger_254_io_result_ready = last_io_enq_ready; // @[Decoupled.scala 365:17]
  assign last_clock = clock;
  assign last_reset = reset;
  assign last_io_enq_valid = last_merger_254_io_result_valid; // @[Decoupled.scala 363:22]
  assign last_io_enq_bits = last_merger_254_io_result_bits; // @[Decoupled.scala 364:21]
  assign last_io_deq_ready = io_stream_out_ready; // @[Stab.scala 180:17]
endmodule
module StreamAggregator(
  input         clock,
  input         reset,
  output        io_stream_in_0_ready,
  input         io_stream_in_0_valid,
  input  [31:0] io_stream_in_0_bits,
  output        io_stream_in_1_ready,
  input         io_stream_in_1_valid,
  input  [31:0] io_stream_in_1_bits,
  output        io_stream_in_2_ready,
  input         io_stream_in_2_valid,
  input  [31:0] io_stream_in_2_bits,
  output        io_stream_in_3_ready,
  input         io_stream_in_3_valid,
  input  [31:0] io_stream_in_3_bits,
  output        io_stream_in_4_ready,
  input         io_stream_in_4_valid,
  input  [31:0] io_stream_in_4_bits,
  output        io_stream_in_5_ready,
  input         io_stream_in_5_valid,
  input  [31:0] io_stream_in_5_bits,
  output        io_stream_in_6_ready,
  input         io_stream_in_6_valid,
  input  [31:0] io_stream_in_6_bits,
  output        io_stream_in_7_ready,
  input         io_stream_in_7_valid,
  input  [31:0] io_stream_in_7_bits,
  output        io_stream_in_8_ready,
  input         io_stream_in_8_valid,
  input  [31:0] io_stream_in_8_bits,
  output        io_stream_in_9_ready,
  input         io_stream_in_9_valid,
  input  [31:0] io_stream_in_9_bits,
  output        io_stream_in_10_ready,
  input         io_stream_in_10_valid,
  input  [31:0] io_stream_in_10_bits,
  output        io_stream_in_11_ready,
  input         io_stream_in_11_valid,
  input  [31:0] io_stream_in_11_bits,
  output        io_stream_in_12_ready,
  input         io_stream_in_12_valid,
  input  [31:0] io_stream_in_12_bits,
  output        io_stream_in_13_ready,
  input         io_stream_in_13_valid,
  input  [31:0] io_stream_in_13_bits,
  output        io_stream_in_14_ready,
  input         io_stream_in_14_valid,
  input  [31:0] io_stream_in_14_bits,
  output        io_stream_in_15_ready,
  input         io_stream_in_15_valid,
  input  [31:0] io_stream_in_15_bits,
  output        io_stream_in_16_ready,
  input         io_stream_in_16_valid,
  input  [31:0] io_stream_in_16_bits,
  output        io_stream_in_17_ready,
  input         io_stream_in_17_valid,
  input  [31:0] io_stream_in_17_bits,
  output        io_stream_in_18_ready,
  input         io_stream_in_18_valid,
  input  [31:0] io_stream_in_18_bits,
  output        io_stream_in_19_ready,
  input         io_stream_in_19_valid,
  input  [31:0] io_stream_in_19_bits,
  output        io_stream_in_20_ready,
  input         io_stream_in_20_valid,
  input  [31:0] io_stream_in_20_bits,
  output        io_stream_in_21_ready,
  input         io_stream_in_21_valid,
  input  [31:0] io_stream_in_21_bits,
  output        io_stream_in_22_ready,
  input         io_stream_in_22_valid,
  input  [31:0] io_stream_in_22_bits,
  output        io_stream_in_23_ready,
  input         io_stream_in_23_valid,
  input  [31:0] io_stream_in_23_bits,
  output        io_stream_in_24_ready,
  input         io_stream_in_24_valid,
  input  [31:0] io_stream_in_24_bits,
  output        io_stream_in_25_ready,
  input         io_stream_in_25_valid,
  input  [31:0] io_stream_in_25_bits,
  output        io_stream_in_26_ready,
  input         io_stream_in_26_valid,
  input  [31:0] io_stream_in_26_bits,
  output        io_stream_in_27_ready,
  input         io_stream_in_27_valid,
  input  [31:0] io_stream_in_27_bits,
  output        io_stream_in_28_ready,
  input         io_stream_in_28_valid,
  input  [31:0] io_stream_in_28_bits,
  output        io_stream_in_29_ready,
  input         io_stream_in_29_valid,
  input  [31:0] io_stream_in_29_bits,
  output        io_stream_in_30_ready,
  input         io_stream_in_30_valid,
  input  [31:0] io_stream_in_30_bits,
  output        io_stream_in_31_ready,
  input         io_stream_in_31_valid,
  input  [31:0] io_stream_in_31_bits,
  output        io_stream_in_32_ready,
  input         io_stream_in_32_valid,
  input  [31:0] io_stream_in_32_bits,
  output        io_stream_in_33_ready,
  input         io_stream_in_33_valid,
  input  [31:0] io_stream_in_33_bits,
  output        io_stream_in_34_ready,
  input         io_stream_in_34_valid,
  input  [31:0] io_stream_in_34_bits,
  output        io_stream_in_35_ready,
  input         io_stream_in_35_valid,
  input  [31:0] io_stream_in_35_bits,
  output        io_stream_in_36_ready,
  input         io_stream_in_36_valid,
  input  [31:0] io_stream_in_36_bits,
  output        io_stream_in_37_ready,
  input         io_stream_in_37_valid,
  input  [31:0] io_stream_in_37_bits,
  output        io_stream_in_38_ready,
  input         io_stream_in_38_valid,
  input  [31:0] io_stream_in_38_bits,
  output        io_stream_in_39_ready,
  input         io_stream_in_39_valid,
  input  [31:0] io_stream_in_39_bits,
  output        io_stream_in_40_ready,
  input         io_stream_in_40_valid,
  input  [31:0] io_stream_in_40_bits,
  output        io_stream_in_41_ready,
  input         io_stream_in_41_valid,
  input  [31:0] io_stream_in_41_bits,
  output        io_stream_in_42_ready,
  input         io_stream_in_42_valid,
  input  [31:0] io_stream_in_42_bits,
  output        io_stream_in_43_ready,
  input         io_stream_in_43_valid,
  input  [31:0] io_stream_in_43_bits,
  output        io_stream_in_44_ready,
  input         io_stream_in_44_valid,
  input  [31:0] io_stream_in_44_bits,
  output        io_stream_in_45_ready,
  input         io_stream_in_45_valid,
  input  [31:0] io_stream_in_45_bits,
  output        io_stream_in_46_ready,
  input         io_stream_in_46_valid,
  input  [31:0] io_stream_in_46_bits,
  output        io_stream_in_47_ready,
  input         io_stream_in_47_valid,
  input  [31:0] io_stream_in_47_bits,
  output        io_stream_in_48_ready,
  input         io_stream_in_48_valid,
  input  [31:0] io_stream_in_48_bits,
  output        io_stream_in_49_ready,
  input         io_stream_in_49_valid,
  input  [31:0] io_stream_in_49_bits,
  output        io_stream_in_50_ready,
  input         io_stream_in_50_valid,
  input  [31:0] io_stream_in_50_bits,
  output        io_stream_in_51_ready,
  input         io_stream_in_51_valid,
  input  [31:0] io_stream_in_51_bits,
  output        io_stream_in_52_ready,
  input         io_stream_in_52_valid,
  input  [31:0] io_stream_in_52_bits,
  output        io_stream_in_53_ready,
  input         io_stream_in_53_valid,
  input  [31:0] io_stream_in_53_bits,
  output        io_stream_in_54_ready,
  input         io_stream_in_54_valid,
  input  [31:0] io_stream_in_54_bits,
  output        io_stream_in_55_ready,
  input         io_stream_in_55_valid,
  input  [31:0] io_stream_in_55_bits,
  output        io_stream_in_56_ready,
  input         io_stream_in_56_valid,
  input  [31:0] io_stream_in_56_bits,
  output        io_stream_in_57_ready,
  input         io_stream_in_57_valid,
  input  [31:0] io_stream_in_57_bits,
  output        io_stream_in_58_ready,
  input         io_stream_in_58_valid,
  input  [31:0] io_stream_in_58_bits,
  output        io_stream_in_59_ready,
  input         io_stream_in_59_valid,
  input  [31:0] io_stream_in_59_bits,
  output        io_stream_in_60_ready,
  input         io_stream_in_60_valid,
  input  [31:0] io_stream_in_60_bits,
  output        io_stream_in_61_ready,
  input         io_stream_in_61_valid,
  input  [31:0] io_stream_in_61_bits,
  output        io_stream_in_62_ready,
  input         io_stream_in_62_valid,
  input  [31:0] io_stream_in_62_bits,
  output        io_stream_in_63_ready,
  input         io_stream_in_63_valid,
  input  [31:0] io_stream_in_63_bits,
  output        io_stream_in_64_ready,
  input         io_stream_in_64_valid,
  input  [31:0] io_stream_in_64_bits,
  output        io_stream_in_65_ready,
  input         io_stream_in_65_valid,
  input  [31:0] io_stream_in_65_bits,
  output        io_stream_in_66_ready,
  input         io_stream_in_66_valid,
  input  [31:0] io_stream_in_66_bits,
  output        io_stream_in_67_ready,
  input         io_stream_in_67_valid,
  input  [31:0] io_stream_in_67_bits,
  output        io_stream_in_68_ready,
  input         io_stream_in_68_valid,
  input  [31:0] io_stream_in_68_bits,
  output        io_stream_in_69_ready,
  input         io_stream_in_69_valid,
  input  [31:0] io_stream_in_69_bits,
  output        io_stream_in_70_ready,
  input         io_stream_in_70_valid,
  input  [31:0] io_stream_in_70_bits,
  output        io_stream_in_71_ready,
  input         io_stream_in_71_valid,
  input  [31:0] io_stream_in_71_bits,
  output        io_stream_in_72_ready,
  input         io_stream_in_72_valid,
  input  [31:0] io_stream_in_72_bits,
  output        io_stream_in_73_ready,
  input         io_stream_in_73_valid,
  input  [31:0] io_stream_in_73_bits,
  output        io_stream_in_74_ready,
  input         io_stream_in_74_valid,
  input  [31:0] io_stream_in_74_bits,
  output        io_stream_in_75_ready,
  input         io_stream_in_75_valid,
  input  [31:0] io_stream_in_75_bits,
  output        io_stream_in_76_ready,
  input         io_stream_in_76_valid,
  input  [31:0] io_stream_in_76_bits,
  output        io_stream_in_77_ready,
  input         io_stream_in_77_valid,
  input  [31:0] io_stream_in_77_bits,
  output        io_stream_in_78_ready,
  input         io_stream_in_78_valid,
  input  [31:0] io_stream_in_78_bits,
  output        io_stream_in_79_ready,
  input         io_stream_in_79_valid,
  input  [31:0] io_stream_in_79_bits,
  output        io_stream_in_80_ready,
  input         io_stream_in_80_valid,
  input  [31:0] io_stream_in_80_bits,
  output        io_stream_in_81_ready,
  input         io_stream_in_81_valid,
  input  [31:0] io_stream_in_81_bits,
  output        io_stream_in_82_ready,
  input         io_stream_in_82_valid,
  input  [31:0] io_stream_in_82_bits,
  output        io_stream_in_83_ready,
  input         io_stream_in_83_valid,
  input  [31:0] io_stream_in_83_bits,
  output        io_stream_in_84_ready,
  input         io_stream_in_84_valid,
  input  [31:0] io_stream_in_84_bits,
  output        io_stream_in_85_ready,
  input         io_stream_in_85_valid,
  input  [31:0] io_stream_in_85_bits,
  output        io_stream_in_86_ready,
  input         io_stream_in_86_valid,
  input  [31:0] io_stream_in_86_bits,
  output        io_stream_in_87_ready,
  input         io_stream_in_87_valid,
  input  [31:0] io_stream_in_87_bits,
  output        io_stream_in_88_ready,
  input         io_stream_in_88_valid,
  input  [31:0] io_stream_in_88_bits,
  output        io_stream_in_89_ready,
  input         io_stream_in_89_valid,
  input  [31:0] io_stream_in_89_bits,
  output        io_stream_in_90_ready,
  input         io_stream_in_90_valid,
  input  [31:0] io_stream_in_90_bits,
  output        io_stream_in_91_ready,
  input         io_stream_in_91_valid,
  input  [31:0] io_stream_in_91_bits,
  output        io_stream_in_92_ready,
  input         io_stream_in_92_valid,
  input  [31:0] io_stream_in_92_bits,
  output        io_stream_in_93_ready,
  input         io_stream_in_93_valid,
  input  [31:0] io_stream_in_93_bits,
  output        io_stream_in_94_ready,
  input         io_stream_in_94_valid,
  input  [31:0] io_stream_in_94_bits,
  output        io_stream_in_95_ready,
  input         io_stream_in_95_valid,
  input  [31:0] io_stream_in_95_bits,
  output        io_stream_in_96_ready,
  input         io_stream_in_96_valid,
  input  [31:0] io_stream_in_96_bits,
  output        io_stream_in_97_ready,
  input         io_stream_in_97_valid,
  input  [31:0] io_stream_in_97_bits,
  output        io_stream_in_98_ready,
  input         io_stream_in_98_valid,
  input  [31:0] io_stream_in_98_bits,
  output        io_stream_in_99_ready,
  input         io_stream_in_99_valid,
  input  [31:0] io_stream_in_99_bits,
  output        io_stream_in_100_ready,
  input         io_stream_in_100_valid,
  input  [31:0] io_stream_in_100_bits,
  output        io_stream_in_101_ready,
  input         io_stream_in_101_valid,
  input  [31:0] io_stream_in_101_bits,
  output        io_stream_in_102_ready,
  input         io_stream_in_102_valid,
  input  [31:0] io_stream_in_102_bits,
  output        io_stream_in_103_ready,
  input         io_stream_in_103_valid,
  input  [31:0] io_stream_in_103_bits,
  output        io_stream_in_104_ready,
  input         io_stream_in_104_valid,
  input  [31:0] io_stream_in_104_bits,
  output        io_stream_in_105_ready,
  input         io_stream_in_105_valid,
  input  [31:0] io_stream_in_105_bits,
  output        io_stream_in_106_ready,
  input         io_stream_in_106_valid,
  input  [31:0] io_stream_in_106_bits,
  output        io_stream_in_107_ready,
  input         io_stream_in_107_valid,
  input  [31:0] io_stream_in_107_bits,
  output        io_stream_in_108_ready,
  input         io_stream_in_108_valid,
  input  [31:0] io_stream_in_108_bits,
  output        io_stream_in_109_ready,
  input         io_stream_in_109_valid,
  input  [31:0] io_stream_in_109_bits,
  output        io_stream_in_110_ready,
  input         io_stream_in_110_valid,
  input  [31:0] io_stream_in_110_bits,
  output        io_stream_in_111_ready,
  input         io_stream_in_111_valid,
  input  [31:0] io_stream_in_111_bits,
  output        io_stream_in_112_ready,
  input         io_stream_in_112_valid,
  input  [31:0] io_stream_in_112_bits,
  output        io_stream_in_113_ready,
  input         io_stream_in_113_valid,
  input  [31:0] io_stream_in_113_bits,
  output        io_stream_in_114_ready,
  input         io_stream_in_114_valid,
  input  [31:0] io_stream_in_114_bits,
  output        io_stream_in_115_ready,
  input         io_stream_in_115_valid,
  input  [31:0] io_stream_in_115_bits,
  output        io_stream_in_116_ready,
  input         io_stream_in_116_valid,
  input  [31:0] io_stream_in_116_bits,
  output        io_stream_in_117_ready,
  input         io_stream_in_117_valid,
  input  [31:0] io_stream_in_117_bits,
  output        io_stream_in_118_ready,
  input         io_stream_in_118_valid,
  input  [31:0] io_stream_in_118_bits,
  output        io_stream_in_119_ready,
  input         io_stream_in_119_valid,
  input  [31:0] io_stream_in_119_bits,
  output        io_stream_in_120_ready,
  input         io_stream_in_120_valid,
  input  [31:0] io_stream_in_120_bits,
  output        io_stream_in_121_ready,
  input         io_stream_in_121_valid,
  input  [31:0] io_stream_in_121_bits,
  output        io_stream_in_122_ready,
  input         io_stream_in_122_valid,
  input  [31:0] io_stream_in_122_bits,
  output        io_stream_in_123_ready,
  input         io_stream_in_123_valid,
  input  [31:0] io_stream_in_123_bits,
  output        io_stream_in_124_ready,
  input         io_stream_in_124_valid,
  input  [31:0] io_stream_in_124_bits,
  output        io_stream_in_125_ready,
  input         io_stream_in_125_valid,
  input  [31:0] io_stream_in_125_bits,
  output        io_stream_in_126_ready,
  input         io_stream_in_126_valid,
  input  [31:0] io_stream_in_126_bits,
  output        io_stream_in_127_ready,
  input         io_stream_in_127_valid,
  input  [31:0] io_stream_in_127_bits,
  output        io_stream_in_128_ready,
  input         io_stream_in_128_valid,
  input  [31:0] io_stream_in_128_bits,
  output        io_stream_in_129_ready,
  input         io_stream_in_129_valid,
  input  [31:0] io_stream_in_129_bits,
  output        io_stream_in_130_ready,
  input         io_stream_in_130_valid,
  input  [31:0] io_stream_in_130_bits,
  output        io_stream_in_131_ready,
  input         io_stream_in_131_valid,
  input  [31:0] io_stream_in_131_bits,
  output        io_stream_in_132_ready,
  input         io_stream_in_132_valid,
  input  [31:0] io_stream_in_132_bits,
  output        io_stream_in_133_ready,
  input         io_stream_in_133_valid,
  input  [31:0] io_stream_in_133_bits,
  output        io_stream_in_134_ready,
  input         io_stream_in_134_valid,
  input  [31:0] io_stream_in_134_bits,
  output        io_stream_in_135_ready,
  input         io_stream_in_135_valid,
  input  [31:0] io_stream_in_135_bits,
  output        io_stream_in_136_ready,
  input         io_stream_in_136_valid,
  input  [31:0] io_stream_in_136_bits,
  output        io_stream_in_137_ready,
  input         io_stream_in_137_valid,
  input  [31:0] io_stream_in_137_bits,
  output        io_stream_in_138_ready,
  input         io_stream_in_138_valid,
  input  [31:0] io_stream_in_138_bits,
  output        io_stream_in_139_ready,
  input         io_stream_in_139_valid,
  input  [31:0] io_stream_in_139_bits,
  output        io_stream_in_140_ready,
  input         io_stream_in_140_valid,
  input  [31:0] io_stream_in_140_bits,
  output        io_stream_in_141_ready,
  input         io_stream_in_141_valid,
  input  [31:0] io_stream_in_141_bits,
  output        io_stream_in_142_ready,
  input         io_stream_in_142_valid,
  input  [31:0] io_stream_in_142_bits,
  output        io_stream_in_143_ready,
  input         io_stream_in_143_valid,
  input  [31:0] io_stream_in_143_bits,
  output        io_stream_in_144_ready,
  input         io_stream_in_144_valid,
  input  [31:0] io_stream_in_144_bits,
  output        io_stream_in_145_ready,
  input         io_stream_in_145_valid,
  input  [31:0] io_stream_in_145_bits,
  output        io_stream_in_146_ready,
  input         io_stream_in_146_valid,
  input  [31:0] io_stream_in_146_bits,
  output        io_stream_in_147_ready,
  input         io_stream_in_147_valid,
  input  [31:0] io_stream_in_147_bits,
  output        io_stream_in_148_ready,
  input         io_stream_in_148_valid,
  input  [31:0] io_stream_in_148_bits,
  output        io_stream_in_149_ready,
  input         io_stream_in_149_valid,
  input  [31:0] io_stream_in_149_bits,
  output        io_stream_in_150_ready,
  input         io_stream_in_150_valid,
  input  [31:0] io_stream_in_150_bits,
  output        io_stream_in_151_ready,
  input         io_stream_in_151_valid,
  input  [31:0] io_stream_in_151_bits,
  output        io_stream_in_152_ready,
  input         io_stream_in_152_valid,
  input  [31:0] io_stream_in_152_bits,
  output        io_stream_in_153_ready,
  input         io_stream_in_153_valid,
  input  [31:0] io_stream_in_153_bits,
  output        io_stream_in_154_ready,
  input         io_stream_in_154_valid,
  input  [31:0] io_stream_in_154_bits,
  output        io_stream_in_155_ready,
  input         io_stream_in_155_valid,
  input  [31:0] io_stream_in_155_bits,
  output        io_stream_in_156_ready,
  input         io_stream_in_156_valid,
  input  [31:0] io_stream_in_156_bits,
  output        io_stream_in_157_ready,
  input         io_stream_in_157_valid,
  input  [31:0] io_stream_in_157_bits,
  output        io_stream_in_158_ready,
  input         io_stream_in_158_valid,
  input  [31:0] io_stream_in_158_bits,
  output        io_stream_in_159_ready,
  input         io_stream_in_159_valid,
  input  [31:0] io_stream_in_159_bits,
  output        io_stream_in_160_ready,
  input         io_stream_in_160_valid,
  input  [31:0] io_stream_in_160_bits,
  output        io_stream_in_161_ready,
  input         io_stream_in_161_valid,
  input  [31:0] io_stream_in_161_bits,
  output        io_stream_in_162_ready,
  input         io_stream_in_162_valid,
  input  [31:0] io_stream_in_162_bits,
  output        io_stream_in_163_ready,
  input         io_stream_in_163_valid,
  input  [31:0] io_stream_in_163_bits,
  output        io_stream_in_164_ready,
  input         io_stream_in_164_valid,
  input  [31:0] io_stream_in_164_bits,
  output        io_stream_in_165_ready,
  input         io_stream_in_165_valid,
  input  [31:0] io_stream_in_165_bits,
  output        io_stream_in_166_ready,
  input         io_stream_in_166_valid,
  input  [31:0] io_stream_in_166_bits,
  output        io_stream_in_167_ready,
  input         io_stream_in_167_valid,
  input  [31:0] io_stream_in_167_bits,
  output        io_stream_in_168_ready,
  input         io_stream_in_168_valid,
  input  [31:0] io_stream_in_168_bits,
  output        io_stream_in_169_ready,
  input         io_stream_in_169_valid,
  input  [31:0] io_stream_in_169_bits,
  output        io_stream_in_170_ready,
  input         io_stream_in_170_valid,
  input  [31:0] io_stream_in_170_bits,
  output        io_stream_in_171_ready,
  input         io_stream_in_171_valid,
  input  [31:0] io_stream_in_171_bits,
  output        io_stream_in_172_ready,
  input         io_stream_in_172_valid,
  input  [31:0] io_stream_in_172_bits,
  output        io_stream_in_173_ready,
  input         io_stream_in_173_valid,
  input  [31:0] io_stream_in_173_bits,
  output        io_stream_in_174_ready,
  input         io_stream_in_174_valid,
  input  [31:0] io_stream_in_174_bits,
  output        io_stream_in_175_ready,
  input         io_stream_in_175_valid,
  input  [31:0] io_stream_in_175_bits,
  output        io_stream_in_176_ready,
  input         io_stream_in_176_valid,
  input  [31:0] io_stream_in_176_bits,
  output        io_stream_in_177_ready,
  input         io_stream_in_177_valid,
  input  [31:0] io_stream_in_177_bits,
  output        io_stream_in_178_ready,
  input         io_stream_in_178_valid,
  input  [31:0] io_stream_in_178_bits,
  output        io_stream_in_179_ready,
  input         io_stream_in_179_valid,
  input  [31:0] io_stream_in_179_bits,
  output        io_stream_in_180_ready,
  input         io_stream_in_180_valid,
  input  [31:0] io_stream_in_180_bits,
  output        io_stream_in_181_ready,
  input         io_stream_in_181_valid,
  input  [31:0] io_stream_in_181_bits,
  output        io_stream_in_182_ready,
  input         io_stream_in_182_valid,
  input  [31:0] io_stream_in_182_bits,
  output        io_stream_in_183_ready,
  input         io_stream_in_183_valid,
  input  [31:0] io_stream_in_183_bits,
  output        io_stream_in_184_ready,
  input         io_stream_in_184_valid,
  input  [31:0] io_stream_in_184_bits,
  output        io_stream_in_185_ready,
  input         io_stream_in_185_valid,
  input  [31:0] io_stream_in_185_bits,
  output        io_stream_in_186_ready,
  input         io_stream_in_186_valid,
  input  [31:0] io_stream_in_186_bits,
  output        io_stream_in_187_ready,
  input         io_stream_in_187_valid,
  input  [31:0] io_stream_in_187_bits,
  output        io_stream_in_188_ready,
  input         io_stream_in_188_valid,
  input  [31:0] io_stream_in_188_bits,
  output        io_stream_in_189_ready,
  input         io_stream_in_189_valid,
  input  [31:0] io_stream_in_189_bits,
  output        io_stream_in_190_ready,
  input         io_stream_in_190_valid,
  input  [31:0] io_stream_in_190_bits,
  output        io_stream_in_191_ready,
  input         io_stream_in_191_valid,
  input  [31:0] io_stream_in_191_bits,
  output        io_stream_in_192_ready,
  input         io_stream_in_192_valid,
  input  [31:0] io_stream_in_192_bits,
  output        io_stream_in_193_ready,
  input         io_stream_in_193_valid,
  input  [31:0] io_stream_in_193_bits,
  output        io_stream_in_194_ready,
  input         io_stream_in_194_valid,
  input  [31:0] io_stream_in_194_bits,
  output        io_stream_in_195_ready,
  input         io_stream_in_195_valid,
  input  [31:0] io_stream_in_195_bits,
  output        io_stream_in_196_ready,
  input         io_stream_in_196_valid,
  input  [31:0] io_stream_in_196_bits,
  output        io_stream_in_197_ready,
  input         io_stream_in_197_valid,
  input  [31:0] io_stream_in_197_bits,
  output        io_stream_in_198_ready,
  input         io_stream_in_198_valid,
  input  [31:0] io_stream_in_198_bits,
  output        io_stream_in_199_ready,
  input         io_stream_in_199_valid,
  input  [31:0] io_stream_in_199_bits,
  output        io_stream_in_200_ready,
  input         io_stream_in_200_valid,
  input  [31:0] io_stream_in_200_bits,
  output        io_stream_in_201_ready,
  input         io_stream_in_201_valid,
  input  [31:0] io_stream_in_201_bits,
  output        io_stream_in_202_ready,
  input         io_stream_in_202_valid,
  input  [31:0] io_stream_in_202_bits,
  output        io_stream_in_203_ready,
  input         io_stream_in_203_valid,
  input  [31:0] io_stream_in_203_bits,
  output        io_stream_in_204_ready,
  input         io_stream_in_204_valid,
  input  [31:0] io_stream_in_204_bits,
  output        io_stream_in_205_ready,
  input         io_stream_in_205_valid,
  input  [31:0] io_stream_in_205_bits,
  output        io_stream_in_206_ready,
  input         io_stream_in_206_valid,
  input  [31:0] io_stream_in_206_bits,
  output        io_stream_in_207_ready,
  input         io_stream_in_207_valid,
  input  [31:0] io_stream_in_207_bits,
  output        io_stream_in_208_ready,
  input         io_stream_in_208_valid,
  input  [31:0] io_stream_in_208_bits,
  output        io_stream_in_209_ready,
  input         io_stream_in_209_valid,
  input  [31:0] io_stream_in_209_bits,
  output        io_stream_in_210_ready,
  input         io_stream_in_210_valid,
  input  [31:0] io_stream_in_210_bits,
  output        io_stream_in_211_ready,
  input         io_stream_in_211_valid,
  input  [31:0] io_stream_in_211_bits,
  output        io_stream_in_212_ready,
  input         io_stream_in_212_valid,
  input  [31:0] io_stream_in_212_bits,
  output        io_stream_in_213_ready,
  input         io_stream_in_213_valid,
  input  [31:0] io_stream_in_213_bits,
  output        io_stream_in_214_ready,
  input         io_stream_in_214_valid,
  input  [31:0] io_stream_in_214_bits,
  output        io_stream_in_215_ready,
  input         io_stream_in_215_valid,
  input  [31:0] io_stream_in_215_bits,
  output        io_stream_in_216_ready,
  input         io_stream_in_216_valid,
  input  [31:0] io_stream_in_216_bits,
  output        io_stream_in_217_ready,
  input         io_stream_in_217_valid,
  input  [31:0] io_stream_in_217_bits,
  output        io_stream_in_218_ready,
  input         io_stream_in_218_valid,
  input  [31:0] io_stream_in_218_bits,
  output        io_stream_in_219_ready,
  input         io_stream_in_219_valid,
  input  [31:0] io_stream_in_219_bits,
  output        io_stream_in_220_ready,
  input         io_stream_in_220_valid,
  input  [31:0] io_stream_in_220_bits,
  output        io_stream_in_221_ready,
  input         io_stream_in_221_valid,
  input  [31:0] io_stream_in_221_bits,
  output        io_stream_in_222_ready,
  input         io_stream_in_222_valid,
  input  [31:0] io_stream_in_222_bits,
  output        io_stream_in_223_ready,
  input         io_stream_in_223_valid,
  input  [31:0] io_stream_in_223_bits,
  output        io_stream_in_224_ready,
  input         io_stream_in_224_valid,
  input  [31:0] io_stream_in_224_bits,
  output        io_stream_in_225_ready,
  input         io_stream_in_225_valid,
  input  [31:0] io_stream_in_225_bits,
  output        io_stream_in_226_ready,
  input         io_stream_in_226_valid,
  input  [31:0] io_stream_in_226_bits,
  output        io_stream_in_227_ready,
  input         io_stream_in_227_valid,
  input  [31:0] io_stream_in_227_bits,
  output        io_stream_in_228_ready,
  input         io_stream_in_228_valid,
  input  [31:0] io_stream_in_228_bits,
  output        io_stream_in_229_ready,
  input         io_stream_in_229_valid,
  input  [31:0] io_stream_in_229_bits,
  output        io_stream_in_230_ready,
  input         io_stream_in_230_valid,
  input  [31:0] io_stream_in_230_bits,
  output        io_stream_in_231_ready,
  input         io_stream_in_231_valid,
  input  [31:0] io_stream_in_231_bits,
  output        io_stream_in_232_ready,
  input         io_stream_in_232_valid,
  input  [31:0] io_stream_in_232_bits,
  output        io_stream_in_233_ready,
  input         io_stream_in_233_valid,
  input  [31:0] io_stream_in_233_bits,
  output        io_stream_in_234_ready,
  input         io_stream_in_234_valid,
  input  [31:0] io_stream_in_234_bits,
  output        io_stream_in_235_ready,
  input         io_stream_in_235_valid,
  input  [31:0] io_stream_in_235_bits,
  output        io_stream_in_236_ready,
  input         io_stream_in_236_valid,
  input  [31:0] io_stream_in_236_bits,
  output        io_stream_in_237_ready,
  input         io_stream_in_237_valid,
  input  [31:0] io_stream_in_237_bits,
  output        io_stream_in_238_ready,
  input         io_stream_in_238_valid,
  input  [31:0] io_stream_in_238_bits,
  output        io_stream_in_239_ready,
  input         io_stream_in_239_valid,
  input  [31:0] io_stream_in_239_bits,
  output        io_stream_in_240_ready,
  input         io_stream_in_240_valid,
  input  [31:0] io_stream_in_240_bits,
  output        io_stream_in_241_ready,
  input         io_stream_in_241_valid,
  input  [31:0] io_stream_in_241_bits,
  output        io_stream_in_242_ready,
  input         io_stream_in_242_valid,
  input  [31:0] io_stream_in_242_bits,
  output        io_stream_in_243_ready,
  input         io_stream_in_243_valid,
  input  [31:0] io_stream_in_243_bits,
  output        io_stream_in_244_ready,
  input         io_stream_in_244_valid,
  input  [31:0] io_stream_in_244_bits,
  output        io_stream_in_245_ready,
  input         io_stream_in_245_valid,
  input  [31:0] io_stream_in_245_bits,
  output        io_stream_in_246_ready,
  input         io_stream_in_246_valid,
  input  [31:0] io_stream_in_246_bits,
  output        io_stream_in_247_ready,
  input         io_stream_in_247_valid,
  input  [31:0] io_stream_in_247_bits,
  output        io_stream_in_248_ready,
  input         io_stream_in_248_valid,
  input  [31:0] io_stream_in_248_bits,
  output        io_stream_in_249_ready,
  input         io_stream_in_249_valid,
  input  [31:0] io_stream_in_249_bits,
  output        io_stream_in_250_ready,
  input         io_stream_in_250_valid,
  input  [31:0] io_stream_in_250_bits,
  output        io_stream_in_251_ready,
  input         io_stream_in_251_valid,
  input  [31:0] io_stream_in_251_bits,
  output        io_stream_in_252_ready,
  input         io_stream_in_252_valid,
  input  [31:0] io_stream_in_252_bits,
  output        io_stream_in_253_ready,
  input         io_stream_in_253_valid,
  input  [31:0] io_stream_in_253_bits,
  output        io_stream_in_254_ready,
  input         io_stream_in_254_valid,
  input  [31:0] io_stream_in_254_bits,
  output        io_stream_in_255_ready,
  input         io_stream_in_255_valid,
  input  [31:0] io_stream_in_255_bits,
  input         io_stream_out_ready,
  output        io_stream_out_valid,
  output [31:0] io_stream_out_bits
);
  wire  merger_clock; // @[Stab.scala 291:22]
  wire  merger_reset; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_0_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_0_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_0_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_1_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_1_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_1_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_2_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_2_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_2_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_3_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_3_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_3_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_4_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_4_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_4_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_5_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_5_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_5_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_6_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_6_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_6_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_7_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_7_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_7_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_8_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_8_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_8_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_9_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_9_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_9_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_10_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_10_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_10_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_11_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_11_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_11_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_12_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_12_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_12_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_13_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_13_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_13_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_14_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_14_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_14_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_15_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_15_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_15_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_16_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_16_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_16_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_17_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_17_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_17_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_18_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_18_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_18_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_19_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_19_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_19_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_20_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_20_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_20_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_21_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_21_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_21_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_22_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_22_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_22_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_23_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_23_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_23_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_24_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_24_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_24_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_25_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_25_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_25_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_26_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_26_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_26_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_27_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_27_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_27_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_28_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_28_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_28_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_29_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_29_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_29_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_30_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_30_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_30_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_31_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_31_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_31_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_32_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_32_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_32_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_33_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_33_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_33_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_34_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_34_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_34_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_35_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_35_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_35_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_36_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_36_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_36_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_37_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_37_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_37_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_38_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_38_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_38_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_39_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_39_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_39_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_40_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_40_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_40_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_41_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_41_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_41_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_42_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_42_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_42_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_43_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_43_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_43_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_44_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_44_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_44_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_45_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_45_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_45_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_46_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_46_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_46_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_47_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_47_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_47_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_48_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_48_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_48_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_49_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_49_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_49_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_50_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_50_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_50_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_51_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_51_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_51_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_52_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_52_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_52_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_53_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_53_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_53_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_54_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_54_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_54_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_55_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_55_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_55_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_56_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_56_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_56_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_57_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_57_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_57_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_58_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_58_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_58_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_59_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_59_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_59_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_60_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_60_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_60_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_61_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_61_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_61_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_62_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_62_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_62_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_63_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_63_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_63_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_64_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_64_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_64_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_65_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_65_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_65_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_66_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_66_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_66_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_67_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_67_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_67_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_68_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_68_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_68_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_69_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_69_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_69_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_70_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_70_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_70_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_71_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_71_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_71_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_72_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_72_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_72_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_73_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_73_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_73_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_74_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_74_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_74_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_75_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_75_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_75_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_76_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_76_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_76_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_77_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_77_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_77_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_78_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_78_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_78_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_79_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_79_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_79_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_80_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_80_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_80_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_81_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_81_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_81_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_82_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_82_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_82_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_83_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_83_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_83_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_84_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_84_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_84_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_85_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_85_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_85_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_86_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_86_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_86_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_87_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_87_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_87_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_88_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_88_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_88_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_89_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_89_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_89_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_90_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_90_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_90_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_91_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_91_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_91_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_92_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_92_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_92_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_93_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_93_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_93_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_94_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_94_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_94_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_95_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_95_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_95_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_96_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_96_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_96_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_97_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_97_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_97_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_98_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_98_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_98_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_99_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_99_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_99_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_100_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_100_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_100_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_101_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_101_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_101_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_102_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_102_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_102_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_103_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_103_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_103_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_104_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_104_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_104_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_105_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_105_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_105_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_106_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_106_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_106_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_107_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_107_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_107_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_108_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_108_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_108_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_109_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_109_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_109_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_110_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_110_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_110_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_111_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_111_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_111_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_112_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_112_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_112_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_113_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_113_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_113_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_114_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_114_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_114_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_115_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_115_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_115_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_116_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_116_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_116_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_117_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_117_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_117_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_118_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_118_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_118_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_119_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_119_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_119_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_120_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_120_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_120_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_121_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_121_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_121_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_122_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_122_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_122_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_123_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_123_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_123_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_124_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_124_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_124_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_125_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_125_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_125_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_126_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_126_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_126_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_127_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_127_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_127_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_128_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_128_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_128_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_129_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_129_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_129_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_130_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_130_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_130_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_131_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_131_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_131_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_132_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_132_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_132_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_133_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_133_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_133_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_134_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_134_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_134_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_135_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_135_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_135_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_136_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_136_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_136_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_137_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_137_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_137_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_138_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_138_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_138_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_139_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_139_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_139_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_140_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_140_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_140_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_141_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_141_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_141_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_142_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_142_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_142_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_143_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_143_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_143_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_144_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_144_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_144_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_145_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_145_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_145_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_146_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_146_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_146_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_147_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_147_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_147_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_148_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_148_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_148_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_149_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_149_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_149_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_150_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_150_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_150_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_151_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_151_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_151_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_152_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_152_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_152_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_153_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_153_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_153_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_154_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_154_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_154_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_155_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_155_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_155_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_156_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_156_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_156_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_157_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_157_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_157_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_158_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_158_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_158_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_159_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_159_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_159_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_160_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_160_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_160_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_161_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_161_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_161_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_162_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_162_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_162_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_163_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_163_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_163_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_164_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_164_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_164_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_165_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_165_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_165_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_166_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_166_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_166_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_167_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_167_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_167_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_168_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_168_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_168_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_169_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_169_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_169_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_170_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_170_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_170_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_171_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_171_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_171_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_172_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_172_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_172_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_173_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_173_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_173_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_174_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_174_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_174_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_175_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_175_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_175_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_176_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_176_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_176_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_177_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_177_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_177_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_178_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_178_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_178_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_179_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_179_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_179_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_180_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_180_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_180_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_181_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_181_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_181_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_182_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_182_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_182_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_183_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_183_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_183_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_184_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_184_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_184_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_185_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_185_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_185_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_186_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_186_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_186_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_187_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_187_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_187_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_188_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_188_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_188_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_189_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_189_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_189_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_190_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_190_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_190_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_191_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_191_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_191_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_192_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_192_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_192_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_193_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_193_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_193_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_194_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_194_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_194_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_195_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_195_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_195_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_196_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_196_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_196_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_197_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_197_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_197_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_198_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_198_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_198_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_199_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_199_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_199_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_200_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_200_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_200_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_201_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_201_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_201_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_202_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_202_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_202_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_203_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_203_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_203_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_204_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_204_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_204_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_205_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_205_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_205_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_206_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_206_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_206_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_207_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_207_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_207_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_208_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_208_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_208_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_209_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_209_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_209_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_210_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_210_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_210_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_211_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_211_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_211_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_212_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_212_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_212_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_213_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_213_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_213_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_214_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_214_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_214_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_215_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_215_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_215_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_216_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_216_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_216_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_217_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_217_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_217_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_218_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_218_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_218_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_219_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_219_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_219_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_220_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_220_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_220_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_221_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_221_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_221_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_222_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_222_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_222_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_223_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_223_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_223_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_224_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_224_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_224_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_225_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_225_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_225_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_226_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_226_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_226_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_227_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_227_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_227_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_228_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_228_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_228_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_229_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_229_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_229_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_230_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_230_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_230_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_231_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_231_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_231_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_232_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_232_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_232_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_233_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_233_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_233_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_234_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_234_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_234_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_235_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_235_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_235_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_236_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_236_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_236_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_237_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_237_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_237_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_238_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_238_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_238_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_239_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_239_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_239_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_240_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_240_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_240_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_241_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_241_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_241_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_242_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_242_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_242_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_243_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_243_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_243_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_244_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_244_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_244_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_245_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_245_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_245_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_246_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_246_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_246_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_247_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_247_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_247_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_248_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_248_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_248_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_249_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_249_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_249_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_250_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_250_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_250_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_251_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_251_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_251_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_252_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_252_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_252_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_253_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_253_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_253_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_254_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_254_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_254_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_255_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_in_255_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_in_255_bits; // @[Stab.scala 291:22]
  wire  merger_io_stream_out_ready; // @[Stab.scala 291:22]
  wire  merger_io_stream_out_valid; // @[Stab.scala 291:22]
  wire [31:0] merger_io_stream_out_bits; // @[Stab.scala 291:22]
  StreamMergerTree merger ( // @[Stab.scala 291:22]
    .clock(merger_clock),
    .reset(merger_reset),
    .io_stream_in_0_ready(merger_io_stream_in_0_ready),
    .io_stream_in_0_valid(merger_io_stream_in_0_valid),
    .io_stream_in_0_bits(merger_io_stream_in_0_bits),
    .io_stream_in_1_ready(merger_io_stream_in_1_ready),
    .io_stream_in_1_valid(merger_io_stream_in_1_valid),
    .io_stream_in_1_bits(merger_io_stream_in_1_bits),
    .io_stream_in_2_ready(merger_io_stream_in_2_ready),
    .io_stream_in_2_valid(merger_io_stream_in_2_valid),
    .io_stream_in_2_bits(merger_io_stream_in_2_bits),
    .io_stream_in_3_ready(merger_io_stream_in_3_ready),
    .io_stream_in_3_valid(merger_io_stream_in_3_valid),
    .io_stream_in_3_bits(merger_io_stream_in_3_bits),
    .io_stream_in_4_ready(merger_io_stream_in_4_ready),
    .io_stream_in_4_valid(merger_io_stream_in_4_valid),
    .io_stream_in_4_bits(merger_io_stream_in_4_bits),
    .io_stream_in_5_ready(merger_io_stream_in_5_ready),
    .io_stream_in_5_valid(merger_io_stream_in_5_valid),
    .io_stream_in_5_bits(merger_io_stream_in_5_bits),
    .io_stream_in_6_ready(merger_io_stream_in_6_ready),
    .io_stream_in_6_valid(merger_io_stream_in_6_valid),
    .io_stream_in_6_bits(merger_io_stream_in_6_bits),
    .io_stream_in_7_ready(merger_io_stream_in_7_ready),
    .io_stream_in_7_valid(merger_io_stream_in_7_valid),
    .io_stream_in_7_bits(merger_io_stream_in_7_bits),
    .io_stream_in_8_ready(merger_io_stream_in_8_ready),
    .io_stream_in_8_valid(merger_io_stream_in_8_valid),
    .io_stream_in_8_bits(merger_io_stream_in_8_bits),
    .io_stream_in_9_ready(merger_io_stream_in_9_ready),
    .io_stream_in_9_valid(merger_io_stream_in_9_valid),
    .io_stream_in_9_bits(merger_io_stream_in_9_bits),
    .io_stream_in_10_ready(merger_io_stream_in_10_ready),
    .io_stream_in_10_valid(merger_io_stream_in_10_valid),
    .io_stream_in_10_bits(merger_io_stream_in_10_bits),
    .io_stream_in_11_ready(merger_io_stream_in_11_ready),
    .io_stream_in_11_valid(merger_io_stream_in_11_valid),
    .io_stream_in_11_bits(merger_io_stream_in_11_bits),
    .io_stream_in_12_ready(merger_io_stream_in_12_ready),
    .io_stream_in_12_valid(merger_io_stream_in_12_valid),
    .io_stream_in_12_bits(merger_io_stream_in_12_bits),
    .io_stream_in_13_ready(merger_io_stream_in_13_ready),
    .io_stream_in_13_valid(merger_io_stream_in_13_valid),
    .io_stream_in_13_bits(merger_io_stream_in_13_bits),
    .io_stream_in_14_ready(merger_io_stream_in_14_ready),
    .io_stream_in_14_valid(merger_io_stream_in_14_valid),
    .io_stream_in_14_bits(merger_io_stream_in_14_bits),
    .io_stream_in_15_ready(merger_io_stream_in_15_ready),
    .io_stream_in_15_valid(merger_io_stream_in_15_valid),
    .io_stream_in_15_bits(merger_io_stream_in_15_bits),
    .io_stream_in_16_ready(merger_io_stream_in_16_ready),
    .io_stream_in_16_valid(merger_io_stream_in_16_valid),
    .io_stream_in_16_bits(merger_io_stream_in_16_bits),
    .io_stream_in_17_ready(merger_io_stream_in_17_ready),
    .io_stream_in_17_valid(merger_io_stream_in_17_valid),
    .io_stream_in_17_bits(merger_io_stream_in_17_bits),
    .io_stream_in_18_ready(merger_io_stream_in_18_ready),
    .io_stream_in_18_valid(merger_io_stream_in_18_valid),
    .io_stream_in_18_bits(merger_io_stream_in_18_bits),
    .io_stream_in_19_ready(merger_io_stream_in_19_ready),
    .io_stream_in_19_valid(merger_io_stream_in_19_valid),
    .io_stream_in_19_bits(merger_io_stream_in_19_bits),
    .io_stream_in_20_ready(merger_io_stream_in_20_ready),
    .io_stream_in_20_valid(merger_io_stream_in_20_valid),
    .io_stream_in_20_bits(merger_io_stream_in_20_bits),
    .io_stream_in_21_ready(merger_io_stream_in_21_ready),
    .io_stream_in_21_valid(merger_io_stream_in_21_valid),
    .io_stream_in_21_bits(merger_io_stream_in_21_bits),
    .io_stream_in_22_ready(merger_io_stream_in_22_ready),
    .io_stream_in_22_valid(merger_io_stream_in_22_valid),
    .io_stream_in_22_bits(merger_io_stream_in_22_bits),
    .io_stream_in_23_ready(merger_io_stream_in_23_ready),
    .io_stream_in_23_valid(merger_io_stream_in_23_valid),
    .io_stream_in_23_bits(merger_io_stream_in_23_bits),
    .io_stream_in_24_ready(merger_io_stream_in_24_ready),
    .io_stream_in_24_valid(merger_io_stream_in_24_valid),
    .io_stream_in_24_bits(merger_io_stream_in_24_bits),
    .io_stream_in_25_ready(merger_io_stream_in_25_ready),
    .io_stream_in_25_valid(merger_io_stream_in_25_valid),
    .io_stream_in_25_bits(merger_io_stream_in_25_bits),
    .io_stream_in_26_ready(merger_io_stream_in_26_ready),
    .io_stream_in_26_valid(merger_io_stream_in_26_valid),
    .io_stream_in_26_bits(merger_io_stream_in_26_bits),
    .io_stream_in_27_ready(merger_io_stream_in_27_ready),
    .io_stream_in_27_valid(merger_io_stream_in_27_valid),
    .io_stream_in_27_bits(merger_io_stream_in_27_bits),
    .io_stream_in_28_ready(merger_io_stream_in_28_ready),
    .io_stream_in_28_valid(merger_io_stream_in_28_valid),
    .io_stream_in_28_bits(merger_io_stream_in_28_bits),
    .io_stream_in_29_ready(merger_io_stream_in_29_ready),
    .io_stream_in_29_valid(merger_io_stream_in_29_valid),
    .io_stream_in_29_bits(merger_io_stream_in_29_bits),
    .io_stream_in_30_ready(merger_io_stream_in_30_ready),
    .io_stream_in_30_valid(merger_io_stream_in_30_valid),
    .io_stream_in_30_bits(merger_io_stream_in_30_bits),
    .io_stream_in_31_ready(merger_io_stream_in_31_ready),
    .io_stream_in_31_valid(merger_io_stream_in_31_valid),
    .io_stream_in_31_bits(merger_io_stream_in_31_bits),
    .io_stream_in_32_ready(merger_io_stream_in_32_ready),
    .io_stream_in_32_valid(merger_io_stream_in_32_valid),
    .io_stream_in_32_bits(merger_io_stream_in_32_bits),
    .io_stream_in_33_ready(merger_io_stream_in_33_ready),
    .io_stream_in_33_valid(merger_io_stream_in_33_valid),
    .io_stream_in_33_bits(merger_io_stream_in_33_bits),
    .io_stream_in_34_ready(merger_io_stream_in_34_ready),
    .io_stream_in_34_valid(merger_io_stream_in_34_valid),
    .io_stream_in_34_bits(merger_io_stream_in_34_bits),
    .io_stream_in_35_ready(merger_io_stream_in_35_ready),
    .io_stream_in_35_valid(merger_io_stream_in_35_valid),
    .io_stream_in_35_bits(merger_io_stream_in_35_bits),
    .io_stream_in_36_ready(merger_io_stream_in_36_ready),
    .io_stream_in_36_valid(merger_io_stream_in_36_valid),
    .io_stream_in_36_bits(merger_io_stream_in_36_bits),
    .io_stream_in_37_ready(merger_io_stream_in_37_ready),
    .io_stream_in_37_valid(merger_io_stream_in_37_valid),
    .io_stream_in_37_bits(merger_io_stream_in_37_bits),
    .io_stream_in_38_ready(merger_io_stream_in_38_ready),
    .io_stream_in_38_valid(merger_io_stream_in_38_valid),
    .io_stream_in_38_bits(merger_io_stream_in_38_bits),
    .io_stream_in_39_ready(merger_io_stream_in_39_ready),
    .io_stream_in_39_valid(merger_io_stream_in_39_valid),
    .io_stream_in_39_bits(merger_io_stream_in_39_bits),
    .io_stream_in_40_ready(merger_io_stream_in_40_ready),
    .io_stream_in_40_valid(merger_io_stream_in_40_valid),
    .io_stream_in_40_bits(merger_io_stream_in_40_bits),
    .io_stream_in_41_ready(merger_io_stream_in_41_ready),
    .io_stream_in_41_valid(merger_io_stream_in_41_valid),
    .io_stream_in_41_bits(merger_io_stream_in_41_bits),
    .io_stream_in_42_ready(merger_io_stream_in_42_ready),
    .io_stream_in_42_valid(merger_io_stream_in_42_valid),
    .io_stream_in_42_bits(merger_io_stream_in_42_bits),
    .io_stream_in_43_ready(merger_io_stream_in_43_ready),
    .io_stream_in_43_valid(merger_io_stream_in_43_valid),
    .io_stream_in_43_bits(merger_io_stream_in_43_bits),
    .io_stream_in_44_ready(merger_io_stream_in_44_ready),
    .io_stream_in_44_valid(merger_io_stream_in_44_valid),
    .io_stream_in_44_bits(merger_io_stream_in_44_bits),
    .io_stream_in_45_ready(merger_io_stream_in_45_ready),
    .io_stream_in_45_valid(merger_io_stream_in_45_valid),
    .io_stream_in_45_bits(merger_io_stream_in_45_bits),
    .io_stream_in_46_ready(merger_io_stream_in_46_ready),
    .io_stream_in_46_valid(merger_io_stream_in_46_valid),
    .io_stream_in_46_bits(merger_io_stream_in_46_bits),
    .io_stream_in_47_ready(merger_io_stream_in_47_ready),
    .io_stream_in_47_valid(merger_io_stream_in_47_valid),
    .io_stream_in_47_bits(merger_io_stream_in_47_bits),
    .io_stream_in_48_ready(merger_io_stream_in_48_ready),
    .io_stream_in_48_valid(merger_io_stream_in_48_valid),
    .io_stream_in_48_bits(merger_io_stream_in_48_bits),
    .io_stream_in_49_ready(merger_io_stream_in_49_ready),
    .io_stream_in_49_valid(merger_io_stream_in_49_valid),
    .io_stream_in_49_bits(merger_io_stream_in_49_bits),
    .io_stream_in_50_ready(merger_io_stream_in_50_ready),
    .io_stream_in_50_valid(merger_io_stream_in_50_valid),
    .io_stream_in_50_bits(merger_io_stream_in_50_bits),
    .io_stream_in_51_ready(merger_io_stream_in_51_ready),
    .io_stream_in_51_valid(merger_io_stream_in_51_valid),
    .io_stream_in_51_bits(merger_io_stream_in_51_bits),
    .io_stream_in_52_ready(merger_io_stream_in_52_ready),
    .io_stream_in_52_valid(merger_io_stream_in_52_valid),
    .io_stream_in_52_bits(merger_io_stream_in_52_bits),
    .io_stream_in_53_ready(merger_io_stream_in_53_ready),
    .io_stream_in_53_valid(merger_io_stream_in_53_valid),
    .io_stream_in_53_bits(merger_io_stream_in_53_bits),
    .io_stream_in_54_ready(merger_io_stream_in_54_ready),
    .io_stream_in_54_valid(merger_io_stream_in_54_valid),
    .io_stream_in_54_bits(merger_io_stream_in_54_bits),
    .io_stream_in_55_ready(merger_io_stream_in_55_ready),
    .io_stream_in_55_valid(merger_io_stream_in_55_valid),
    .io_stream_in_55_bits(merger_io_stream_in_55_bits),
    .io_stream_in_56_ready(merger_io_stream_in_56_ready),
    .io_stream_in_56_valid(merger_io_stream_in_56_valid),
    .io_stream_in_56_bits(merger_io_stream_in_56_bits),
    .io_stream_in_57_ready(merger_io_stream_in_57_ready),
    .io_stream_in_57_valid(merger_io_stream_in_57_valid),
    .io_stream_in_57_bits(merger_io_stream_in_57_bits),
    .io_stream_in_58_ready(merger_io_stream_in_58_ready),
    .io_stream_in_58_valid(merger_io_stream_in_58_valid),
    .io_stream_in_58_bits(merger_io_stream_in_58_bits),
    .io_stream_in_59_ready(merger_io_stream_in_59_ready),
    .io_stream_in_59_valid(merger_io_stream_in_59_valid),
    .io_stream_in_59_bits(merger_io_stream_in_59_bits),
    .io_stream_in_60_ready(merger_io_stream_in_60_ready),
    .io_stream_in_60_valid(merger_io_stream_in_60_valid),
    .io_stream_in_60_bits(merger_io_stream_in_60_bits),
    .io_stream_in_61_ready(merger_io_stream_in_61_ready),
    .io_stream_in_61_valid(merger_io_stream_in_61_valid),
    .io_stream_in_61_bits(merger_io_stream_in_61_bits),
    .io_stream_in_62_ready(merger_io_stream_in_62_ready),
    .io_stream_in_62_valid(merger_io_stream_in_62_valid),
    .io_stream_in_62_bits(merger_io_stream_in_62_bits),
    .io_stream_in_63_ready(merger_io_stream_in_63_ready),
    .io_stream_in_63_valid(merger_io_stream_in_63_valid),
    .io_stream_in_63_bits(merger_io_stream_in_63_bits),
    .io_stream_in_64_ready(merger_io_stream_in_64_ready),
    .io_stream_in_64_valid(merger_io_stream_in_64_valid),
    .io_stream_in_64_bits(merger_io_stream_in_64_bits),
    .io_stream_in_65_ready(merger_io_stream_in_65_ready),
    .io_stream_in_65_valid(merger_io_stream_in_65_valid),
    .io_stream_in_65_bits(merger_io_stream_in_65_bits),
    .io_stream_in_66_ready(merger_io_stream_in_66_ready),
    .io_stream_in_66_valid(merger_io_stream_in_66_valid),
    .io_stream_in_66_bits(merger_io_stream_in_66_bits),
    .io_stream_in_67_ready(merger_io_stream_in_67_ready),
    .io_stream_in_67_valid(merger_io_stream_in_67_valid),
    .io_stream_in_67_bits(merger_io_stream_in_67_bits),
    .io_stream_in_68_ready(merger_io_stream_in_68_ready),
    .io_stream_in_68_valid(merger_io_stream_in_68_valid),
    .io_stream_in_68_bits(merger_io_stream_in_68_bits),
    .io_stream_in_69_ready(merger_io_stream_in_69_ready),
    .io_stream_in_69_valid(merger_io_stream_in_69_valid),
    .io_stream_in_69_bits(merger_io_stream_in_69_bits),
    .io_stream_in_70_ready(merger_io_stream_in_70_ready),
    .io_stream_in_70_valid(merger_io_stream_in_70_valid),
    .io_stream_in_70_bits(merger_io_stream_in_70_bits),
    .io_stream_in_71_ready(merger_io_stream_in_71_ready),
    .io_stream_in_71_valid(merger_io_stream_in_71_valid),
    .io_stream_in_71_bits(merger_io_stream_in_71_bits),
    .io_stream_in_72_ready(merger_io_stream_in_72_ready),
    .io_stream_in_72_valid(merger_io_stream_in_72_valid),
    .io_stream_in_72_bits(merger_io_stream_in_72_bits),
    .io_stream_in_73_ready(merger_io_stream_in_73_ready),
    .io_stream_in_73_valid(merger_io_stream_in_73_valid),
    .io_stream_in_73_bits(merger_io_stream_in_73_bits),
    .io_stream_in_74_ready(merger_io_stream_in_74_ready),
    .io_stream_in_74_valid(merger_io_stream_in_74_valid),
    .io_stream_in_74_bits(merger_io_stream_in_74_bits),
    .io_stream_in_75_ready(merger_io_stream_in_75_ready),
    .io_stream_in_75_valid(merger_io_stream_in_75_valid),
    .io_stream_in_75_bits(merger_io_stream_in_75_bits),
    .io_stream_in_76_ready(merger_io_stream_in_76_ready),
    .io_stream_in_76_valid(merger_io_stream_in_76_valid),
    .io_stream_in_76_bits(merger_io_stream_in_76_bits),
    .io_stream_in_77_ready(merger_io_stream_in_77_ready),
    .io_stream_in_77_valid(merger_io_stream_in_77_valid),
    .io_stream_in_77_bits(merger_io_stream_in_77_bits),
    .io_stream_in_78_ready(merger_io_stream_in_78_ready),
    .io_stream_in_78_valid(merger_io_stream_in_78_valid),
    .io_stream_in_78_bits(merger_io_stream_in_78_bits),
    .io_stream_in_79_ready(merger_io_stream_in_79_ready),
    .io_stream_in_79_valid(merger_io_stream_in_79_valid),
    .io_stream_in_79_bits(merger_io_stream_in_79_bits),
    .io_stream_in_80_ready(merger_io_stream_in_80_ready),
    .io_stream_in_80_valid(merger_io_stream_in_80_valid),
    .io_stream_in_80_bits(merger_io_stream_in_80_bits),
    .io_stream_in_81_ready(merger_io_stream_in_81_ready),
    .io_stream_in_81_valid(merger_io_stream_in_81_valid),
    .io_stream_in_81_bits(merger_io_stream_in_81_bits),
    .io_stream_in_82_ready(merger_io_stream_in_82_ready),
    .io_stream_in_82_valid(merger_io_stream_in_82_valid),
    .io_stream_in_82_bits(merger_io_stream_in_82_bits),
    .io_stream_in_83_ready(merger_io_stream_in_83_ready),
    .io_stream_in_83_valid(merger_io_stream_in_83_valid),
    .io_stream_in_83_bits(merger_io_stream_in_83_bits),
    .io_stream_in_84_ready(merger_io_stream_in_84_ready),
    .io_stream_in_84_valid(merger_io_stream_in_84_valid),
    .io_stream_in_84_bits(merger_io_stream_in_84_bits),
    .io_stream_in_85_ready(merger_io_stream_in_85_ready),
    .io_stream_in_85_valid(merger_io_stream_in_85_valid),
    .io_stream_in_85_bits(merger_io_stream_in_85_bits),
    .io_stream_in_86_ready(merger_io_stream_in_86_ready),
    .io_stream_in_86_valid(merger_io_stream_in_86_valid),
    .io_stream_in_86_bits(merger_io_stream_in_86_bits),
    .io_stream_in_87_ready(merger_io_stream_in_87_ready),
    .io_stream_in_87_valid(merger_io_stream_in_87_valid),
    .io_stream_in_87_bits(merger_io_stream_in_87_bits),
    .io_stream_in_88_ready(merger_io_stream_in_88_ready),
    .io_stream_in_88_valid(merger_io_stream_in_88_valid),
    .io_stream_in_88_bits(merger_io_stream_in_88_bits),
    .io_stream_in_89_ready(merger_io_stream_in_89_ready),
    .io_stream_in_89_valid(merger_io_stream_in_89_valid),
    .io_stream_in_89_bits(merger_io_stream_in_89_bits),
    .io_stream_in_90_ready(merger_io_stream_in_90_ready),
    .io_stream_in_90_valid(merger_io_stream_in_90_valid),
    .io_stream_in_90_bits(merger_io_stream_in_90_bits),
    .io_stream_in_91_ready(merger_io_stream_in_91_ready),
    .io_stream_in_91_valid(merger_io_stream_in_91_valid),
    .io_stream_in_91_bits(merger_io_stream_in_91_bits),
    .io_stream_in_92_ready(merger_io_stream_in_92_ready),
    .io_stream_in_92_valid(merger_io_stream_in_92_valid),
    .io_stream_in_92_bits(merger_io_stream_in_92_bits),
    .io_stream_in_93_ready(merger_io_stream_in_93_ready),
    .io_stream_in_93_valid(merger_io_stream_in_93_valid),
    .io_stream_in_93_bits(merger_io_stream_in_93_bits),
    .io_stream_in_94_ready(merger_io_stream_in_94_ready),
    .io_stream_in_94_valid(merger_io_stream_in_94_valid),
    .io_stream_in_94_bits(merger_io_stream_in_94_bits),
    .io_stream_in_95_ready(merger_io_stream_in_95_ready),
    .io_stream_in_95_valid(merger_io_stream_in_95_valid),
    .io_stream_in_95_bits(merger_io_stream_in_95_bits),
    .io_stream_in_96_ready(merger_io_stream_in_96_ready),
    .io_stream_in_96_valid(merger_io_stream_in_96_valid),
    .io_stream_in_96_bits(merger_io_stream_in_96_bits),
    .io_stream_in_97_ready(merger_io_stream_in_97_ready),
    .io_stream_in_97_valid(merger_io_stream_in_97_valid),
    .io_stream_in_97_bits(merger_io_stream_in_97_bits),
    .io_stream_in_98_ready(merger_io_stream_in_98_ready),
    .io_stream_in_98_valid(merger_io_stream_in_98_valid),
    .io_stream_in_98_bits(merger_io_stream_in_98_bits),
    .io_stream_in_99_ready(merger_io_stream_in_99_ready),
    .io_stream_in_99_valid(merger_io_stream_in_99_valid),
    .io_stream_in_99_bits(merger_io_stream_in_99_bits),
    .io_stream_in_100_ready(merger_io_stream_in_100_ready),
    .io_stream_in_100_valid(merger_io_stream_in_100_valid),
    .io_stream_in_100_bits(merger_io_stream_in_100_bits),
    .io_stream_in_101_ready(merger_io_stream_in_101_ready),
    .io_stream_in_101_valid(merger_io_stream_in_101_valid),
    .io_stream_in_101_bits(merger_io_stream_in_101_bits),
    .io_stream_in_102_ready(merger_io_stream_in_102_ready),
    .io_stream_in_102_valid(merger_io_stream_in_102_valid),
    .io_stream_in_102_bits(merger_io_stream_in_102_bits),
    .io_stream_in_103_ready(merger_io_stream_in_103_ready),
    .io_stream_in_103_valid(merger_io_stream_in_103_valid),
    .io_stream_in_103_bits(merger_io_stream_in_103_bits),
    .io_stream_in_104_ready(merger_io_stream_in_104_ready),
    .io_stream_in_104_valid(merger_io_stream_in_104_valid),
    .io_stream_in_104_bits(merger_io_stream_in_104_bits),
    .io_stream_in_105_ready(merger_io_stream_in_105_ready),
    .io_stream_in_105_valid(merger_io_stream_in_105_valid),
    .io_stream_in_105_bits(merger_io_stream_in_105_bits),
    .io_stream_in_106_ready(merger_io_stream_in_106_ready),
    .io_stream_in_106_valid(merger_io_stream_in_106_valid),
    .io_stream_in_106_bits(merger_io_stream_in_106_bits),
    .io_stream_in_107_ready(merger_io_stream_in_107_ready),
    .io_stream_in_107_valid(merger_io_stream_in_107_valid),
    .io_stream_in_107_bits(merger_io_stream_in_107_bits),
    .io_stream_in_108_ready(merger_io_stream_in_108_ready),
    .io_stream_in_108_valid(merger_io_stream_in_108_valid),
    .io_stream_in_108_bits(merger_io_stream_in_108_bits),
    .io_stream_in_109_ready(merger_io_stream_in_109_ready),
    .io_stream_in_109_valid(merger_io_stream_in_109_valid),
    .io_stream_in_109_bits(merger_io_stream_in_109_bits),
    .io_stream_in_110_ready(merger_io_stream_in_110_ready),
    .io_stream_in_110_valid(merger_io_stream_in_110_valid),
    .io_stream_in_110_bits(merger_io_stream_in_110_bits),
    .io_stream_in_111_ready(merger_io_stream_in_111_ready),
    .io_stream_in_111_valid(merger_io_stream_in_111_valid),
    .io_stream_in_111_bits(merger_io_stream_in_111_bits),
    .io_stream_in_112_ready(merger_io_stream_in_112_ready),
    .io_stream_in_112_valid(merger_io_stream_in_112_valid),
    .io_stream_in_112_bits(merger_io_stream_in_112_bits),
    .io_stream_in_113_ready(merger_io_stream_in_113_ready),
    .io_stream_in_113_valid(merger_io_stream_in_113_valid),
    .io_stream_in_113_bits(merger_io_stream_in_113_bits),
    .io_stream_in_114_ready(merger_io_stream_in_114_ready),
    .io_stream_in_114_valid(merger_io_stream_in_114_valid),
    .io_stream_in_114_bits(merger_io_stream_in_114_bits),
    .io_stream_in_115_ready(merger_io_stream_in_115_ready),
    .io_stream_in_115_valid(merger_io_stream_in_115_valid),
    .io_stream_in_115_bits(merger_io_stream_in_115_bits),
    .io_stream_in_116_ready(merger_io_stream_in_116_ready),
    .io_stream_in_116_valid(merger_io_stream_in_116_valid),
    .io_stream_in_116_bits(merger_io_stream_in_116_bits),
    .io_stream_in_117_ready(merger_io_stream_in_117_ready),
    .io_stream_in_117_valid(merger_io_stream_in_117_valid),
    .io_stream_in_117_bits(merger_io_stream_in_117_bits),
    .io_stream_in_118_ready(merger_io_stream_in_118_ready),
    .io_stream_in_118_valid(merger_io_stream_in_118_valid),
    .io_stream_in_118_bits(merger_io_stream_in_118_bits),
    .io_stream_in_119_ready(merger_io_stream_in_119_ready),
    .io_stream_in_119_valid(merger_io_stream_in_119_valid),
    .io_stream_in_119_bits(merger_io_stream_in_119_bits),
    .io_stream_in_120_ready(merger_io_stream_in_120_ready),
    .io_stream_in_120_valid(merger_io_stream_in_120_valid),
    .io_stream_in_120_bits(merger_io_stream_in_120_bits),
    .io_stream_in_121_ready(merger_io_stream_in_121_ready),
    .io_stream_in_121_valid(merger_io_stream_in_121_valid),
    .io_stream_in_121_bits(merger_io_stream_in_121_bits),
    .io_stream_in_122_ready(merger_io_stream_in_122_ready),
    .io_stream_in_122_valid(merger_io_stream_in_122_valid),
    .io_stream_in_122_bits(merger_io_stream_in_122_bits),
    .io_stream_in_123_ready(merger_io_stream_in_123_ready),
    .io_stream_in_123_valid(merger_io_stream_in_123_valid),
    .io_stream_in_123_bits(merger_io_stream_in_123_bits),
    .io_stream_in_124_ready(merger_io_stream_in_124_ready),
    .io_stream_in_124_valid(merger_io_stream_in_124_valid),
    .io_stream_in_124_bits(merger_io_stream_in_124_bits),
    .io_stream_in_125_ready(merger_io_stream_in_125_ready),
    .io_stream_in_125_valid(merger_io_stream_in_125_valid),
    .io_stream_in_125_bits(merger_io_stream_in_125_bits),
    .io_stream_in_126_ready(merger_io_stream_in_126_ready),
    .io_stream_in_126_valid(merger_io_stream_in_126_valid),
    .io_stream_in_126_bits(merger_io_stream_in_126_bits),
    .io_stream_in_127_ready(merger_io_stream_in_127_ready),
    .io_stream_in_127_valid(merger_io_stream_in_127_valid),
    .io_stream_in_127_bits(merger_io_stream_in_127_bits),
    .io_stream_in_128_ready(merger_io_stream_in_128_ready),
    .io_stream_in_128_valid(merger_io_stream_in_128_valid),
    .io_stream_in_128_bits(merger_io_stream_in_128_bits),
    .io_stream_in_129_ready(merger_io_stream_in_129_ready),
    .io_stream_in_129_valid(merger_io_stream_in_129_valid),
    .io_stream_in_129_bits(merger_io_stream_in_129_bits),
    .io_stream_in_130_ready(merger_io_stream_in_130_ready),
    .io_stream_in_130_valid(merger_io_stream_in_130_valid),
    .io_stream_in_130_bits(merger_io_stream_in_130_bits),
    .io_stream_in_131_ready(merger_io_stream_in_131_ready),
    .io_stream_in_131_valid(merger_io_stream_in_131_valid),
    .io_stream_in_131_bits(merger_io_stream_in_131_bits),
    .io_stream_in_132_ready(merger_io_stream_in_132_ready),
    .io_stream_in_132_valid(merger_io_stream_in_132_valid),
    .io_stream_in_132_bits(merger_io_stream_in_132_bits),
    .io_stream_in_133_ready(merger_io_stream_in_133_ready),
    .io_stream_in_133_valid(merger_io_stream_in_133_valid),
    .io_stream_in_133_bits(merger_io_stream_in_133_bits),
    .io_stream_in_134_ready(merger_io_stream_in_134_ready),
    .io_stream_in_134_valid(merger_io_stream_in_134_valid),
    .io_stream_in_134_bits(merger_io_stream_in_134_bits),
    .io_stream_in_135_ready(merger_io_stream_in_135_ready),
    .io_stream_in_135_valid(merger_io_stream_in_135_valid),
    .io_stream_in_135_bits(merger_io_stream_in_135_bits),
    .io_stream_in_136_ready(merger_io_stream_in_136_ready),
    .io_stream_in_136_valid(merger_io_stream_in_136_valid),
    .io_stream_in_136_bits(merger_io_stream_in_136_bits),
    .io_stream_in_137_ready(merger_io_stream_in_137_ready),
    .io_stream_in_137_valid(merger_io_stream_in_137_valid),
    .io_stream_in_137_bits(merger_io_stream_in_137_bits),
    .io_stream_in_138_ready(merger_io_stream_in_138_ready),
    .io_stream_in_138_valid(merger_io_stream_in_138_valid),
    .io_stream_in_138_bits(merger_io_stream_in_138_bits),
    .io_stream_in_139_ready(merger_io_stream_in_139_ready),
    .io_stream_in_139_valid(merger_io_stream_in_139_valid),
    .io_stream_in_139_bits(merger_io_stream_in_139_bits),
    .io_stream_in_140_ready(merger_io_stream_in_140_ready),
    .io_stream_in_140_valid(merger_io_stream_in_140_valid),
    .io_stream_in_140_bits(merger_io_stream_in_140_bits),
    .io_stream_in_141_ready(merger_io_stream_in_141_ready),
    .io_stream_in_141_valid(merger_io_stream_in_141_valid),
    .io_stream_in_141_bits(merger_io_stream_in_141_bits),
    .io_stream_in_142_ready(merger_io_stream_in_142_ready),
    .io_stream_in_142_valid(merger_io_stream_in_142_valid),
    .io_stream_in_142_bits(merger_io_stream_in_142_bits),
    .io_stream_in_143_ready(merger_io_stream_in_143_ready),
    .io_stream_in_143_valid(merger_io_stream_in_143_valid),
    .io_stream_in_143_bits(merger_io_stream_in_143_bits),
    .io_stream_in_144_ready(merger_io_stream_in_144_ready),
    .io_stream_in_144_valid(merger_io_stream_in_144_valid),
    .io_stream_in_144_bits(merger_io_stream_in_144_bits),
    .io_stream_in_145_ready(merger_io_stream_in_145_ready),
    .io_stream_in_145_valid(merger_io_stream_in_145_valid),
    .io_stream_in_145_bits(merger_io_stream_in_145_bits),
    .io_stream_in_146_ready(merger_io_stream_in_146_ready),
    .io_stream_in_146_valid(merger_io_stream_in_146_valid),
    .io_stream_in_146_bits(merger_io_stream_in_146_bits),
    .io_stream_in_147_ready(merger_io_stream_in_147_ready),
    .io_stream_in_147_valid(merger_io_stream_in_147_valid),
    .io_stream_in_147_bits(merger_io_stream_in_147_bits),
    .io_stream_in_148_ready(merger_io_stream_in_148_ready),
    .io_stream_in_148_valid(merger_io_stream_in_148_valid),
    .io_stream_in_148_bits(merger_io_stream_in_148_bits),
    .io_stream_in_149_ready(merger_io_stream_in_149_ready),
    .io_stream_in_149_valid(merger_io_stream_in_149_valid),
    .io_stream_in_149_bits(merger_io_stream_in_149_bits),
    .io_stream_in_150_ready(merger_io_stream_in_150_ready),
    .io_stream_in_150_valid(merger_io_stream_in_150_valid),
    .io_stream_in_150_bits(merger_io_stream_in_150_bits),
    .io_stream_in_151_ready(merger_io_stream_in_151_ready),
    .io_stream_in_151_valid(merger_io_stream_in_151_valid),
    .io_stream_in_151_bits(merger_io_stream_in_151_bits),
    .io_stream_in_152_ready(merger_io_stream_in_152_ready),
    .io_stream_in_152_valid(merger_io_stream_in_152_valid),
    .io_stream_in_152_bits(merger_io_stream_in_152_bits),
    .io_stream_in_153_ready(merger_io_stream_in_153_ready),
    .io_stream_in_153_valid(merger_io_stream_in_153_valid),
    .io_stream_in_153_bits(merger_io_stream_in_153_bits),
    .io_stream_in_154_ready(merger_io_stream_in_154_ready),
    .io_stream_in_154_valid(merger_io_stream_in_154_valid),
    .io_stream_in_154_bits(merger_io_stream_in_154_bits),
    .io_stream_in_155_ready(merger_io_stream_in_155_ready),
    .io_stream_in_155_valid(merger_io_stream_in_155_valid),
    .io_stream_in_155_bits(merger_io_stream_in_155_bits),
    .io_stream_in_156_ready(merger_io_stream_in_156_ready),
    .io_stream_in_156_valid(merger_io_stream_in_156_valid),
    .io_stream_in_156_bits(merger_io_stream_in_156_bits),
    .io_stream_in_157_ready(merger_io_stream_in_157_ready),
    .io_stream_in_157_valid(merger_io_stream_in_157_valid),
    .io_stream_in_157_bits(merger_io_stream_in_157_bits),
    .io_stream_in_158_ready(merger_io_stream_in_158_ready),
    .io_stream_in_158_valid(merger_io_stream_in_158_valid),
    .io_stream_in_158_bits(merger_io_stream_in_158_bits),
    .io_stream_in_159_ready(merger_io_stream_in_159_ready),
    .io_stream_in_159_valid(merger_io_stream_in_159_valid),
    .io_stream_in_159_bits(merger_io_stream_in_159_bits),
    .io_stream_in_160_ready(merger_io_stream_in_160_ready),
    .io_stream_in_160_valid(merger_io_stream_in_160_valid),
    .io_stream_in_160_bits(merger_io_stream_in_160_bits),
    .io_stream_in_161_ready(merger_io_stream_in_161_ready),
    .io_stream_in_161_valid(merger_io_stream_in_161_valid),
    .io_stream_in_161_bits(merger_io_stream_in_161_bits),
    .io_stream_in_162_ready(merger_io_stream_in_162_ready),
    .io_stream_in_162_valid(merger_io_stream_in_162_valid),
    .io_stream_in_162_bits(merger_io_stream_in_162_bits),
    .io_stream_in_163_ready(merger_io_stream_in_163_ready),
    .io_stream_in_163_valid(merger_io_stream_in_163_valid),
    .io_stream_in_163_bits(merger_io_stream_in_163_bits),
    .io_stream_in_164_ready(merger_io_stream_in_164_ready),
    .io_stream_in_164_valid(merger_io_stream_in_164_valid),
    .io_stream_in_164_bits(merger_io_stream_in_164_bits),
    .io_stream_in_165_ready(merger_io_stream_in_165_ready),
    .io_stream_in_165_valid(merger_io_stream_in_165_valid),
    .io_stream_in_165_bits(merger_io_stream_in_165_bits),
    .io_stream_in_166_ready(merger_io_stream_in_166_ready),
    .io_stream_in_166_valid(merger_io_stream_in_166_valid),
    .io_stream_in_166_bits(merger_io_stream_in_166_bits),
    .io_stream_in_167_ready(merger_io_stream_in_167_ready),
    .io_stream_in_167_valid(merger_io_stream_in_167_valid),
    .io_stream_in_167_bits(merger_io_stream_in_167_bits),
    .io_stream_in_168_ready(merger_io_stream_in_168_ready),
    .io_stream_in_168_valid(merger_io_stream_in_168_valid),
    .io_stream_in_168_bits(merger_io_stream_in_168_bits),
    .io_stream_in_169_ready(merger_io_stream_in_169_ready),
    .io_stream_in_169_valid(merger_io_stream_in_169_valid),
    .io_stream_in_169_bits(merger_io_stream_in_169_bits),
    .io_stream_in_170_ready(merger_io_stream_in_170_ready),
    .io_stream_in_170_valid(merger_io_stream_in_170_valid),
    .io_stream_in_170_bits(merger_io_stream_in_170_bits),
    .io_stream_in_171_ready(merger_io_stream_in_171_ready),
    .io_stream_in_171_valid(merger_io_stream_in_171_valid),
    .io_stream_in_171_bits(merger_io_stream_in_171_bits),
    .io_stream_in_172_ready(merger_io_stream_in_172_ready),
    .io_stream_in_172_valid(merger_io_stream_in_172_valid),
    .io_stream_in_172_bits(merger_io_stream_in_172_bits),
    .io_stream_in_173_ready(merger_io_stream_in_173_ready),
    .io_stream_in_173_valid(merger_io_stream_in_173_valid),
    .io_stream_in_173_bits(merger_io_stream_in_173_bits),
    .io_stream_in_174_ready(merger_io_stream_in_174_ready),
    .io_stream_in_174_valid(merger_io_stream_in_174_valid),
    .io_stream_in_174_bits(merger_io_stream_in_174_bits),
    .io_stream_in_175_ready(merger_io_stream_in_175_ready),
    .io_stream_in_175_valid(merger_io_stream_in_175_valid),
    .io_stream_in_175_bits(merger_io_stream_in_175_bits),
    .io_stream_in_176_ready(merger_io_stream_in_176_ready),
    .io_stream_in_176_valid(merger_io_stream_in_176_valid),
    .io_stream_in_176_bits(merger_io_stream_in_176_bits),
    .io_stream_in_177_ready(merger_io_stream_in_177_ready),
    .io_stream_in_177_valid(merger_io_stream_in_177_valid),
    .io_stream_in_177_bits(merger_io_stream_in_177_bits),
    .io_stream_in_178_ready(merger_io_stream_in_178_ready),
    .io_stream_in_178_valid(merger_io_stream_in_178_valid),
    .io_stream_in_178_bits(merger_io_stream_in_178_bits),
    .io_stream_in_179_ready(merger_io_stream_in_179_ready),
    .io_stream_in_179_valid(merger_io_stream_in_179_valid),
    .io_stream_in_179_bits(merger_io_stream_in_179_bits),
    .io_stream_in_180_ready(merger_io_stream_in_180_ready),
    .io_stream_in_180_valid(merger_io_stream_in_180_valid),
    .io_stream_in_180_bits(merger_io_stream_in_180_bits),
    .io_stream_in_181_ready(merger_io_stream_in_181_ready),
    .io_stream_in_181_valid(merger_io_stream_in_181_valid),
    .io_stream_in_181_bits(merger_io_stream_in_181_bits),
    .io_stream_in_182_ready(merger_io_stream_in_182_ready),
    .io_stream_in_182_valid(merger_io_stream_in_182_valid),
    .io_stream_in_182_bits(merger_io_stream_in_182_bits),
    .io_stream_in_183_ready(merger_io_stream_in_183_ready),
    .io_stream_in_183_valid(merger_io_stream_in_183_valid),
    .io_stream_in_183_bits(merger_io_stream_in_183_bits),
    .io_stream_in_184_ready(merger_io_stream_in_184_ready),
    .io_stream_in_184_valid(merger_io_stream_in_184_valid),
    .io_stream_in_184_bits(merger_io_stream_in_184_bits),
    .io_stream_in_185_ready(merger_io_stream_in_185_ready),
    .io_stream_in_185_valid(merger_io_stream_in_185_valid),
    .io_stream_in_185_bits(merger_io_stream_in_185_bits),
    .io_stream_in_186_ready(merger_io_stream_in_186_ready),
    .io_stream_in_186_valid(merger_io_stream_in_186_valid),
    .io_stream_in_186_bits(merger_io_stream_in_186_bits),
    .io_stream_in_187_ready(merger_io_stream_in_187_ready),
    .io_stream_in_187_valid(merger_io_stream_in_187_valid),
    .io_stream_in_187_bits(merger_io_stream_in_187_bits),
    .io_stream_in_188_ready(merger_io_stream_in_188_ready),
    .io_stream_in_188_valid(merger_io_stream_in_188_valid),
    .io_stream_in_188_bits(merger_io_stream_in_188_bits),
    .io_stream_in_189_ready(merger_io_stream_in_189_ready),
    .io_stream_in_189_valid(merger_io_stream_in_189_valid),
    .io_stream_in_189_bits(merger_io_stream_in_189_bits),
    .io_stream_in_190_ready(merger_io_stream_in_190_ready),
    .io_stream_in_190_valid(merger_io_stream_in_190_valid),
    .io_stream_in_190_bits(merger_io_stream_in_190_bits),
    .io_stream_in_191_ready(merger_io_stream_in_191_ready),
    .io_stream_in_191_valid(merger_io_stream_in_191_valid),
    .io_stream_in_191_bits(merger_io_stream_in_191_bits),
    .io_stream_in_192_ready(merger_io_stream_in_192_ready),
    .io_stream_in_192_valid(merger_io_stream_in_192_valid),
    .io_stream_in_192_bits(merger_io_stream_in_192_bits),
    .io_stream_in_193_ready(merger_io_stream_in_193_ready),
    .io_stream_in_193_valid(merger_io_stream_in_193_valid),
    .io_stream_in_193_bits(merger_io_stream_in_193_bits),
    .io_stream_in_194_ready(merger_io_stream_in_194_ready),
    .io_stream_in_194_valid(merger_io_stream_in_194_valid),
    .io_stream_in_194_bits(merger_io_stream_in_194_bits),
    .io_stream_in_195_ready(merger_io_stream_in_195_ready),
    .io_stream_in_195_valid(merger_io_stream_in_195_valid),
    .io_stream_in_195_bits(merger_io_stream_in_195_bits),
    .io_stream_in_196_ready(merger_io_stream_in_196_ready),
    .io_stream_in_196_valid(merger_io_stream_in_196_valid),
    .io_stream_in_196_bits(merger_io_stream_in_196_bits),
    .io_stream_in_197_ready(merger_io_stream_in_197_ready),
    .io_stream_in_197_valid(merger_io_stream_in_197_valid),
    .io_stream_in_197_bits(merger_io_stream_in_197_bits),
    .io_stream_in_198_ready(merger_io_stream_in_198_ready),
    .io_stream_in_198_valid(merger_io_stream_in_198_valid),
    .io_stream_in_198_bits(merger_io_stream_in_198_bits),
    .io_stream_in_199_ready(merger_io_stream_in_199_ready),
    .io_stream_in_199_valid(merger_io_stream_in_199_valid),
    .io_stream_in_199_bits(merger_io_stream_in_199_bits),
    .io_stream_in_200_ready(merger_io_stream_in_200_ready),
    .io_stream_in_200_valid(merger_io_stream_in_200_valid),
    .io_stream_in_200_bits(merger_io_stream_in_200_bits),
    .io_stream_in_201_ready(merger_io_stream_in_201_ready),
    .io_stream_in_201_valid(merger_io_stream_in_201_valid),
    .io_stream_in_201_bits(merger_io_stream_in_201_bits),
    .io_stream_in_202_ready(merger_io_stream_in_202_ready),
    .io_stream_in_202_valid(merger_io_stream_in_202_valid),
    .io_stream_in_202_bits(merger_io_stream_in_202_bits),
    .io_stream_in_203_ready(merger_io_stream_in_203_ready),
    .io_stream_in_203_valid(merger_io_stream_in_203_valid),
    .io_stream_in_203_bits(merger_io_stream_in_203_bits),
    .io_stream_in_204_ready(merger_io_stream_in_204_ready),
    .io_stream_in_204_valid(merger_io_stream_in_204_valid),
    .io_stream_in_204_bits(merger_io_stream_in_204_bits),
    .io_stream_in_205_ready(merger_io_stream_in_205_ready),
    .io_stream_in_205_valid(merger_io_stream_in_205_valid),
    .io_stream_in_205_bits(merger_io_stream_in_205_bits),
    .io_stream_in_206_ready(merger_io_stream_in_206_ready),
    .io_stream_in_206_valid(merger_io_stream_in_206_valid),
    .io_stream_in_206_bits(merger_io_stream_in_206_bits),
    .io_stream_in_207_ready(merger_io_stream_in_207_ready),
    .io_stream_in_207_valid(merger_io_stream_in_207_valid),
    .io_stream_in_207_bits(merger_io_stream_in_207_bits),
    .io_stream_in_208_ready(merger_io_stream_in_208_ready),
    .io_stream_in_208_valid(merger_io_stream_in_208_valid),
    .io_stream_in_208_bits(merger_io_stream_in_208_bits),
    .io_stream_in_209_ready(merger_io_stream_in_209_ready),
    .io_stream_in_209_valid(merger_io_stream_in_209_valid),
    .io_stream_in_209_bits(merger_io_stream_in_209_bits),
    .io_stream_in_210_ready(merger_io_stream_in_210_ready),
    .io_stream_in_210_valid(merger_io_stream_in_210_valid),
    .io_stream_in_210_bits(merger_io_stream_in_210_bits),
    .io_stream_in_211_ready(merger_io_stream_in_211_ready),
    .io_stream_in_211_valid(merger_io_stream_in_211_valid),
    .io_stream_in_211_bits(merger_io_stream_in_211_bits),
    .io_stream_in_212_ready(merger_io_stream_in_212_ready),
    .io_stream_in_212_valid(merger_io_stream_in_212_valid),
    .io_stream_in_212_bits(merger_io_stream_in_212_bits),
    .io_stream_in_213_ready(merger_io_stream_in_213_ready),
    .io_stream_in_213_valid(merger_io_stream_in_213_valid),
    .io_stream_in_213_bits(merger_io_stream_in_213_bits),
    .io_stream_in_214_ready(merger_io_stream_in_214_ready),
    .io_stream_in_214_valid(merger_io_stream_in_214_valid),
    .io_stream_in_214_bits(merger_io_stream_in_214_bits),
    .io_stream_in_215_ready(merger_io_stream_in_215_ready),
    .io_stream_in_215_valid(merger_io_stream_in_215_valid),
    .io_stream_in_215_bits(merger_io_stream_in_215_bits),
    .io_stream_in_216_ready(merger_io_stream_in_216_ready),
    .io_stream_in_216_valid(merger_io_stream_in_216_valid),
    .io_stream_in_216_bits(merger_io_stream_in_216_bits),
    .io_stream_in_217_ready(merger_io_stream_in_217_ready),
    .io_stream_in_217_valid(merger_io_stream_in_217_valid),
    .io_stream_in_217_bits(merger_io_stream_in_217_bits),
    .io_stream_in_218_ready(merger_io_stream_in_218_ready),
    .io_stream_in_218_valid(merger_io_stream_in_218_valid),
    .io_stream_in_218_bits(merger_io_stream_in_218_bits),
    .io_stream_in_219_ready(merger_io_stream_in_219_ready),
    .io_stream_in_219_valid(merger_io_stream_in_219_valid),
    .io_stream_in_219_bits(merger_io_stream_in_219_bits),
    .io_stream_in_220_ready(merger_io_stream_in_220_ready),
    .io_stream_in_220_valid(merger_io_stream_in_220_valid),
    .io_stream_in_220_bits(merger_io_stream_in_220_bits),
    .io_stream_in_221_ready(merger_io_stream_in_221_ready),
    .io_stream_in_221_valid(merger_io_stream_in_221_valid),
    .io_stream_in_221_bits(merger_io_stream_in_221_bits),
    .io_stream_in_222_ready(merger_io_stream_in_222_ready),
    .io_stream_in_222_valid(merger_io_stream_in_222_valid),
    .io_stream_in_222_bits(merger_io_stream_in_222_bits),
    .io_stream_in_223_ready(merger_io_stream_in_223_ready),
    .io_stream_in_223_valid(merger_io_stream_in_223_valid),
    .io_stream_in_223_bits(merger_io_stream_in_223_bits),
    .io_stream_in_224_ready(merger_io_stream_in_224_ready),
    .io_stream_in_224_valid(merger_io_stream_in_224_valid),
    .io_stream_in_224_bits(merger_io_stream_in_224_bits),
    .io_stream_in_225_ready(merger_io_stream_in_225_ready),
    .io_stream_in_225_valid(merger_io_stream_in_225_valid),
    .io_stream_in_225_bits(merger_io_stream_in_225_bits),
    .io_stream_in_226_ready(merger_io_stream_in_226_ready),
    .io_stream_in_226_valid(merger_io_stream_in_226_valid),
    .io_stream_in_226_bits(merger_io_stream_in_226_bits),
    .io_stream_in_227_ready(merger_io_stream_in_227_ready),
    .io_stream_in_227_valid(merger_io_stream_in_227_valid),
    .io_stream_in_227_bits(merger_io_stream_in_227_bits),
    .io_stream_in_228_ready(merger_io_stream_in_228_ready),
    .io_stream_in_228_valid(merger_io_stream_in_228_valid),
    .io_stream_in_228_bits(merger_io_stream_in_228_bits),
    .io_stream_in_229_ready(merger_io_stream_in_229_ready),
    .io_stream_in_229_valid(merger_io_stream_in_229_valid),
    .io_stream_in_229_bits(merger_io_stream_in_229_bits),
    .io_stream_in_230_ready(merger_io_stream_in_230_ready),
    .io_stream_in_230_valid(merger_io_stream_in_230_valid),
    .io_stream_in_230_bits(merger_io_stream_in_230_bits),
    .io_stream_in_231_ready(merger_io_stream_in_231_ready),
    .io_stream_in_231_valid(merger_io_stream_in_231_valid),
    .io_stream_in_231_bits(merger_io_stream_in_231_bits),
    .io_stream_in_232_ready(merger_io_stream_in_232_ready),
    .io_stream_in_232_valid(merger_io_stream_in_232_valid),
    .io_stream_in_232_bits(merger_io_stream_in_232_bits),
    .io_stream_in_233_ready(merger_io_stream_in_233_ready),
    .io_stream_in_233_valid(merger_io_stream_in_233_valid),
    .io_stream_in_233_bits(merger_io_stream_in_233_bits),
    .io_stream_in_234_ready(merger_io_stream_in_234_ready),
    .io_stream_in_234_valid(merger_io_stream_in_234_valid),
    .io_stream_in_234_bits(merger_io_stream_in_234_bits),
    .io_stream_in_235_ready(merger_io_stream_in_235_ready),
    .io_stream_in_235_valid(merger_io_stream_in_235_valid),
    .io_stream_in_235_bits(merger_io_stream_in_235_bits),
    .io_stream_in_236_ready(merger_io_stream_in_236_ready),
    .io_stream_in_236_valid(merger_io_stream_in_236_valid),
    .io_stream_in_236_bits(merger_io_stream_in_236_bits),
    .io_stream_in_237_ready(merger_io_stream_in_237_ready),
    .io_stream_in_237_valid(merger_io_stream_in_237_valid),
    .io_stream_in_237_bits(merger_io_stream_in_237_bits),
    .io_stream_in_238_ready(merger_io_stream_in_238_ready),
    .io_stream_in_238_valid(merger_io_stream_in_238_valid),
    .io_stream_in_238_bits(merger_io_stream_in_238_bits),
    .io_stream_in_239_ready(merger_io_stream_in_239_ready),
    .io_stream_in_239_valid(merger_io_stream_in_239_valid),
    .io_stream_in_239_bits(merger_io_stream_in_239_bits),
    .io_stream_in_240_ready(merger_io_stream_in_240_ready),
    .io_stream_in_240_valid(merger_io_stream_in_240_valid),
    .io_stream_in_240_bits(merger_io_stream_in_240_bits),
    .io_stream_in_241_ready(merger_io_stream_in_241_ready),
    .io_stream_in_241_valid(merger_io_stream_in_241_valid),
    .io_stream_in_241_bits(merger_io_stream_in_241_bits),
    .io_stream_in_242_ready(merger_io_stream_in_242_ready),
    .io_stream_in_242_valid(merger_io_stream_in_242_valid),
    .io_stream_in_242_bits(merger_io_stream_in_242_bits),
    .io_stream_in_243_ready(merger_io_stream_in_243_ready),
    .io_stream_in_243_valid(merger_io_stream_in_243_valid),
    .io_stream_in_243_bits(merger_io_stream_in_243_bits),
    .io_stream_in_244_ready(merger_io_stream_in_244_ready),
    .io_stream_in_244_valid(merger_io_stream_in_244_valid),
    .io_stream_in_244_bits(merger_io_stream_in_244_bits),
    .io_stream_in_245_ready(merger_io_stream_in_245_ready),
    .io_stream_in_245_valid(merger_io_stream_in_245_valid),
    .io_stream_in_245_bits(merger_io_stream_in_245_bits),
    .io_stream_in_246_ready(merger_io_stream_in_246_ready),
    .io_stream_in_246_valid(merger_io_stream_in_246_valid),
    .io_stream_in_246_bits(merger_io_stream_in_246_bits),
    .io_stream_in_247_ready(merger_io_stream_in_247_ready),
    .io_stream_in_247_valid(merger_io_stream_in_247_valid),
    .io_stream_in_247_bits(merger_io_stream_in_247_bits),
    .io_stream_in_248_ready(merger_io_stream_in_248_ready),
    .io_stream_in_248_valid(merger_io_stream_in_248_valid),
    .io_stream_in_248_bits(merger_io_stream_in_248_bits),
    .io_stream_in_249_ready(merger_io_stream_in_249_ready),
    .io_stream_in_249_valid(merger_io_stream_in_249_valid),
    .io_stream_in_249_bits(merger_io_stream_in_249_bits),
    .io_stream_in_250_ready(merger_io_stream_in_250_ready),
    .io_stream_in_250_valid(merger_io_stream_in_250_valid),
    .io_stream_in_250_bits(merger_io_stream_in_250_bits),
    .io_stream_in_251_ready(merger_io_stream_in_251_ready),
    .io_stream_in_251_valid(merger_io_stream_in_251_valid),
    .io_stream_in_251_bits(merger_io_stream_in_251_bits),
    .io_stream_in_252_ready(merger_io_stream_in_252_ready),
    .io_stream_in_252_valid(merger_io_stream_in_252_valid),
    .io_stream_in_252_bits(merger_io_stream_in_252_bits),
    .io_stream_in_253_ready(merger_io_stream_in_253_ready),
    .io_stream_in_253_valid(merger_io_stream_in_253_valid),
    .io_stream_in_253_bits(merger_io_stream_in_253_bits),
    .io_stream_in_254_ready(merger_io_stream_in_254_ready),
    .io_stream_in_254_valid(merger_io_stream_in_254_valid),
    .io_stream_in_254_bits(merger_io_stream_in_254_bits),
    .io_stream_in_255_ready(merger_io_stream_in_255_ready),
    .io_stream_in_255_valid(merger_io_stream_in_255_valid),
    .io_stream_in_255_bits(merger_io_stream_in_255_bits),
    .io_stream_out_ready(merger_io_stream_out_ready),
    .io_stream_out_valid(merger_io_stream_out_valid),
    .io_stream_out_bits(merger_io_stream_out_bits)
  );
  assign io_stream_in_0_ready = merger_io_stream_in_0_ready; // @[Stab.scala 292:64]
  assign io_stream_in_1_ready = merger_io_stream_in_1_ready; // @[Stab.scala 292:64]
  assign io_stream_in_2_ready = merger_io_stream_in_2_ready; // @[Stab.scala 292:64]
  assign io_stream_in_3_ready = merger_io_stream_in_3_ready; // @[Stab.scala 292:64]
  assign io_stream_in_4_ready = merger_io_stream_in_4_ready; // @[Stab.scala 292:64]
  assign io_stream_in_5_ready = merger_io_stream_in_5_ready; // @[Stab.scala 292:64]
  assign io_stream_in_6_ready = merger_io_stream_in_6_ready; // @[Stab.scala 292:64]
  assign io_stream_in_7_ready = merger_io_stream_in_7_ready; // @[Stab.scala 292:64]
  assign io_stream_in_8_ready = merger_io_stream_in_8_ready; // @[Stab.scala 292:64]
  assign io_stream_in_9_ready = merger_io_stream_in_9_ready; // @[Stab.scala 292:64]
  assign io_stream_in_10_ready = merger_io_stream_in_10_ready; // @[Stab.scala 292:64]
  assign io_stream_in_11_ready = merger_io_stream_in_11_ready; // @[Stab.scala 292:64]
  assign io_stream_in_12_ready = merger_io_stream_in_12_ready; // @[Stab.scala 292:64]
  assign io_stream_in_13_ready = merger_io_stream_in_13_ready; // @[Stab.scala 292:64]
  assign io_stream_in_14_ready = merger_io_stream_in_14_ready; // @[Stab.scala 292:64]
  assign io_stream_in_15_ready = merger_io_stream_in_15_ready; // @[Stab.scala 292:64]
  assign io_stream_in_16_ready = merger_io_stream_in_16_ready; // @[Stab.scala 292:64]
  assign io_stream_in_17_ready = merger_io_stream_in_17_ready; // @[Stab.scala 292:64]
  assign io_stream_in_18_ready = merger_io_stream_in_18_ready; // @[Stab.scala 292:64]
  assign io_stream_in_19_ready = merger_io_stream_in_19_ready; // @[Stab.scala 292:64]
  assign io_stream_in_20_ready = merger_io_stream_in_20_ready; // @[Stab.scala 292:64]
  assign io_stream_in_21_ready = merger_io_stream_in_21_ready; // @[Stab.scala 292:64]
  assign io_stream_in_22_ready = merger_io_stream_in_22_ready; // @[Stab.scala 292:64]
  assign io_stream_in_23_ready = merger_io_stream_in_23_ready; // @[Stab.scala 292:64]
  assign io_stream_in_24_ready = merger_io_stream_in_24_ready; // @[Stab.scala 292:64]
  assign io_stream_in_25_ready = merger_io_stream_in_25_ready; // @[Stab.scala 292:64]
  assign io_stream_in_26_ready = merger_io_stream_in_26_ready; // @[Stab.scala 292:64]
  assign io_stream_in_27_ready = merger_io_stream_in_27_ready; // @[Stab.scala 292:64]
  assign io_stream_in_28_ready = merger_io_stream_in_28_ready; // @[Stab.scala 292:64]
  assign io_stream_in_29_ready = merger_io_stream_in_29_ready; // @[Stab.scala 292:64]
  assign io_stream_in_30_ready = merger_io_stream_in_30_ready; // @[Stab.scala 292:64]
  assign io_stream_in_31_ready = merger_io_stream_in_31_ready; // @[Stab.scala 292:64]
  assign io_stream_in_32_ready = merger_io_stream_in_32_ready; // @[Stab.scala 292:64]
  assign io_stream_in_33_ready = merger_io_stream_in_33_ready; // @[Stab.scala 292:64]
  assign io_stream_in_34_ready = merger_io_stream_in_34_ready; // @[Stab.scala 292:64]
  assign io_stream_in_35_ready = merger_io_stream_in_35_ready; // @[Stab.scala 292:64]
  assign io_stream_in_36_ready = merger_io_stream_in_36_ready; // @[Stab.scala 292:64]
  assign io_stream_in_37_ready = merger_io_stream_in_37_ready; // @[Stab.scala 292:64]
  assign io_stream_in_38_ready = merger_io_stream_in_38_ready; // @[Stab.scala 292:64]
  assign io_stream_in_39_ready = merger_io_stream_in_39_ready; // @[Stab.scala 292:64]
  assign io_stream_in_40_ready = merger_io_stream_in_40_ready; // @[Stab.scala 292:64]
  assign io_stream_in_41_ready = merger_io_stream_in_41_ready; // @[Stab.scala 292:64]
  assign io_stream_in_42_ready = merger_io_stream_in_42_ready; // @[Stab.scala 292:64]
  assign io_stream_in_43_ready = merger_io_stream_in_43_ready; // @[Stab.scala 292:64]
  assign io_stream_in_44_ready = merger_io_stream_in_44_ready; // @[Stab.scala 292:64]
  assign io_stream_in_45_ready = merger_io_stream_in_45_ready; // @[Stab.scala 292:64]
  assign io_stream_in_46_ready = merger_io_stream_in_46_ready; // @[Stab.scala 292:64]
  assign io_stream_in_47_ready = merger_io_stream_in_47_ready; // @[Stab.scala 292:64]
  assign io_stream_in_48_ready = merger_io_stream_in_48_ready; // @[Stab.scala 292:64]
  assign io_stream_in_49_ready = merger_io_stream_in_49_ready; // @[Stab.scala 292:64]
  assign io_stream_in_50_ready = merger_io_stream_in_50_ready; // @[Stab.scala 292:64]
  assign io_stream_in_51_ready = merger_io_stream_in_51_ready; // @[Stab.scala 292:64]
  assign io_stream_in_52_ready = merger_io_stream_in_52_ready; // @[Stab.scala 292:64]
  assign io_stream_in_53_ready = merger_io_stream_in_53_ready; // @[Stab.scala 292:64]
  assign io_stream_in_54_ready = merger_io_stream_in_54_ready; // @[Stab.scala 292:64]
  assign io_stream_in_55_ready = merger_io_stream_in_55_ready; // @[Stab.scala 292:64]
  assign io_stream_in_56_ready = merger_io_stream_in_56_ready; // @[Stab.scala 292:64]
  assign io_stream_in_57_ready = merger_io_stream_in_57_ready; // @[Stab.scala 292:64]
  assign io_stream_in_58_ready = merger_io_stream_in_58_ready; // @[Stab.scala 292:64]
  assign io_stream_in_59_ready = merger_io_stream_in_59_ready; // @[Stab.scala 292:64]
  assign io_stream_in_60_ready = merger_io_stream_in_60_ready; // @[Stab.scala 292:64]
  assign io_stream_in_61_ready = merger_io_stream_in_61_ready; // @[Stab.scala 292:64]
  assign io_stream_in_62_ready = merger_io_stream_in_62_ready; // @[Stab.scala 292:64]
  assign io_stream_in_63_ready = merger_io_stream_in_63_ready; // @[Stab.scala 292:64]
  assign io_stream_in_64_ready = merger_io_stream_in_64_ready; // @[Stab.scala 292:64]
  assign io_stream_in_65_ready = merger_io_stream_in_65_ready; // @[Stab.scala 292:64]
  assign io_stream_in_66_ready = merger_io_stream_in_66_ready; // @[Stab.scala 292:64]
  assign io_stream_in_67_ready = merger_io_stream_in_67_ready; // @[Stab.scala 292:64]
  assign io_stream_in_68_ready = merger_io_stream_in_68_ready; // @[Stab.scala 292:64]
  assign io_stream_in_69_ready = merger_io_stream_in_69_ready; // @[Stab.scala 292:64]
  assign io_stream_in_70_ready = merger_io_stream_in_70_ready; // @[Stab.scala 292:64]
  assign io_stream_in_71_ready = merger_io_stream_in_71_ready; // @[Stab.scala 292:64]
  assign io_stream_in_72_ready = merger_io_stream_in_72_ready; // @[Stab.scala 292:64]
  assign io_stream_in_73_ready = merger_io_stream_in_73_ready; // @[Stab.scala 292:64]
  assign io_stream_in_74_ready = merger_io_stream_in_74_ready; // @[Stab.scala 292:64]
  assign io_stream_in_75_ready = merger_io_stream_in_75_ready; // @[Stab.scala 292:64]
  assign io_stream_in_76_ready = merger_io_stream_in_76_ready; // @[Stab.scala 292:64]
  assign io_stream_in_77_ready = merger_io_stream_in_77_ready; // @[Stab.scala 292:64]
  assign io_stream_in_78_ready = merger_io_stream_in_78_ready; // @[Stab.scala 292:64]
  assign io_stream_in_79_ready = merger_io_stream_in_79_ready; // @[Stab.scala 292:64]
  assign io_stream_in_80_ready = merger_io_stream_in_80_ready; // @[Stab.scala 292:64]
  assign io_stream_in_81_ready = merger_io_stream_in_81_ready; // @[Stab.scala 292:64]
  assign io_stream_in_82_ready = merger_io_stream_in_82_ready; // @[Stab.scala 292:64]
  assign io_stream_in_83_ready = merger_io_stream_in_83_ready; // @[Stab.scala 292:64]
  assign io_stream_in_84_ready = merger_io_stream_in_84_ready; // @[Stab.scala 292:64]
  assign io_stream_in_85_ready = merger_io_stream_in_85_ready; // @[Stab.scala 292:64]
  assign io_stream_in_86_ready = merger_io_stream_in_86_ready; // @[Stab.scala 292:64]
  assign io_stream_in_87_ready = merger_io_stream_in_87_ready; // @[Stab.scala 292:64]
  assign io_stream_in_88_ready = merger_io_stream_in_88_ready; // @[Stab.scala 292:64]
  assign io_stream_in_89_ready = merger_io_stream_in_89_ready; // @[Stab.scala 292:64]
  assign io_stream_in_90_ready = merger_io_stream_in_90_ready; // @[Stab.scala 292:64]
  assign io_stream_in_91_ready = merger_io_stream_in_91_ready; // @[Stab.scala 292:64]
  assign io_stream_in_92_ready = merger_io_stream_in_92_ready; // @[Stab.scala 292:64]
  assign io_stream_in_93_ready = merger_io_stream_in_93_ready; // @[Stab.scala 292:64]
  assign io_stream_in_94_ready = merger_io_stream_in_94_ready; // @[Stab.scala 292:64]
  assign io_stream_in_95_ready = merger_io_stream_in_95_ready; // @[Stab.scala 292:64]
  assign io_stream_in_96_ready = merger_io_stream_in_96_ready; // @[Stab.scala 292:64]
  assign io_stream_in_97_ready = merger_io_stream_in_97_ready; // @[Stab.scala 292:64]
  assign io_stream_in_98_ready = merger_io_stream_in_98_ready; // @[Stab.scala 292:64]
  assign io_stream_in_99_ready = merger_io_stream_in_99_ready; // @[Stab.scala 292:64]
  assign io_stream_in_100_ready = merger_io_stream_in_100_ready; // @[Stab.scala 292:64]
  assign io_stream_in_101_ready = merger_io_stream_in_101_ready; // @[Stab.scala 292:64]
  assign io_stream_in_102_ready = merger_io_stream_in_102_ready; // @[Stab.scala 292:64]
  assign io_stream_in_103_ready = merger_io_stream_in_103_ready; // @[Stab.scala 292:64]
  assign io_stream_in_104_ready = merger_io_stream_in_104_ready; // @[Stab.scala 292:64]
  assign io_stream_in_105_ready = merger_io_stream_in_105_ready; // @[Stab.scala 292:64]
  assign io_stream_in_106_ready = merger_io_stream_in_106_ready; // @[Stab.scala 292:64]
  assign io_stream_in_107_ready = merger_io_stream_in_107_ready; // @[Stab.scala 292:64]
  assign io_stream_in_108_ready = merger_io_stream_in_108_ready; // @[Stab.scala 292:64]
  assign io_stream_in_109_ready = merger_io_stream_in_109_ready; // @[Stab.scala 292:64]
  assign io_stream_in_110_ready = merger_io_stream_in_110_ready; // @[Stab.scala 292:64]
  assign io_stream_in_111_ready = merger_io_stream_in_111_ready; // @[Stab.scala 292:64]
  assign io_stream_in_112_ready = merger_io_stream_in_112_ready; // @[Stab.scala 292:64]
  assign io_stream_in_113_ready = merger_io_stream_in_113_ready; // @[Stab.scala 292:64]
  assign io_stream_in_114_ready = merger_io_stream_in_114_ready; // @[Stab.scala 292:64]
  assign io_stream_in_115_ready = merger_io_stream_in_115_ready; // @[Stab.scala 292:64]
  assign io_stream_in_116_ready = merger_io_stream_in_116_ready; // @[Stab.scala 292:64]
  assign io_stream_in_117_ready = merger_io_stream_in_117_ready; // @[Stab.scala 292:64]
  assign io_stream_in_118_ready = merger_io_stream_in_118_ready; // @[Stab.scala 292:64]
  assign io_stream_in_119_ready = merger_io_stream_in_119_ready; // @[Stab.scala 292:64]
  assign io_stream_in_120_ready = merger_io_stream_in_120_ready; // @[Stab.scala 292:64]
  assign io_stream_in_121_ready = merger_io_stream_in_121_ready; // @[Stab.scala 292:64]
  assign io_stream_in_122_ready = merger_io_stream_in_122_ready; // @[Stab.scala 292:64]
  assign io_stream_in_123_ready = merger_io_stream_in_123_ready; // @[Stab.scala 292:64]
  assign io_stream_in_124_ready = merger_io_stream_in_124_ready; // @[Stab.scala 292:64]
  assign io_stream_in_125_ready = merger_io_stream_in_125_ready; // @[Stab.scala 292:64]
  assign io_stream_in_126_ready = merger_io_stream_in_126_ready; // @[Stab.scala 292:64]
  assign io_stream_in_127_ready = merger_io_stream_in_127_ready; // @[Stab.scala 292:64]
  assign io_stream_in_128_ready = merger_io_stream_in_128_ready; // @[Stab.scala 292:64]
  assign io_stream_in_129_ready = merger_io_stream_in_129_ready; // @[Stab.scala 292:64]
  assign io_stream_in_130_ready = merger_io_stream_in_130_ready; // @[Stab.scala 292:64]
  assign io_stream_in_131_ready = merger_io_stream_in_131_ready; // @[Stab.scala 292:64]
  assign io_stream_in_132_ready = merger_io_stream_in_132_ready; // @[Stab.scala 292:64]
  assign io_stream_in_133_ready = merger_io_stream_in_133_ready; // @[Stab.scala 292:64]
  assign io_stream_in_134_ready = merger_io_stream_in_134_ready; // @[Stab.scala 292:64]
  assign io_stream_in_135_ready = merger_io_stream_in_135_ready; // @[Stab.scala 292:64]
  assign io_stream_in_136_ready = merger_io_stream_in_136_ready; // @[Stab.scala 292:64]
  assign io_stream_in_137_ready = merger_io_stream_in_137_ready; // @[Stab.scala 292:64]
  assign io_stream_in_138_ready = merger_io_stream_in_138_ready; // @[Stab.scala 292:64]
  assign io_stream_in_139_ready = merger_io_stream_in_139_ready; // @[Stab.scala 292:64]
  assign io_stream_in_140_ready = merger_io_stream_in_140_ready; // @[Stab.scala 292:64]
  assign io_stream_in_141_ready = merger_io_stream_in_141_ready; // @[Stab.scala 292:64]
  assign io_stream_in_142_ready = merger_io_stream_in_142_ready; // @[Stab.scala 292:64]
  assign io_stream_in_143_ready = merger_io_stream_in_143_ready; // @[Stab.scala 292:64]
  assign io_stream_in_144_ready = merger_io_stream_in_144_ready; // @[Stab.scala 292:64]
  assign io_stream_in_145_ready = merger_io_stream_in_145_ready; // @[Stab.scala 292:64]
  assign io_stream_in_146_ready = merger_io_stream_in_146_ready; // @[Stab.scala 292:64]
  assign io_stream_in_147_ready = merger_io_stream_in_147_ready; // @[Stab.scala 292:64]
  assign io_stream_in_148_ready = merger_io_stream_in_148_ready; // @[Stab.scala 292:64]
  assign io_stream_in_149_ready = merger_io_stream_in_149_ready; // @[Stab.scala 292:64]
  assign io_stream_in_150_ready = merger_io_stream_in_150_ready; // @[Stab.scala 292:64]
  assign io_stream_in_151_ready = merger_io_stream_in_151_ready; // @[Stab.scala 292:64]
  assign io_stream_in_152_ready = merger_io_stream_in_152_ready; // @[Stab.scala 292:64]
  assign io_stream_in_153_ready = merger_io_stream_in_153_ready; // @[Stab.scala 292:64]
  assign io_stream_in_154_ready = merger_io_stream_in_154_ready; // @[Stab.scala 292:64]
  assign io_stream_in_155_ready = merger_io_stream_in_155_ready; // @[Stab.scala 292:64]
  assign io_stream_in_156_ready = merger_io_stream_in_156_ready; // @[Stab.scala 292:64]
  assign io_stream_in_157_ready = merger_io_stream_in_157_ready; // @[Stab.scala 292:64]
  assign io_stream_in_158_ready = merger_io_stream_in_158_ready; // @[Stab.scala 292:64]
  assign io_stream_in_159_ready = merger_io_stream_in_159_ready; // @[Stab.scala 292:64]
  assign io_stream_in_160_ready = merger_io_stream_in_160_ready; // @[Stab.scala 292:64]
  assign io_stream_in_161_ready = merger_io_stream_in_161_ready; // @[Stab.scala 292:64]
  assign io_stream_in_162_ready = merger_io_stream_in_162_ready; // @[Stab.scala 292:64]
  assign io_stream_in_163_ready = merger_io_stream_in_163_ready; // @[Stab.scala 292:64]
  assign io_stream_in_164_ready = merger_io_stream_in_164_ready; // @[Stab.scala 292:64]
  assign io_stream_in_165_ready = merger_io_stream_in_165_ready; // @[Stab.scala 292:64]
  assign io_stream_in_166_ready = merger_io_stream_in_166_ready; // @[Stab.scala 292:64]
  assign io_stream_in_167_ready = merger_io_stream_in_167_ready; // @[Stab.scala 292:64]
  assign io_stream_in_168_ready = merger_io_stream_in_168_ready; // @[Stab.scala 292:64]
  assign io_stream_in_169_ready = merger_io_stream_in_169_ready; // @[Stab.scala 292:64]
  assign io_stream_in_170_ready = merger_io_stream_in_170_ready; // @[Stab.scala 292:64]
  assign io_stream_in_171_ready = merger_io_stream_in_171_ready; // @[Stab.scala 292:64]
  assign io_stream_in_172_ready = merger_io_stream_in_172_ready; // @[Stab.scala 292:64]
  assign io_stream_in_173_ready = merger_io_stream_in_173_ready; // @[Stab.scala 292:64]
  assign io_stream_in_174_ready = merger_io_stream_in_174_ready; // @[Stab.scala 292:64]
  assign io_stream_in_175_ready = merger_io_stream_in_175_ready; // @[Stab.scala 292:64]
  assign io_stream_in_176_ready = merger_io_stream_in_176_ready; // @[Stab.scala 292:64]
  assign io_stream_in_177_ready = merger_io_stream_in_177_ready; // @[Stab.scala 292:64]
  assign io_stream_in_178_ready = merger_io_stream_in_178_ready; // @[Stab.scala 292:64]
  assign io_stream_in_179_ready = merger_io_stream_in_179_ready; // @[Stab.scala 292:64]
  assign io_stream_in_180_ready = merger_io_stream_in_180_ready; // @[Stab.scala 292:64]
  assign io_stream_in_181_ready = merger_io_stream_in_181_ready; // @[Stab.scala 292:64]
  assign io_stream_in_182_ready = merger_io_stream_in_182_ready; // @[Stab.scala 292:64]
  assign io_stream_in_183_ready = merger_io_stream_in_183_ready; // @[Stab.scala 292:64]
  assign io_stream_in_184_ready = merger_io_stream_in_184_ready; // @[Stab.scala 292:64]
  assign io_stream_in_185_ready = merger_io_stream_in_185_ready; // @[Stab.scala 292:64]
  assign io_stream_in_186_ready = merger_io_stream_in_186_ready; // @[Stab.scala 292:64]
  assign io_stream_in_187_ready = merger_io_stream_in_187_ready; // @[Stab.scala 292:64]
  assign io_stream_in_188_ready = merger_io_stream_in_188_ready; // @[Stab.scala 292:64]
  assign io_stream_in_189_ready = merger_io_stream_in_189_ready; // @[Stab.scala 292:64]
  assign io_stream_in_190_ready = merger_io_stream_in_190_ready; // @[Stab.scala 292:64]
  assign io_stream_in_191_ready = merger_io_stream_in_191_ready; // @[Stab.scala 292:64]
  assign io_stream_in_192_ready = merger_io_stream_in_192_ready; // @[Stab.scala 292:64]
  assign io_stream_in_193_ready = merger_io_stream_in_193_ready; // @[Stab.scala 292:64]
  assign io_stream_in_194_ready = merger_io_stream_in_194_ready; // @[Stab.scala 292:64]
  assign io_stream_in_195_ready = merger_io_stream_in_195_ready; // @[Stab.scala 292:64]
  assign io_stream_in_196_ready = merger_io_stream_in_196_ready; // @[Stab.scala 292:64]
  assign io_stream_in_197_ready = merger_io_stream_in_197_ready; // @[Stab.scala 292:64]
  assign io_stream_in_198_ready = merger_io_stream_in_198_ready; // @[Stab.scala 292:64]
  assign io_stream_in_199_ready = merger_io_stream_in_199_ready; // @[Stab.scala 292:64]
  assign io_stream_in_200_ready = merger_io_stream_in_200_ready; // @[Stab.scala 292:64]
  assign io_stream_in_201_ready = merger_io_stream_in_201_ready; // @[Stab.scala 292:64]
  assign io_stream_in_202_ready = merger_io_stream_in_202_ready; // @[Stab.scala 292:64]
  assign io_stream_in_203_ready = merger_io_stream_in_203_ready; // @[Stab.scala 292:64]
  assign io_stream_in_204_ready = merger_io_stream_in_204_ready; // @[Stab.scala 292:64]
  assign io_stream_in_205_ready = merger_io_stream_in_205_ready; // @[Stab.scala 292:64]
  assign io_stream_in_206_ready = merger_io_stream_in_206_ready; // @[Stab.scala 292:64]
  assign io_stream_in_207_ready = merger_io_stream_in_207_ready; // @[Stab.scala 292:64]
  assign io_stream_in_208_ready = merger_io_stream_in_208_ready; // @[Stab.scala 292:64]
  assign io_stream_in_209_ready = merger_io_stream_in_209_ready; // @[Stab.scala 292:64]
  assign io_stream_in_210_ready = merger_io_stream_in_210_ready; // @[Stab.scala 292:64]
  assign io_stream_in_211_ready = merger_io_stream_in_211_ready; // @[Stab.scala 292:64]
  assign io_stream_in_212_ready = merger_io_stream_in_212_ready; // @[Stab.scala 292:64]
  assign io_stream_in_213_ready = merger_io_stream_in_213_ready; // @[Stab.scala 292:64]
  assign io_stream_in_214_ready = merger_io_stream_in_214_ready; // @[Stab.scala 292:64]
  assign io_stream_in_215_ready = merger_io_stream_in_215_ready; // @[Stab.scala 292:64]
  assign io_stream_in_216_ready = merger_io_stream_in_216_ready; // @[Stab.scala 292:64]
  assign io_stream_in_217_ready = merger_io_stream_in_217_ready; // @[Stab.scala 292:64]
  assign io_stream_in_218_ready = merger_io_stream_in_218_ready; // @[Stab.scala 292:64]
  assign io_stream_in_219_ready = merger_io_stream_in_219_ready; // @[Stab.scala 292:64]
  assign io_stream_in_220_ready = merger_io_stream_in_220_ready; // @[Stab.scala 292:64]
  assign io_stream_in_221_ready = merger_io_stream_in_221_ready; // @[Stab.scala 292:64]
  assign io_stream_in_222_ready = merger_io_stream_in_222_ready; // @[Stab.scala 292:64]
  assign io_stream_in_223_ready = merger_io_stream_in_223_ready; // @[Stab.scala 292:64]
  assign io_stream_in_224_ready = merger_io_stream_in_224_ready; // @[Stab.scala 292:64]
  assign io_stream_in_225_ready = merger_io_stream_in_225_ready; // @[Stab.scala 292:64]
  assign io_stream_in_226_ready = merger_io_stream_in_226_ready; // @[Stab.scala 292:64]
  assign io_stream_in_227_ready = merger_io_stream_in_227_ready; // @[Stab.scala 292:64]
  assign io_stream_in_228_ready = merger_io_stream_in_228_ready; // @[Stab.scala 292:64]
  assign io_stream_in_229_ready = merger_io_stream_in_229_ready; // @[Stab.scala 292:64]
  assign io_stream_in_230_ready = merger_io_stream_in_230_ready; // @[Stab.scala 292:64]
  assign io_stream_in_231_ready = merger_io_stream_in_231_ready; // @[Stab.scala 292:64]
  assign io_stream_in_232_ready = merger_io_stream_in_232_ready; // @[Stab.scala 292:64]
  assign io_stream_in_233_ready = merger_io_stream_in_233_ready; // @[Stab.scala 292:64]
  assign io_stream_in_234_ready = merger_io_stream_in_234_ready; // @[Stab.scala 292:64]
  assign io_stream_in_235_ready = merger_io_stream_in_235_ready; // @[Stab.scala 292:64]
  assign io_stream_in_236_ready = merger_io_stream_in_236_ready; // @[Stab.scala 292:64]
  assign io_stream_in_237_ready = merger_io_stream_in_237_ready; // @[Stab.scala 292:64]
  assign io_stream_in_238_ready = merger_io_stream_in_238_ready; // @[Stab.scala 292:64]
  assign io_stream_in_239_ready = merger_io_stream_in_239_ready; // @[Stab.scala 292:64]
  assign io_stream_in_240_ready = merger_io_stream_in_240_ready; // @[Stab.scala 292:64]
  assign io_stream_in_241_ready = merger_io_stream_in_241_ready; // @[Stab.scala 292:64]
  assign io_stream_in_242_ready = merger_io_stream_in_242_ready; // @[Stab.scala 292:64]
  assign io_stream_in_243_ready = merger_io_stream_in_243_ready; // @[Stab.scala 292:64]
  assign io_stream_in_244_ready = merger_io_stream_in_244_ready; // @[Stab.scala 292:64]
  assign io_stream_in_245_ready = merger_io_stream_in_245_ready; // @[Stab.scala 292:64]
  assign io_stream_in_246_ready = merger_io_stream_in_246_ready; // @[Stab.scala 292:64]
  assign io_stream_in_247_ready = merger_io_stream_in_247_ready; // @[Stab.scala 292:64]
  assign io_stream_in_248_ready = merger_io_stream_in_248_ready; // @[Stab.scala 292:64]
  assign io_stream_in_249_ready = merger_io_stream_in_249_ready; // @[Stab.scala 292:64]
  assign io_stream_in_250_ready = merger_io_stream_in_250_ready; // @[Stab.scala 292:64]
  assign io_stream_in_251_ready = merger_io_stream_in_251_ready; // @[Stab.scala 292:64]
  assign io_stream_in_252_ready = merger_io_stream_in_252_ready; // @[Stab.scala 292:64]
  assign io_stream_in_253_ready = merger_io_stream_in_253_ready; // @[Stab.scala 292:64]
  assign io_stream_in_254_ready = merger_io_stream_in_254_ready; // @[Stab.scala 292:64]
  assign io_stream_in_255_ready = merger_io_stream_in_255_ready; // @[Stab.scala 292:64]
  assign io_stream_out_valid = merger_io_stream_out_valid; // @[Stab.scala 294:17]
  assign io_stream_out_bits = merger_io_stream_out_bits; // @[Stab.scala 294:17]
  assign merger_clock = clock;
  assign merger_reset = reset;
  assign merger_io_stream_in_0_valid = io_stream_in_0_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_0_bits = io_stream_in_0_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_1_valid = io_stream_in_1_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_1_bits = io_stream_in_1_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_2_valid = io_stream_in_2_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_2_bits = io_stream_in_2_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_3_valid = io_stream_in_3_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_3_bits = io_stream_in_3_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_4_valid = io_stream_in_4_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_4_bits = io_stream_in_4_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_5_valid = io_stream_in_5_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_5_bits = io_stream_in_5_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_6_valid = io_stream_in_6_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_6_bits = io_stream_in_6_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_7_valid = io_stream_in_7_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_7_bits = io_stream_in_7_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_8_valid = io_stream_in_8_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_8_bits = io_stream_in_8_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_9_valid = io_stream_in_9_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_9_bits = io_stream_in_9_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_10_valid = io_stream_in_10_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_10_bits = io_stream_in_10_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_11_valid = io_stream_in_11_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_11_bits = io_stream_in_11_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_12_valid = io_stream_in_12_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_12_bits = io_stream_in_12_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_13_valid = io_stream_in_13_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_13_bits = io_stream_in_13_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_14_valid = io_stream_in_14_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_14_bits = io_stream_in_14_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_15_valid = io_stream_in_15_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_15_bits = io_stream_in_15_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_16_valid = io_stream_in_16_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_16_bits = io_stream_in_16_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_17_valid = io_stream_in_17_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_17_bits = io_stream_in_17_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_18_valid = io_stream_in_18_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_18_bits = io_stream_in_18_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_19_valid = io_stream_in_19_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_19_bits = io_stream_in_19_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_20_valid = io_stream_in_20_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_20_bits = io_stream_in_20_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_21_valid = io_stream_in_21_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_21_bits = io_stream_in_21_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_22_valid = io_stream_in_22_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_22_bits = io_stream_in_22_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_23_valid = io_stream_in_23_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_23_bits = io_stream_in_23_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_24_valid = io_stream_in_24_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_24_bits = io_stream_in_24_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_25_valid = io_stream_in_25_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_25_bits = io_stream_in_25_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_26_valid = io_stream_in_26_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_26_bits = io_stream_in_26_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_27_valid = io_stream_in_27_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_27_bits = io_stream_in_27_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_28_valid = io_stream_in_28_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_28_bits = io_stream_in_28_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_29_valid = io_stream_in_29_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_29_bits = io_stream_in_29_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_30_valid = io_stream_in_30_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_30_bits = io_stream_in_30_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_31_valid = io_stream_in_31_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_31_bits = io_stream_in_31_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_32_valid = io_stream_in_32_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_32_bits = io_stream_in_32_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_33_valid = io_stream_in_33_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_33_bits = io_stream_in_33_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_34_valid = io_stream_in_34_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_34_bits = io_stream_in_34_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_35_valid = io_stream_in_35_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_35_bits = io_stream_in_35_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_36_valid = io_stream_in_36_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_36_bits = io_stream_in_36_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_37_valid = io_stream_in_37_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_37_bits = io_stream_in_37_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_38_valid = io_stream_in_38_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_38_bits = io_stream_in_38_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_39_valid = io_stream_in_39_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_39_bits = io_stream_in_39_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_40_valid = io_stream_in_40_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_40_bits = io_stream_in_40_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_41_valid = io_stream_in_41_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_41_bits = io_stream_in_41_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_42_valid = io_stream_in_42_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_42_bits = io_stream_in_42_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_43_valid = io_stream_in_43_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_43_bits = io_stream_in_43_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_44_valid = io_stream_in_44_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_44_bits = io_stream_in_44_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_45_valid = io_stream_in_45_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_45_bits = io_stream_in_45_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_46_valid = io_stream_in_46_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_46_bits = io_stream_in_46_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_47_valid = io_stream_in_47_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_47_bits = io_stream_in_47_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_48_valid = io_stream_in_48_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_48_bits = io_stream_in_48_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_49_valid = io_stream_in_49_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_49_bits = io_stream_in_49_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_50_valid = io_stream_in_50_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_50_bits = io_stream_in_50_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_51_valid = io_stream_in_51_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_51_bits = io_stream_in_51_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_52_valid = io_stream_in_52_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_52_bits = io_stream_in_52_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_53_valid = io_stream_in_53_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_53_bits = io_stream_in_53_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_54_valid = io_stream_in_54_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_54_bits = io_stream_in_54_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_55_valid = io_stream_in_55_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_55_bits = io_stream_in_55_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_56_valid = io_stream_in_56_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_56_bits = io_stream_in_56_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_57_valid = io_stream_in_57_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_57_bits = io_stream_in_57_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_58_valid = io_stream_in_58_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_58_bits = io_stream_in_58_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_59_valid = io_stream_in_59_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_59_bits = io_stream_in_59_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_60_valid = io_stream_in_60_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_60_bits = io_stream_in_60_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_61_valid = io_stream_in_61_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_61_bits = io_stream_in_61_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_62_valid = io_stream_in_62_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_62_bits = io_stream_in_62_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_63_valid = io_stream_in_63_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_63_bits = io_stream_in_63_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_64_valid = io_stream_in_64_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_64_bits = io_stream_in_64_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_65_valid = io_stream_in_65_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_65_bits = io_stream_in_65_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_66_valid = io_stream_in_66_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_66_bits = io_stream_in_66_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_67_valid = io_stream_in_67_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_67_bits = io_stream_in_67_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_68_valid = io_stream_in_68_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_68_bits = io_stream_in_68_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_69_valid = io_stream_in_69_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_69_bits = io_stream_in_69_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_70_valid = io_stream_in_70_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_70_bits = io_stream_in_70_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_71_valid = io_stream_in_71_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_71_bits = io_stream_in_71_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_72_valid = io_stream_in_72_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_72_bits = io_stream_in_72_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_73_valid = io_stream_in_73_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_73_bits = io_stream_in_73_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_74_valid = io_stream_in_74_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_74_bits = io_stream_in_74_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_75_valid = io_stream_in_75_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_75_bits = io_stream_in_75_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_76_valid = io_stream_in_76_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_76_bits = io_stream_in_76_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_77_valid = io_stream_in_77_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_77_bits = io_stream_in_77_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_78_valid = io_stream_in_78_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_78_bits = io_stream_in_78_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_79_valid = io_stream_in_79_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_79_bits = io_stream_in_79_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_80_valid = io_stream_in_80_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_80_bits = io_stream_in_80_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_81_valid = io_stream_in_81_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_81_bits = io_stream_in_81_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_82_valid = io_stream_in_82_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_82_bits = io_stream_in_82_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_83_valid = io_stream_in_83_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_83_bits = io_stream_in_83_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_84_valid = io_stream_in_84_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_84_bits = io_stream_in_84_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_85_valid = io_stream_in_85_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_85_bits = io_stream_in_85_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_86_valid = io_stream_in_86_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_86_bits = io_stream_in_86_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_87_valid = io_stream_in_87_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_87_bits = io_stream_in_87_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_88_valid = io_stream_in_88_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_88_bits = io_stream_in_88_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_89_valid = io_stream_in_89_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_89_bits = io_stream_in_89_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_90_valid = io_stream_in_90_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_90_bits = io_stream_in_90_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_91_valid = io_stream_in_91_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_91_bits = io_stream_in_91_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_92_valid = io_stream_in_92_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_92_bits = io_stream_in_92_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_93_valid = io_stream_in_93_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_93_bits = io_stream_in_93_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_94_valid = io_stream_in_94_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_94_bits = io_stream_in_94_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_95_valid = io_stream_in_95_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_95_bits = io_stream_in_95_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_96_valid = io_stream_in_96_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_96_bits = io_stream_in_96_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_97_valid = io_stream_in_97_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_97_bits = io_stream_in_97_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_98_valid = io_stream_in_98_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_98_bits = io_stream_in_98_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_99_valid = io_stream_in_99_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_99_bits = io_stream_in_99_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_100_valid = io_stream_in_100_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_100_bits = io_stream_in_100_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_101_valid = io_stream_in_101_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_101_bits = io_stream_in_101_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_102_valid = io_stream_in_102_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_102_bits = io_stream_in_102_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_103_valid = io_stream_in_103_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_103_bits = io_stream_in_103_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_104_valid = io_stream_in_104_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_104_bits = io_stream_in_104_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_105_valid = io_stream_in_105_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_105_bits = io_stream_in_105_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_106_valid = io_stream_in_106_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_106_bits = io_stream_in_106_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_107_valid = io_stream_in_107_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_107_bits = io_stream_in_107_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_108_valid = io_stream_in_108_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_108_bits = io_stream_in_108_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_109_valid = io_stream_in_109_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_109_bits = io_stream_in_109_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_110_valid = io_stream_in_110_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_110_bits = io_stream_in_110_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_111_valid = io_stream_in_111_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_111_bits = io_stream_in_111_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_112_valid = io_stream_in_112_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_112_bits = io_stream_in_112_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_113_valid = io_stream_in_113_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_113_bits = io_stream_in_113_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_114_valid = io_stream_in_114_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_114_bits = io_stream_in_114_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_115_valid = io_stream_in_115_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_115_bits = io_stream_in_115_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_116_valid = io_stream_in_116_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_116_bits = io_stream_in_116_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_117_valid = io_stream_in_117_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_117_bits = io_stream_in_117_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_118_valid = io_stream_in_118_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_118_bits = io_stream_in_118_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_119_valid = io_stream_in_119_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_119_bits = io_stream_in_119_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_120_valid = io_stream_in_120_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_120_bits = io_stream_in_120_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_121_valid = io_stream_in_121_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_121_bits = io_stream_in_121_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_122_valid = io_stream_in_122_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_122_bits = io_stream_in_122_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_123_valid = io_stream_in_123_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_123_bits = io_stream_in_123_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_124_valid = io_stream_in_124_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_124_bits = io_stream_in_124_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_125_valid = io_stream_in_125_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_125_bits = io_stream_in_125_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_126_valid = io_stream_in_126_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_126_bits = io_stream_in_126_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_127_valid = io_stream_in_127_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_127_bits = io_stream_in_127_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_128_valid = io_stream_in_128_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_128_bits = io_stream_in_128_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_129_valid = io_stream_in_129_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_129_bits = io_stream_in_129_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_130_valid = io_stream_in_130_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_130_bits = io_stream_in_130_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_131_valid = io_stream_in_131_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_131_bits = io_stream_in_131_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_132_valid = io_stream_in_132_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_132_bits = io_stream_in_132_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_133_valid = io_stream_in_133_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_133_bits = io_stream_in_133_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_134_valid = io_stream_in_134_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_134_bits = io_stream_in_134_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_135_valid = io_stream_in_135_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_135_bits = io_stream_in_135_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_136_valid = io_stream_in_136_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_136_bits = io_stream_in_136_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_137_valid = io_stream_in_137_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_137_bits = io_stream_in_137_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_138_valid = io_stream_in_138_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_138_bits = io_stream_in_138_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_139_valid = io_stream_in_139_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_139_bits = io_stream_in_139_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_140_valid = io_stream_in_140_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_140_bits = io_stream_in_140_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_141_valid = io_stream_in_141_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_141_bits = io_stream_in_141_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_142_valid = io_stream_in_142_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_142_bits = io_stream_in_142_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_143_valid = io_stream_in_143_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_143_bits = io_stream_in_143_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_144_valid = io_stream_in_144_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_144_bits = io_stream_in_144_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_145_valid = io_stream_in_145_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_145_bits = io_stream_in_145_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_146_valid = io_stream_in_146_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_146_bits = io_stream_in_146_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_147_valid = io_stream_in_147_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_147_bits = io_stream_in_147_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_148_valid = io_stream_in_148_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_148_bits = io_stream_in_148_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_149_valid = io_stream_in_149_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_149_bits = io_stream_in_149_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_150_valid = io_stream_in_150_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_150_bits = io_stream_in_150_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_151_valid = io_stream_in_151_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_151_bits = io_stream_in_151_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_152_valid = io_stream_in_152_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_152_bits = io_stream_in_152_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_153_valid = io_stream_in_153_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_153_bits = io_stream_in_153_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_154_valid = io_stream_in_154_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_154_bits = io_stream_in_154_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_155_valid = io_stream_in_155_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_155_bits = io_stream_in_155_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_156_valid = io_stream_in_156_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_156_bits = io_stream_in_156_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_157_valid = io_stream_in_157_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_157_bits = io_stream_in_157_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_158_valid = io_stream_in_158_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_158_bits = io_stream_in_158_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_159_valid = io_stream_in_159_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_159_bits = io_stream_in_159_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_160_valid = io_stream_in_160_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_160_bits = io_stream_in_160_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_161_valid = io_stream_in_161_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_161_bits = io_stream_in_161_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_162_valid = io_stream_in_162_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_162_bits = io_stream_in_162_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_163_valid = io_stream_in_163_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_163_bits = io_stream_in_163_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_164_valid = io_stream_in_164_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_164_bits = io_stream_in_164_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_165_valid = io_stream_in_165_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_165_bits = io_stream_in_165_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_166_valid = io_stream_in_166_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_166_bits = io_stream_in_166_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_167_valid = io_stream_in_167_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_167_bits = io_stream_in_167_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_168_valid = io_stream_in_168_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_168_bits = io_stream_in_168_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_169_valid = io_stream_in_169_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_169_bits = io_stream_in_169_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_170_valid = io_stream_in_170_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_170_bits = io_stream_in_170_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_171_valid = io_stream_in_171_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_171_bits = io_stream_in_171_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_172_valid = io_stream_in_172_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_172_bits = io_stream_in_172_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_173_valid = io_stream_in_173_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_173_bits = io_stream_in_173_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_174_valid = io_stream_in_174_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_174_bits = io_stream_in_174_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_175_valid = io_stream_in_175_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_175_bits = io_stream_in_175_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_176_valid = io_stream_in_176_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_176_bits = io_stream_in_176_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_177_valid = io_stream_in_177_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_177_bits = io_stream_in_177_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_178_valid = io_stream_in_178_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_178_bits = io_stream_in_178_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_179_valid = io_stream_in_179_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_179_bits = io_stream_in_179_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_180_valid = io_stream_in_180_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_180_bits = io_stream_in_180_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_181_valid = io_stream_in_181_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_181_bits = io_stream_in_181_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_182_valid = io_stream_in_182_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_182_bits = io_stream_in_182_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_183_valid = io_stream_in_183_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_183_bits = io_stream_in_183_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_184_valid = io_stream_in_184_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_184_bits = io_stream_in_184_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_185_valid = io_stream_in_185_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_185_bits = io_stream_in_185_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_186_valid = io_stream_in_186_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_186_bits = io_stream_in_186_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_187_valid = io_stream_in_187_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_187_bits = io_stream_in_187_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_188_valid = io_stream_in_188_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_188_bits = io_stream_in_188_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_189_valid = io_stream_in_189_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_189_bits = io_stream_in_189_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_190_valid = io_stream_in_190_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_190_bits = io_stream_in_190_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_191_valid = io_stream_in_191_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_191_bits = io_stream_in_191_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_192_valid = io_stream_in_192_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_192_bits = io_stream_in_192_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_193_valid = io_stream_in_193_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_193_bits = io_stream_in_193_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_194_valid = io_stream_in_194_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_194_bits = io_stream_in_194_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_195_valid = io_stream_in_195_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_195_bits = io_stream_in_195_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_196_valid = io_stream_in_196_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_196_bits = io_stream_in_196_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_197_valid = io_stream_in_197_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_197_bits = io_stream_in_197_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_198_valid = io_stream_in_198_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_198_bits = io_stream_in_198_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_199_valid = io_stream_in_199_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_199_bits = io_stream_in_199_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_200_valid = io_stream_in_200_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_200_bits = io_stream_in_200_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_201_valid = io_stream_in_201_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_201_bits = io_stream_in_201_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_202_valid = io_stream_in_202_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_202_bits = io_stream_in_202_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_203_valid = io_stream_in_203_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_203_bits = io_stream_in_203_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_204_valid = io_stream_in_204_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_204_bits = io_stream_in_204_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_205_valid = io_stream_in_205_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_205_bits = io_stream_in_205_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_206_valid = io_stream_in_206_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_206_bits = io_stream_in_206_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_207_valid = io_stream_in_207_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_207_bits = io_stream_in_207_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_208_valid = io_stream_in_208_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_208_bits = io_stream_in_208_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_209_valid = io_stream_in_209_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_209_bits = io_stream_in_209_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_210_valid = io_stream_in_210_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_210_bits = io_stream_in_210_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_211_valid = io_stream_in_211_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_211_bits = io_stream_in_211_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_212_valid = io_stream_in_212_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_212_bits = io_stream_in_212_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_213_valid = io_stream_in_213_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_213_bits = io_stream_in_213_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_214_valid = io_stream_in_214_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_214_bits = io_stream_in_214_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_215_valid = io_stream_in_215_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_215_bits = io_stream_in_215_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_216_valid = io_stream_in_216_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_216_bits = io_stream_in_216_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_217_valid = io_stream_in_217_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_217_bits = io_stream_in_217_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_218_valid = io_stream_in_218_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_218_bits = io_stream_in_218_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_219_valid = io_stream_in_219_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_219_bits = io_stream_in_219_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_220_valid = io_stream_in_220_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_220_bits = io_stream_in_220_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_221_valid = io_stream_in_221_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_221_bits = io_stream_in_221_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_222_valid = io_stream_in_222_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_222_bits = io_stream_in_222_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_223_valid = io_stream_in_223_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_223_bits = io_stream_in_223_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_224_valid = io_stream_in_224_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_224_bits = io_stream_in_224_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_225_valid = io_stream_in_225_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_225_bits = io_stream_in_225_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_226_valid = io_stream_in_226_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_226_bits = io_stream_in_226_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_227_valid = io_stream_in_227_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_227_bits = io_stream_in_227_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_228_valid = io_stream_in_228_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_228_bits = io_stream_in_228_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_229_valid = io_stream_in_229_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_229_bits = io_stream_in_229_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_230_valid = io_stream_in_230_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_230_bits = io_stream_in_230_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_231_valid = io_stream_in_231_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_231_bits = io_stream_in_231_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_232_valid = io_stream_in_232_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_232_bits = io_stream_in_232_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_233_valid = io_stream_in_233_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_233_bits = io_stream_in_233_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_234_valid = io_stream_in_234_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_234_bits = io_stream_in_234_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_235_valid = io_stream_in_235_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_235_bits = io_stream_in_235_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_236_valid = io_stream_in_236_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_236_bits = io_stream_in_236_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_237_valid = io_stream_in_237_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_237_bits = io_stream_in_237_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_238_valid = io_stream_in_238_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_238_bits = io_stream_in_238_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_239_valid = io_stream_in_239_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_239_bits = io_stream_in_239_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_240_valid = io_stream_in_240_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_240_bits = io_stream_in_240_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_241_valid = io_stream_in_241_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_241_bits = io_stream_in_241_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_242_valid = io_stream_in_242_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_242_bits = io_stream_in_242_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_243_valid = io_stream_in_243_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_243_bits = io_stream_in_243_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_244_valid = io_stream_in_244_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_244_bits = io_stream_in_244_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_245_valid = io_stream_in_245_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_245_bits = io_stream_in_245_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_246_valid = io_stream_in_246_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_246_bits = io_stream_in_246_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_247_valid = io_stream_in_247_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_247_bits = io_stream_in_247_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_248_valid = io_stream_in_248_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_248_bits = io_stream_in_248_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_249_valid = io_stream_in_249_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_249_bits = io_stream_in_249_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_250_valid = io_stream_in_250_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_250_bits = io_stream_in_250_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_251_valid = io_stream_in_251_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_251_bits = io_stream_in_251_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_252_valid = io_stream_in_252_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_252_bits = io_stream_in_252_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_253_valid = io_stream_in_253_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_253_bits = io_stream_in_253_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_254_valid = io_stream_in_254_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_254_bits = io_stream_in_254_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_in_255_valid = io_stream_in_255_valid; // @[Stab.scala 292:64]
  assign merger_io_stream_in_255_bits = io_stream_in_255_bits; // @[Stab.scala 292:64]
  assign merger_io_stream_out_ready = io_stream_out_ready; // @[Stab.scala 294:17]
endmodule
module MatrixMultiplierStreaming(
  input         clock,
  input         reset,
  output        io_value_in_ready,
  input         io_value_in_valid,
  input  [31:0] io_value_in_bits,
  output        io_weight_in_ready,
  input         io_weight_in_valid,
  input  [31:0] io_weight_in_bits,
  input         io_value_out_ready,
  output        io_value_out_valid,
  output [31:0] io_value_out_bits
);
  wire  core_clock; // @[Stab.scala 312:20]
  wire  core_reset; // @[Stab.scala 312:20]
  wire  core_io_weight_in_0_ready; // @[Stab.scala 312:20]
  wire  core_io_weight_in_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_weight_in_0_bits; // @[Stab.scala 312:20]
  wire  core_io_weight_in_1_ready; // @[Stab.scala 312:20]
  wire  core_io_weight_in_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_weight_in_1_bits; // @[Stab.scala 312:20]
  wire  core_io_weight_in_2_ready; // @[Stab.scala 312:20]
  wire  core_io_weight_in_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_weight_in_2_bits; // @[Stab.scala 312:20]
  wire  core_io_weight_in_3_ready; // @[Stab.scala 312:20]
  wire  core_io_weight_in_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_weight_in_3_bits; // @[Stab.scala 312:20]
  wire  core_io_weight_in_4_ready; // @[Stab.scala 312:20]
  wire  core_io_weight_in_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_weight_in_4_bits; // @[Stab.scala 312:20]
  wire  core_io_weight_in_5_ready; // @[Stab.scala 312:20]
  wire  core_io_weight_in_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_weight_in_5_bits; // @[Stab.scala 312:20]
  wire  core_io_weight_in_6_ready; // @[Stab.scala 312:20]
  wire  core_io_weight_in_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_weight_in_6_bits; // @[Stab.scala 312:20]
  wire  core_io_weight_in_7_ready; // @[Stab.scala 312:20]
  wire  core_io_weight_in_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_weight_in_7_bits; // @[Stab.scala 312:20]
  wire  core_io_weight_in_8_ready; // @[Stab.scala 312:20]
  wire  core_io_weight_in_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_weight_in_8_bits; // @[Stab.scala 312:20]
  wire  core_io_weight_in_9_ready; // @[Stab.scala 312:20]
  wire  core_io_weight_in_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_weight_in_9_bits; // @[Stab.scala 312:20]
  wire  core_io_weight_in_10_ready; // @[Stab.scala 312:20]
  wire  core_io_weight_in_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_weight_in_10_bits; // @[Stab.scala 312:20]
  wire  core_io_weight_in_11_ready; // @[Stab.scala 312:20]
  wire  core_io_weight_in_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_weight_in_11_bits; // @[Stab.scala 312:20]
  wire  core_io_weight_in_12_ready; // @[Stab.scala 312:20]
  wire  core_io_weight_in_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_weight_in_12_bits; // @[Stab.scala 312:20]
  wire  core_io_weight_in_13_ready; // @[Stab.scala 312:20]
  wire  core_io_weight_in_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_weight_in_13_bits; // @[Stab.scala 312:20]
  wire  core_io_weight_in_14_ready; // @[Stab.scala 312:20]
  wire  core_io_weight_in_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_weight_in_14_bits; // @[Stab.scala 312:20]
  wire  core_io_weight_in_15_ready; // @[Stab.scala 312:20]
  wire  core_io_weight_in_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_weight_in_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_in_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_in_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_in_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_in_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_in_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_in_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_in_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_in_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_in_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_in_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_in_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_in_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_in_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_in_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_in_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_in_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_in_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_in_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_in_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_in_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_in_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_in_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_in_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_in_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_in_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_in_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_in_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_in_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_in_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_in_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_in_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_in_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_in_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_in_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_in_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_in_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_in_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_in_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_in_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_in_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_in_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_in_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_in_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_in_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_in_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_in_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_in_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_in_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_0_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_0_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_0_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_0_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_0_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_0_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_0_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_0_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_0_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_0_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_0_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_0_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_0_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_0_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_0_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_0_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_0_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_1_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_1_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_1_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_1_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_1_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_1_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_1_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_1_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_1_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_1_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_1_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_1_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_1_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_1_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_1_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_1_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_1_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_2_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_2_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_2_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_2_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_2_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_2_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_2_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_2_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_2_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_2_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_2_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_2_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_2_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_2_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_2_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_2_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_2_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_3_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_3_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_3_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_3_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_3_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_3_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_3_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_3_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_3_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_3_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_3_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_3_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_3_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_3_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_3_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_3_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_3_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_4_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_4_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_4_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_4_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_4_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_4_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_4_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_4_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_4_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_4_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_4_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_4_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_4_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_4_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_4_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_4_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_4_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_5_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_5_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_5_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_5_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_5_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_5_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_5_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_5_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_5_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_5_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_5_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_5_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_5_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_5_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_5_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_5_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_5_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_6_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_6_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_6_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_6_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_6_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_6_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_6_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_6_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_6_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_6_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_6_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_6_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_6_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_6_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_6_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_6_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_6_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_7_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_7_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_7_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_7_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_7_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_7_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_7_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_7_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_7_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_7_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_7_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_7_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_7_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_7_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_7_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_7_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_7_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_8_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_8_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_8_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_8_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_8_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_8_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_8_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_8_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_8_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_8_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_8_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_8_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_8_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_8_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_8_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_8_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_8_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_9_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_9_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_9_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_9_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_9_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_9_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_9_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_9_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_9_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_9_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_9_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_9_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_9_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_9_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_9_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_9_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_9_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_10_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_10_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_10_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_10_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_10_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_10_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_10_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_10_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_10_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_10_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_10_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_10_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_10_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_10_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_10_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_10_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_10_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_11_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_11_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_11_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_11_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_11_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_11_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_11_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_11_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_11_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_11_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_11_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_11_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_11_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_11_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_11_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_11_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_11_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_12_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_12_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_12_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_12_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_12_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_12_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_12_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_12_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_12_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_12_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_12_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_12_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_12_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_12_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_12_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_12_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_12_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_13_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_13_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_13_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_13_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_13_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_13_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_13_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_13_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_13_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_13_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_13_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_13_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_13_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_13_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_13_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_13_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_13_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_14_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_14_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_14_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_14_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_14_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_14_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_14_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_14_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_14_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_14_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_14_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_14_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_14_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_14_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_14_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_14_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_14_15_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_0_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_0_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_15_0_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_1_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_1_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_15_1_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_2_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_2_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_15_2_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_3_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_3_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_15_3_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_4_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_4_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_15_4_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_5_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_5_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_15_5_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_6_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_6_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_15_6_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_7_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_7_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_15_7_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_8_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_8_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_15_8_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_9_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_9_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_15_9_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_10_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_10_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_15_10_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_11_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_11_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_15_11_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_12_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_12_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_15_12_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_13_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_13_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_15_13_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_14_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_14_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_15_14_bits; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_15_ready; // @[Stab.scala 312:20]
  wire  core_io_value_out_15_15_valid; // @[Stab.scala 312:20]
  wire [31:0] core_io_value_out_15_15_bits; // @[Stab.scala 312:20]
  wire  wsplit_clock; // @[Stab.scala 314:22]
  wire  wsplit_reset; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_in_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_in_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_in_bits; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_0_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_0_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_out_0_bits; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_1_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_1_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_out_1_bits; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_2_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_2_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_out_2_bits; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_3_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_3_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_out_3_bits; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_4_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_4_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_out_4_bits; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_5_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_5_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_out_5_bits; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_6_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_6_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_out_6_bits; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_7_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_7_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_out_7_bits; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_8_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_8_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_out_8_bits; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_9_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_9_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_out_9_bits; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_10_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_10_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_out_10_bits; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_11_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_11_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_out_11_bits; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_12_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_12_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_out_12_bits; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_13_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_13_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_out_13_bits; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_14_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_14_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_out_14_bits; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_15_ready; // @[Stab.scala 314:22]
  wire  wsplit_io_stream_out_15_valid; // @[Stab.scala 314:22]
  wire [31:0] wsplit_io_stream_out_15_bits; // @[Stab.scala 314:22]
  wire  vsplit_clock; // @[Stab.scala 315:22]
  wire  vsplit_reset; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_in_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_in_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_in_bits; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_0_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_0_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_out_0_bits; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_1_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_1_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_out_1_bits; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_2_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_2_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_out_2_bits; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_3_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_3_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_out_3_bits; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_4_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_4_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_out_4_bits; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_5_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_5_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_out_5_bits; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_6_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_6_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_out_6_bits; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_7_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_7_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_out_7_bits; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_8_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_8_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_out_8_bits; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_9_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_9_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_out_9_bits; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_10_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_10_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_out_10_bits; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_11_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_11_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_out_11_bits; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_12_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_12_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_out_12_bits; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_13_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_13_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_out_13_bits; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_14_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_14_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_out_14_bits; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_15_ready; // @[Stab.scala 315:22]
  wire  vsplit_io_stream_out_15_valid; // @[Stab.scala 315:22]
  wire [31:0] vsplit_io_stream_out_15_bits; // @[Stab.scala 315:22]
  wire  rmerge_clock; // @[Stab.scala 317:22]
  wire  rmerge_reset; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_0_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_0_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_0_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_1_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_1_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_1_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_2_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_2_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_2_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_3_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_3_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_3_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_4_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_4_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_4_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_5_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_5_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_5_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_6_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_6_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_6_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_7_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_7_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_7_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_8_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_8_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_8_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_9_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_9_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_9_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_10_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_10_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_10_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_11_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_11_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_11_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_12_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_12_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_12_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_13_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_13_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_13_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_14_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_14_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_14_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_15_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_15_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_15_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_16_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_16_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_16_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_17_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_17_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_17_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_18_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_18_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_18_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_19_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_19_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_19_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_20_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_20_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_20_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_21_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_21_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_21_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_22_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_22_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_22_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_23_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_23_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_23_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_24_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_24_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_24_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_25_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_25_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_25_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_26_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_26_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_26_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_27_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_27_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_27_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_28_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_28_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_28_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_29_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_29_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_29_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_30_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_30_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_30_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_31_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_31_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_31_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_32_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_32_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_32_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_33_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_33_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_33_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_34_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_34_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_34_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_35_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_35_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_35_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_36_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_36_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_36_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_37_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_37_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_37_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_38_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_38_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_38_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_39_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_39_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_39_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_40_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_40_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_40_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_41_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_41_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_41_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_42_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_42_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_42_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_43_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_43_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_43_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_44_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_44_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_44_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_45_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_45_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_45_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_46_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_46_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_46_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_47_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_47_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_47_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_48_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_48_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_48_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_49_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_49_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_49_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_50_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_50_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_50_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_51_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_51_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_51_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_52_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_52_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_52_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_53_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_53_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_53_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_54_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_54_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_54_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_55_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_55_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_55_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_56_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_56_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_56_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_57_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_57_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_57_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_58_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_58_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_58_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_59_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_59_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_59_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_60_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_60_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_60_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_61_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_61_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_61_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_62_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_62_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_62_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_63_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_63_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_63_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_64_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_64_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_64_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_65_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_65_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_65_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_66_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_66_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_66_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_67_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_67_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_67_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_68_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_68_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_68_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_69_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_69_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_69_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_70_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_70_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_70_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_71_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_71_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_71_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_72_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_72_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_72_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_73_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_73_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_73_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_74_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_74_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_74_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_75_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_75_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_75_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_76_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_76_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_76_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_77_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_77_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_77_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_78_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_78_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_78_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_79_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_79_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_79_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_80_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_80_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_80_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_81_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_81_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_81_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_82_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_82_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_82_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_83_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_83_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_83_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_84_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_84_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_84_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_85_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_85_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_85_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_86_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_86_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_86_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_87_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_87_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_87_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_88_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_88_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_88_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_89_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_89_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_89_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_90_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_90_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_90_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_91_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_91_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_91_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_92_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_92_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_92_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_93_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_93_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_93_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_94_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_94_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_94_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_95_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_95_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_95_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_96_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_96_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_96_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_97_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_97_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_97_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_98_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_98_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_98_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_99_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_99_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_99_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_100_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_100_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_100_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_101_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_101_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_101_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_102_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_102_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_102_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_103_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_103_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_103_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_104_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_104_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_104_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_105_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_105_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_105_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_106_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_106_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_106_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_107_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_107_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_107_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_108_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_108_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_108_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_109_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_109_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_109_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_110_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_110_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_110_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_111_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_111_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_111_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_112_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_112_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_112_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_113_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_113_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_113_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_114_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_114_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_114_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_115_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_115_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_115_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_116_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_116_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_116_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_117_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_117_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_117_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_118_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_118_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_118_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_119_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_119_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_119_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_120_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_120_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_120_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_121_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_121_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_121_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_122_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_122_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_122_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_123_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_123_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_123_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_124_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_124_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_124_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_125_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_125_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_125_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_126_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_126_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_126_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_127_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_127_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_127_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_128_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_128_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_128_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_129_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_129_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_129_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_130_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_130_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_130_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_131_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_131_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_131_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_132_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_132_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_132_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_133_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_133_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_133_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_134_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_134_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_134_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_135_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_135_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_135_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_136_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_136_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_136_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_137_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_137_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_137_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_138_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_138_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_138_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_139_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_139_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_139_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_140_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_140_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_140_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_141_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_141_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_141_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_142_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_142_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_142_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_143_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_143_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_143_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_144_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_144_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_144_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_145_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_145_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_145_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_146_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_146_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_146_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_147_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_147_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_147_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_148_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_148_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_148_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_149_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_149_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_149_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_150_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_150_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_150_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_151_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_151_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_151_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_152_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_152_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_152_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_153_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_153_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_153_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_154_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_154_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_154_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_155_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_155_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_155_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_156_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_156_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_156_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_157_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_157_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_157_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_158_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_158_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_158_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_159_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_159_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_159_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_160_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_160_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_160_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_161_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_161_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_161_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_162_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_162_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_162_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_163_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_163_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_163_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_164_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_164_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_164_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_165_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_165_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_165_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_166_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_166_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_166_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_167_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_167_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_167_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_168_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_168_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_168_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_169_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_169_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_169_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_170_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_170_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_170_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_171_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_171_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_171_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_172_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_172_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_172_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_173_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_173_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_173_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_174_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_174_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_174_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_175_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_175_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_175_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_176_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_176_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_176_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_177_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_177_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_177_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_178_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_178_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_178_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_179_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_179_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_179_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_180_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_180_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_180_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_181_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_181_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_181_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_182_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_182_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_182_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_183_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_183_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_183_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_184_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_184_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_184_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_185_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_185_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_185_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_186_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_186_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_186_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_187_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_187_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_187_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_188_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_188_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_188_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_189_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_189_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_189_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_190_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_190_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_190_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_191_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_191_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_191_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_192_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_192_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_192_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_193_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_193_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_193_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_194_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_194_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_194_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_195_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_195_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_195_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_196_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_196_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_196_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_197_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_197_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_197_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_198_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_198_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_198_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_199_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_199_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_199_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_200_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_200_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_200_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_201_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_201_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_201_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_202_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_202_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_202_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_203_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_203_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_203_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_204_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_204_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_204_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_205_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_205_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_205_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_206_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_206_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_206_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_207_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_207_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_207_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_208_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_208_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_208_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_209_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_209_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_209_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_210_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_210_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_210_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_211_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_211_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_211_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_212_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_212_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_212_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_213_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_213_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_213_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_214_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_214_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_214_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_215_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_215_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_215_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_216_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_216_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_216_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_217_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_217_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_217_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_218_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_218_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_218_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_219_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_219_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_219_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_220_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_220_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_220_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_221_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_221_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_221_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_222_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_222_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_222_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_223_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_223_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_223_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_224_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_224_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_224_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_225_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_225_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_225_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_226_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_226_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_226_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_227_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_227_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_227_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_228_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_228_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_228_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_229_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_229_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_229_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_230_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_230_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_230_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_231_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_231_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_231_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_232_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_232_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_232_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_233_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_233_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_233_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_234_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_234_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_234_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_235_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_235_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_235_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_236_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_236_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_236_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_237_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_237_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_237_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_238_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_238_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_238_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_239_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_239_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_239_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_240_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_240_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_240_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_241_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_241_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_241_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_242_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_242_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_242_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_243_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_243_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_243_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_244_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_244_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_244_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_245_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_245_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_245_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_246_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_246_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_246_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_247_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_247_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_247_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_248_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_248_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_248_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_249_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_249_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_249_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_250_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_250_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_250_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_251_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_251_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_251_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_252_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_252_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_252_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_253_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_253_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_253_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_254_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_254_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_254_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_255_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_in_255_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_in_255_bits; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_out_ready; // @[Stab.scala 317:22]
  wire  rmerge_io_stream_out_valid; // @[Stab.scala 317:22]
  wire [31:0] rmerge_io_stream_out_bits; // @[Stab.scala 317:22]
  BareMatrixMultiplier core ( // @[Stab.scala 312:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_weight_in_0_ready(core_io_weight_in_0_ready),
    .io_weight_in_0_valid(core_io_weight_in_0_valid),
    .io_weight_in_0_bits(core_io_weight_in_0_bits),
    .io_weight_in_1_ready(core_io_weight_in_1_ready),
    .io_weight_in_1_valid(core_io_weight_in_1_valid),
    .io_weight_in_1_bits(core_io_weight_in_1_bits),
    .io_weight_in_2_ready(core_io_weight_in_2_ready),
    .io_weight_in_2_valid(core_io_weight_in_2_valid),
    .io_weight_in_2_bits(core_io_weight_in_2_bits),
    .io_weight_in_3_ready(core_io_weight_in_3_ready),
    .io_weight_in_3_valid(core_io_weight_in_3_valid),
    .io_weight_in_3_bits(core_io_weight_in_3_bits),
    .io_weight_in_4_ready(core_io_weight_in_4_ready),
    .io_weight_in_4_valid(core_io_weight_in_4_valid),
    .io_weight_in_4_bits(core_io_weight_in_4_bits),
    .io_weight_in_5_ready(core_io_weight_in_5_ready),
    .io_weight_in_5_valid(core_io_weight_in_5_valid),
    .io_weight_in_5_bits(core_io_weight_in_5_bits),
    .io_weight_in_6_ready(core_io_weight_in_6_ready),
    .io_weight_in_6_valid(core_io_weight_in_6_valid),
    .io_weight_in_6_bits(core_io_weight_in_6_bits),
    .io_weight_in_7_ready(core_io_weight_in_7_ready),
    .io_weight_in_7_valid(core_io_weight_in_7_valid),
    .io_weight_in_7_bits(core_io_weight_in_7_bits),
    .io_weight_in_8_ready(core_io_weight_in_8_ready),
    .io_weight_in_8_valid(core_io_weight_in_8_valid),
    .io_weight_in_8_bits(core_io_weight_in_8_bits),
    .io_weight_in_9_ready(core_io_weight_in_9_ready),
    .io_weight_in_9_valid(core_io_weight_in_9_valid),
    .io_weight_in_9_bits(core_io_weight_in_9_bits),
    .io_weight_in_10_ready(core_io_weight_in_10_ready),
    .io_weight_in_10_valid(core_io_weight_in_10_valid),
    .io_weight_in_10_bits(core_io_weight_in_10_bits),
    .io_weight_in_11_ready(core_io_weight_in_11_ready),
    .io_weight_in_11_valid(core_io_weight_in_11_valid),
    .io_weight_in_11_bits(core_io_weight_in_11_bits),
    .io_weight_in_12_ready(core_io_weight_in_12_ready),
    .io_weight_in_12_valid(core_io_weight_in_12_valid),
    .io_weight_in_12_bits(core_io_weight_in_12_bits),
    .io_weight_in_13_ready(core_io_weight_in_13_ready),
    .io_weight_in_13_valid(core_io_weight_in_13_valid),
    .io_weight_in_13_bits(core_io_weight_in_13_bits),
    .io_weight_in_14_ready(core_io_weight_in_14_ready),
    .io_weight_in_14_valid(core_io_weight_in_14_valid),
    .io_weight_in_14_bits(core_io_weight_in_14_bits),
    .io_weight_in_15_ready(core_io_weight_in_15_ready),
    .io_weight_in_15_valid(core_io_weight_in_15_valid),
    .io_weight_in_15_bits(core_io_weight_in_15_bits),
    .io_value_in_0_ready(core_io_value_in_0_ready),
    .io_value_in_0_valid(core_io_value_in_0_valid),
    .io_value_in_0_bits(core_io_value_in_0_bits),
    .io_value_in_1_ready(core_io_value_in_1_ready),
    .io_value_in_1_valid(core_io_value_in_1_valid),
    .io_value_in_1_bits(core_io_value_in_1_bits),
    .io_value_in_2_ready(core_io_value_in_2_ready),
    .io_value_in_2_valid(core_io_value_in_2_valid),
    .io_value_in_2_bits(core_io_value_in_2_bits),
    .io_value_in_3_ready(core_io_value_in_3_ready),
    .io_value_in_3_valid(core_io_value_in_3_valid),
    .io_value_in_3_bits(core_io_value_in_3_bits),
    .io_value_in_4_ready(core_io_value_in_4_ready),
    .io_value_in_4_valid(core_io_value_in_4_valid),
    .io_value_in_4_bits(core_io_value_in_4_bits),
    .io_value_in_5_ready(core_io_value_in_5_ready),
    .io_value_in_5_valid(core_io_value_in_5_valid),
    .io_value_in_5_bits(core_io_value_in_5_bits),
    .io_value_in_6_ready(core_io_value_in_6_ready),
    .io_value_in_6_valid(core_io_value_in_6_valid),
    .io_value_in_6_bits(core_io_value_in_6_bits),
    .io_value_in_7_ready(core_io_value_in_7_ready),
    .io_value_in_7_valid(core_io_value_in_7_valid),
    .io_value_in_7_bits(core_io_value_in_7_bits),
    .io_value_in_8_ready(core_io_value_in_8_ready),
    .io_value_in_8_valid(core_io_value_in_8_valid),
    .io_value_in_8_bits(core_io_value_in_8_bits),
    .io_value_in_9_ready(core_io_value_in_9_ready),
    .io_value_in_9_valid(core_io_value_in_9_valid),
    .io_value_in_9_bits(core_io_value_in_9_bits),
    .io_value_in_10_ready(core_io_value_in_10_ready),
    .io_value_in_10_valid(core_io_value_in_10_valid),
    .io_value_in_10_bits(core_io_value_in_10_bits),
    .io_value_in_11_ready(core_io_value_in_11_ready),
    .io_value_in_11_valid(core_io_value_in_11_valid),
    .io_value_in_11_bits(core_io_value_in_11_bits),
    .io_value_in_12_ready(core_io_value_in_12_ready),
    .io_value_in_12_valid(core_io_value_in_12_valid),
    .io_value_in_12_bits(core_io_value_in_12_bits),
    .io_value_in_13_ready(core_io_value_in_13_ready),
    .io_value_in_13_valid(core_io_value_in_13_valid),
    .io_value_in_13_bits(core_io_value_in_13_bits),
    .io_value_in_14_ready(core_io_value_in_14_ready),
    .io_value_in_14_valid(core_io_value_in_14_valid),
    .io_value_in_14_bits(core_io_value_in_14_bits),
    .io_value_in_15_ready(core_io_value_in_15_ready),
    .io_value_in_15_valid(core_io_value_in_15_valid),
    .io_value_in_15_bits(core_io_value_in_15_bits),
    .io_value_out_0_0_ready(core_io_value_out_0_0_ready),
    .io_value_out_0_0_valid(core_io_value_out_0_0_valid),
    .io_value_out_0_0_bits(core_io_value_out_0_0_bits),
    .io_value_out_0_1_ready(core_io_value_out_0_1_ready),
    .io_value_out_0_1_valid(core_io_value_out_0_1_valid),
    .io_value_out_0_1_bits(core_io_value_out_0_1_bits),
    .io_value_out_0_2_ready(core_io_value_out_0_2_ready),
    .io_value_out_0_2_valid(core_io_value_out_0_2_valid),
    .io_value_out_0_2_bits(core_io_value_out_0_2_bits),
    .io_value_out_0_3_ready(core_io_value_out_0_3_ready),
    .io_value_out_0_3_valid(core_io_value_out_0_3_valid),
    .io_value_out_0_3_bits(core_io_value_out_0_3_bits),
    .io_value_out_0_4_ready(core_io_value_out_0_4_ready),
    .io_value_out_0_4_valid(core_io_value_out_0_4_valid),
    .io_value_out_0_4_bits(core_io_value_out_0_4_bits),
    .io_value_out_0_5_ready(core_io_value_out_0_5_ready),
    .io_value_out_0_5_valid(core_io_value_out_0_5_valid),
    .io_value_out_0_5_bits(core_io_value_out_0_5_bits),
    .io_value_out_0_6_ready(core_io_value_out_0_6_ready),
    .io_value_out_0_6_valid(core_io_value_out_0_6_valid),
    .io_value_out_0_6_bits(core_io_value_out_0_6_bits),
    .io_value_out_0_7_ready(core_io_value_out_0_7_ready),
    .io_value_out_0_7_valid(core_io_value_out_0_7_valid),
    .io_value_out_0_7_bits(core_io_value_out_0_7_bits),
    .io_value_out_0_8_ready(core_io_value_out_0_8_ready),
    .io_value_out_0_8_valid(core_io_value_out_0_8_valid),
    .io_value_out_0_8_bits(core_io_value_out_0_8_bits),
    .io_value_out_0_9_ready(core_io_value_out_0_9_ready),
    .io_value_out_0_9_valid(core_io_value_out_0_9_valid),
    .io_value_out_0_9_bits(core_io_value_out_0_9_bits),
    .io_value_out_0_10_ready(core_io_value_out_0_10_ready),
    .io_value_out_0_10_valid(core_io_value_out_0_10_valid),
    .io_value_out_0_10_bits(core_io_value_out_0_10_bits),
    .io_value_out_0_11_ready(core_io_value_out_0_11_ready),
    .io_value_out_0_11_valid(core_io_value_out_0_11_valid),
    .io_value_out_0_11_bits(core_io_value_out_0_11_bits),
    .io_value_out_0_12_ready(core_io_value_out_0_12_ready),
    .io_value_out_0_12_valid(core_io_value_out_0_12_valid),
    .io_value_out_0_12_bits(core_io_value_out_0_12_bits),
    .io_value_out_0_13_ready(core_io_value_out_0_13_ready),
    .io_value_out_0_13_valid(core_io_value_out_0_13_valid),
    .io_value_out_0_13_bits(core_io_value_out_0_13_bits),
    .io_value_out_0_14_ready(core_io_value_out_0_14_ready),
    .io_value_out_0_14_valid(core_io_value_out_0_14_valid),
    .io_value_out_0_14_bits(core_io_value_out_0_14_bits),
    .io_value_out_0_15_ready(core_io_value_out_0_15_ready),
    .io_value_out_0_15_valid(core_io_value_out_0_15_valid),
    .io_value_out_0_15_bits(core_io_value_out_0_15_bits),
    .io_value_out_1_0_ready(core_io_value_out_1_0_ready),
    .io_value_out_1_0_valid(core_io_value_out_1_0_valid),
    .io_value_out_1_0_bits(core_io_value_out_1_0_bits),
    .io_value_out_1_1_ready(core_io_value_out_1_1_ready),
    .io_value_out_1_1_valid(core_io_value_out_1_1_valid),
    .io_value_out_1_1_bits(core_io_value_out_1_1_bits),
    .io_value_out_1_2_ready(core_io_value_out_1_2_ready),
    .io_value_out_1_2_valid(core_io_value_out_1_2_valid),
    .io_value_out_1_2_bits(core_io_value_out_1_2_bits),
    .io_value_out_1_3_ready(core_io_value_out_1_3_ready),
    .io_value_out_1_3_valid(core_io_value_out_1_3_valid),
    .io_value_out_1_3_bits(core_io_value_out_1_3_bits),
    .io_value_out_1_4_ready(core_io_value_out_1_4_ready),
    .io_value_out_1_4_valid(core_io_value_out_1_4_valid),
    .io_value_out_1_4_bits(core_io_value_out_1_4_bits),
    .io_value_out_1_5_ready(core_io_value_out_1_5_ready),
    .io_value_out_1_5_valid(core_io_value_out_1_5_valid),
    .io_value_out_1_5_bits(core_io_value_out_1_5_bits),
    .io_value_out_1_6_ready(core_io_value_out_1_6_ready),
    .io_value_out_1_6_valid(core_io_value_out_1_6_valid),
    .io_value_out_1_6_bits(core_io_value_out_1_6_bits),
    .io_value_out_1_7_ready(core_io_value_out_1_7_ready),
    .io_value_out_1_7_valid(core_io_value_out_1_7_valid),
    .io_value_out_1_7_bits(core_io_value_out_1_7_bits),
    .io_value_out_1_8_ready(core_io_value_out_1_8_ready),
    .io_value_out_1_8_valid(core_io_value_out_1_8_valid),
    .io_value_out_1_8_bits(core_io_value_out_1_8_bits),
    .io_value_out_1_9_ready(core_io_value_out_1_9_ready),
    .io_value_out_1_9_valid(core_io_value_out_1_9_valid),
    .io_value_out_1_9_bits(core_io_value_out_1_9_bits),
    .io_value_out_1_10_ready(core_io_value_out_1_10_ready),
    .io_value_out_1_10_valid(core_io_value_out_1_10_valid),
    .io_value_out_1_10_bits(core_io_value_out_1_10_bits),
    .io_value_out_1_11_ready(core_io_value_out_1_11_ready),
    .io_value_out_1_11_valid(core_io_value_out_1_11_valid),
    .io_value_out_1_11_bits(core_io_value_out_1_11_bits),
    .io_value_out_1_12_ready(core_io_value_out_1_12_ready),
    .io_value_out_1_12_valid(core_io_value_out_1_12_valid),
    .io_value_out_1_12_bits(core_io_value_out_1_12_bits),
    .io_value_out_1_13_ready(core_io_value_out_1_13_ready),
    .io_value_out_1_13_valid(core_io_value_out_1_13_valid),
    .io_value_out_1_13_bits(core_io_value_out_1_13_bits),
    .io_value_out_1_14_ready(core_io_value_out_1_14_ready),
    .io_value_out_1_14_valid(core_io_value_out_1_14_valid),
    .io_value_out_1_14_bits(core_io_value_out_1_14_bits),
    .io_value_out_1_15_ready(core_io_value_out_1_15_ready),
    .io_value_out_1_15_valid(core_io_value_out_1_15_valid),
    .io_value_out_1_15_bits(core_io_value_out_1_15_bits),
    .io_value_out_2_0_ready(core_io_value_out_2_0_ready),
    .io_value_out_2_0_valid(core_io_value_out_2_0_valid),
    .io_value_out_2_0_bits(core_io_value_out_2_0_bits),
    .io_value_out_2_1_ready(core_io_value_out_2_1_ready),
    .io_value_out_2_1_valid(core_io_value_out_2_1_valid),
    .io_value_out_2_1_bits(core_io_value_out_2_1_bits),
    .io_value_out_2_2_ready(core_io_value_out_2_2_ready),
    .io_value_out_2_2_valid(core_io_value_out_2_2_valid),
    .io_value_out_2_2_bits(core_io_value_out_2_2_bits),
    .io_value_out_2_3_ready(core_io_value_out_2_3_ready),
    .io_value_out_2_3_valid(core_io_value_out_2_3_valid),
    .io_value_out_2_3_bits(core_io_value_out_2_3_bits),
    .io_value_out_2_4_ready(core_io_value_out_2_4_ready),
    .io_value_out_2_4_valid(core_io_value_out_2_4_valid),
    .io_value_out_2_4_bits(core_io_value_out_2_4_bits),
    .io_value_out_2_5_ready(core_io_value_out_2_5_ready),
    .io_value_out_2_5_valid(core_io_value_out_2_5_valid),
    .io_value_out_2_5_bits(core_io_value_out_2_5_bits),
    .io_value_out_2_6_ready(core_io_value_out_2_6_ready),
    .io_value_out_2_6_valid(core_io_value_out_2_6_valid),
    .io_value_out_2_6_bits(core_io_value_out_2_6_bits),
    .io_value_out_2_7_ready(core_io_value_out_2_7_ready),
    .io_value_out_2_7_valid(core_io_value_out_2_7_valid),
    .io_value_out_2_7_bits(core_io_value_out_2_7_bits),
    .io_value_out_2_8_ready(core_io_value_out_2_8_ready),
    .io_value_out_2_8_valid(core_io_value_out_2_8_valid),
    .io_value_out_2_8_bits(core_io_value_out_2_8_bits),
    .io_value_out_2_9_ready(core_io_value_out_2_9_ready),
    .io_value_out_2_9_valid(core_io_value_out_2_9_valid),
    .io_value_out_2_9_bits(core_io_value_out_2_9_bits),
    .io_value_out_2_10_ready(core_io_value_out_2_10_ready),
    .io_value_out_2_10_valid(core_io_value_out_2_10_valid),
    .io_value_out_2_10_bits(core_io_value_out_2_10_bits),
    .io_value_out_2_11_ready(core_io_value_out_2_11_ready),
    .io_value_out_2_11_valid(core_io_value_out_2_11_valid),
    .io_value_out_2_11_bits(core_io_value_out_2_11_bits),
    .io_value_out_2_12_ready(core_io_value_out_2_12_ready),
    .io_value_out_2_12_valid(core_io_value_out_2_12_valid),
    .io_value_out_2_12_bits(core_io_value_out_2_12_bits),
    .io_value_out_2_13_ready(core_io_value_out_2_13_ready),
    .io_value_out_2_13_valid(core_io_value_out_2_13_valid),
    .io_value_out_2_13_bits(core_io_value_out_2_13_bits),
    .io_value_out_2_14_ready(core_io_value_out_2_14_ready),
    .io_value_out_2_14_valid(core_io_value_out_2_14_valid),
    .io_value_out_2_14_bits(core_io_value_out_2_14_bits),
    .io_value_out_2_15_ready(core_io_value_out_2_15_ready),
    .io_value_out_2_15_valid(core_io_value_out_2_15_valid),
    .io_value_out_2_15_bits(core_io_value_out_2_15_bits),
    .io_value_out_3_0_ready(core_io_value_out_3_0_ready),
    .io_value_out_3_0_valid(core_io_value_out_3_0_valid),
    .io_value_out_3_0_bits(core_io_value_out_3_0_bits),
    .io_value_out_3_1_ready(core_io_value_out_3_1_ready),
    .io_value_out_3_1_valid(core_io_value_out_3_1_valid),
    .io_value_out_3_1_bits(core_io_value_out_3_1_bits),
    .io_value_out_3_2_ready(core_io_value_out_3_2_ready),
    .io_value_out_3_2_valid(core_io_value_out_3_2_valid),
    .io_value_out_3_2_bits(core_io_value_out_3_2_bits),
    .io_value_out_3_3_ready(core_io_value_out_3_3_ready),
    .io_value_out_3_3_valid(core_io_value_out_3_3_valid),
    .io_value_out_3_3_bits(core_io_value_out_3_3_bits),
    .io_value_out_3_4_ready(core_io_value_out_3_4_ready),
    .io_value_out_3_4_valid(core_io_value_out_3_4_valid),
    .io_value_out_3_4_bits(core_io_value_out_3_4_bits),
    .io_value_out_3_5_ready(core_io_value_out_3_5_ready),
    .io_value_out_3_5_valid(core_io_value_out_3_5_valid),
    .io_value_out_3_5_bits(core_io_value_out_3_5_bits),
    .io_value_out_3_6_ready(core_io_value_out_3_6_ready),
    .io_value_out_3_6_valid(core_io_value_out_3_6_valid),
    .io_value_out_3_6_bits(core_io_value_out_3_6_bits),
    .io_value_out_3_7_ready(core_io_value_out_3_7_ready),
    .io_value_out_3_7_valid(core_io_value_out_3_7_valid),
    .io_value_out_3_7_bits(core_io_value_out_3_7_bits),
    .io_value_out_3_8_ready(core_io_value_out_3_8_ready),
    .io_value_out_3_8_valid(core_io_value_out_3_8_valid),
    .io_value_out_3_8_bits(core_io_value_out_3_8_bits),
    .io_value_out_3_9_ready(core_io_value_out_3_9_ready),
    .io_value_out_3_9_valid(core_io_value_out_3_9_valid),
    .io_value_out_3_9_bits(core_io_value_out_3_9_bits),
    .io_value_out_3_10_ready(core_io_value_out_3_10_ready),
    .io_value_out_3_10_valid(core_io_value_out_3_10_valid),
    .io_value_out_3_10_bits(core_io_value_out_3_10_bits),
    .io_value_out_3_11_ready(core_io_value_out_3_11_ready),
    .io_value_out_3_11_valid(core_io_value_out_3_11_valid),
    .io_value_out_3_11_bits(core_io_value_out_3_11_bits),
    .io_value_out_3_12_ready(core_io_value_out_3_12_ready),
    .io_value_out_3_12_valid(core_io_value_out_3_12_valid),
    .io_value_out_3_12_bits(core_io_value_out_3_12_bits),
    .io_value_out_3_13_ready(core_io_value_out_3_13_ready),
    .io_value_out_3_13_valid(core_io_value_out_3_13_valid),
    .io_value_out_3_13_bits(core_io_value_out_3_13_bits),
    .io_value_out_3_14_ready(core_io_value_out_3_14_ready),
    .io_value_out_3_14_valid(core_io_value_out_3_14_valid),
    .io_value_out_3_14_bits(core_io_value_out_3_14_bits),
    .io_value_out_3_15_ready(core_io_value_out_3_15_ready),
    .io_value_out_3_15_valid(core_io_value_out_3_15_valid),
    .io_value_out_3_15_bits(core_io_value_out_3_15_bits),
    .io_value_out_4_0_ready(core_io_value_out_4_0_ready),
    .io_value_out_4_0_valid(core_io_value_out_4_0_valid),
    .io_value_out_4_0_bits(core_io_value_out_4_0_bits),
    .io_value_out_4_1_ready(core_io_value_out_4_1_ready),
    .io_value_out_4_1_valid(core_io_value_out_4_1_valid),
    .io_value_out_4_1_bits(core_io_value_out_4_1_bits),
    .io_value_out_4_2_ready(core_io_value_out_4_2_ready),
    .io_value_out_4_2_valid(core_io_value_out_4_2_valid),
    .io_value_out_4_2_bits(core_io_value_out_4_2_bits),
    .io_value_out_4_3_ready(core_io_value_out_4_3_ready),
    .io_value_out_4_3_valid(core_io_value_out_4_3_valid),
    .io_value_out_4_3_bits(core_io_value_out_4_3_bits),
    .io_value_out_4_4_ready(core_io_value_out_4_4_ready),
    .io_value_out_4_4_valid(core_io_value_out_4_4_valid),
    .io_value_out_4_4_bits(core_io_value_out_4_4_bits),
    .io_value_out_4_5_ready(core_io_value_out_4_5_ready),
    .io_value_out_4_5_valid(core_io_value_out_4_5_valid),
    .io_value_out_4_5_bits(core_io_value_out_4_5_bits),
    .io_value_out_4_6_ready(core_io_value_out_4_6_ready),
    .io_value_out_4_6_valid(core_io_value_out_4_6_valid),
    .io_value_out_4_6_bits(core_io_value_out_4_6_bits),
    .io_value_out_4_7_ready(core_io_value_out_4_7_ready),
    .io_value_out_4_7_valid(core_io_value_out_4_7_valid),
    .io_value_out_4_7_bits(core_io_value_out_4_7_bits),
    .io_value_out_4_8_ready(core_io_value_out_4_8_ready),
    .io_value_out_4_8_valid(core_io_value_out_4_8_valid),
    .io_value_out_4_8_bits(core_io_value_out_4_8_bits),
    .io_value_out_4_9_ready(core_io_value_out_4_9_ready),
    .io_value_out_4_9_valid(core_io_value_out_4_9_valid),
    .io_value_out_4_9_bits(core_io_value_out_4_9_bits),
    .io_value_out_4_10_ready(core_io_value_out_4_10_ready),
    .io_value_out_4_10_valid(core_io_value_out_4_10_valid),
    .io_value_out_4_10_bits(core_io_value_out_4_10_bits),
    .io_value_out_4_11_ready(core_io_value_out_4_11_ready),
    .io_value_out_4_11_valid(core_io_value_out_4_11_valid),
    .io_value_out_4_11_bits(core_io_value_out_4_11_bits),
    .io_value_out_4_12_ready(core_io_value_out_4_12_ready),
    .io_value_out_4_12_valid(core_io_value_out_4_12_valid),
    .io_value_out_4_12_bits(core_io_value_out_4_12_bits),
    .io_value_out_4_13_ready(core_io_value_out_4_13_ready),
    .io_value_out_4_13_valid(core_io_value_out_4_13_valid),
    .io_value_out_4_13_bits(core_io_value_out_4_13_bits),
    .io_value_out_4_14_ready(core_io_value_out_4_14_ready),
    .io_value_out_4_14_valid(core_io_value_out_4_14_valid),
    .io_value_out_4_14_bits(core_io_value_out_4_14_bits),
    .io_value_out_4_15_ready(core_io_value_out_4_15_ready),
    .io_value_out_4_15_valid(core_io_value_out_4_15_valid),
    .io_value_out_4_15_bits(core_io_value_out_4_15_bits),
    .io_value_out_5_0_ready(core_io_value_out_5_0_ready),
    .io_value_out_5_0_valid(core_io_value_out_5_0_valid),
    .io_value_out_5_0_bits(core_io_value_out_5_0_bits),
    .io_value_out_5_1_ready(core_io_value_out_5_1_ready),
    .io_value_out_5_1_valid(core_io_value_out_5_1_valid),
    .io_value_out_5_1_bits(core_io_value_out_5_1_bits),
    .io_value_out_5_2_ready(core_io_value_out_5_2_ready),
    .io_value_out_5_2_valid(core_io_value_out_5_2_valid),
    .io_value_out_5_2_bits(core_io_value_out_5_2_bits),
    .io_value_out_5_3_ready(core_io_value_out_5_3_ready),
    .io_value_out_5_3_valid(core_io_value_out_5_3_valid),
    .io_value_out_5_3_bits(core_io_value_out_5_3_bits),
    .io_value_out_5_4_ready(core_io_value_out_5_4_ready),
    .io_value_out_5_4_valid(core_io_value_out_5_4_valid),
    .io_value_out_5_4_bits(core_io_value_out_5_4_bits),
    .io_value_out_5_5_ready(core_io_value_out_5_5_ready),
    .io_value_out_5_5_valid(core_io_value_out_5_5_valid),
    .io_value_out_5_5_bits(core_io_value_out_5_5_bits),
    .io_value_out_5_6_ready(core_io_value_out_5_6_ready),
    .io_value_out_5_6_valid(core_io_value_out_5_6_valid),
    .io_value_out_5_6_bits(core_io_value_out_5_6_bits),
    .io_value_out_5_7_ready(core_io_value_out_5_7_ready),
    .io_value_out_5_7_valid(core_io_value_out_5_7_valid),
    .io_value_out_5_7_bits(core_io_value_out_5_7_bits),
    .io_value_out_5_8_ready(core_io_value_out_5_8_ready),
    .io_value_out_5_8_valid(core_io_value_out_5_8_valid),
    .io_value_out_5_8_bits(core_io_value_out_5_8_bits),
    .io_value_out_5_9_ready(core_io_value_out_5_9_ready),
    .io_value_out_5_9_valid(core_io_value_out_5_9_valid),
    .io_value_out_5_9_bits(core_io_value_out_5_9_bits),
    .io_value_out_5_10_ready(core_io_value_out_5_10_ready),
    .io_value_out_5_10_valid(core_io_value_out_5_10_valid),
    .io_value_out_5_10_bits(core_io_value_out_5_10_bits),
    .io_value_out_5_11_ready(core_io_value_out_5_11_ready),
    .io_value_out_5_11_valid(core_io_value_out_5_11_valid),
    .io_value_out_5_11_bits(core_io_value_out_5_11_bits),
    .io_value_out_5_12_ready(core_io_value_out_5_12_ready),
    .io_value_out_5_12_valid(core_io_value_out_5_12_valid),
    .io_value_out_5_12_bits(core_io_value_out_5_12_bits),
    .io_value_out_5_13_ready(core_io_value_out_5_13_ready),
    .io_value_out_5_13_valid(core_io_value_out_5_13_valid),
    .io_value_out_5_13_bits(core_io_value_out_5_13_bits),
    .io_value_out_5_14_ready(core_io_value_out_5_14_ready),
    .io_value_out_5_14_valid(core_io_value_out_5_14_valid),
    .io_value_out_5_14_bits(core_io_value_out_5_14_bits),
    .io_value_out_5_15_ready(core_io_value_out_5_15_ready),
    .io_value_out_5_15_valid(core_io_value_out_5_15_valid),
    .io_value_out_5_15_bits(core_io_value_out_5_15_bits),
    .io_value_out_6_0_ready(core_io_value_out_6_0_ready),
    .io_value_out_6_0_valid(core_io_value_out_6_0_valid),
    .io_value_out_6_0_bits(core_io_value_out_6_0_bits),
    .io_value_out_6_1_ready(core_io_value_out_6_1_ready),
    .io_value_out_6_1_valid(core_io_value_out_6_1_valid),
    .io_value_out_6_1_bits(core_io_value_out_6_1_bits),
    .io_value_out_6_2_ready(core_io_value_out_6_2_ready),
    .io_value_out_6_2_valid(core_io_value_out_6_2_valid),
    .io_value_out_6_2_bits(core_io_value_out_6_2_bits),
    .io_value_out_6_3_ready(core_io_value_out_6_3_ready),
    .io_value_out_6_3_valid(core_io_value_out_6_3_valid),
    .io_value_out_6_3_bits(core_io_value_out_6_3_bits),
    .io_value_out_6_4_ready(core_io_value_out_6_4_ready),
    .io_value_out_6_4_valid(core_io_value_out_6_4_valid),
    .io_value_out_6_4_bits(core_io_value_out_6_4_bits),
    .io_value_out_6_5_ready(core_io_value_out_6_5_ready),
    .io_value_out_6_5_valid(core_io_value_out_6_5_valid),
    .io_value_out_6_5_bits(core_io_value_out_6_5_bits),
    .io_value_out_6_6_ready(core_io_value_out_6_6_ready),
    .io_value_out_6_6_valid(core_io_value_out_6_6_valid),
    .io_value_out_6_6_bits(core_io_value_out_6_6_bits),
    .io_value_out_6_7_ready(core_io_value_out_6_7_ready),
    .io_value_out_6_7_valid(core_io_value_out_6_7_valid),
    .io_value_out_6_7_bits(core_io_value_out_6_7_bits),
    .io_value_out_6_8_ready(core_io_value_out_6_8_ready),
    .io_value_out_6_8_valid(core_io_value_out_6_8_valid),
    .io_value_out_6_8_bits(core_io_value_out_6_8_bits),
    .io_value_out_6_9_ready(core_io_value_out_6_9_ready),
    .io_value_out_6_9_valid(core_io_value_out_6_9_valid),
    .io_value_out_6_9_bits(core_io_value_out_6_9_bits),
    .io_value_out_6_10_ready(core_io_value_out_6_10_ready),
    .io_value_out_6_10_valid(core_io_value_out_6_10_valid),
    .io_value_out_6_10_bits(core_io_value_out_6_10_bits),
    .io_value_out_6_11_ready(core_io_value_out_6_11_ready),
    .io_value_out_6_11_valid(core_io_value_out_6_11_valid),
    .io_value_out_6_11_bits(core_io_value_out_6_11_bits),
    .io_value_out_6_12_ready(core_io_value_out_6_12_ready),
    .io_value_out_6_12_valid(core_io_value_out_6_12_valid),
    .io_value_out_6_12_bits(core_io_value_out_6_12_bits),
    .io_value_out_6_13_ready(core_io_value_out_6_13_ready),
    .io_value_out_6_13_valid(core_io_value_out_6_13_valid),
    .io_value_out_6_13_bits(core_io_value_out_6_13_bits),
    .io_value_out_6_14_ready(core_io_value_out_6_14_ready),
    .io_value_out_6_14_valid(core_io_value_out_6_14_valid),
    .io_value_out_6_14_bits(core_io_value_out_6_14_bits),
    .io_value_out_6_15_ready(core_io_value_out_6_15_ready),
    .io_value_out_6_15_valid(core_io_value_out_6_15_valid),
    .io_value_out_6_15_bits(core_io_value_out_6_15_bits),
    .io_value_out_7_0_ready(core_io_value_out_7_0_ready),
    .io_value_out_7_0_valid(core_io_value_out_7_0_valid),
    .io_value_out_7_0_bits(core_io_value_out_7_0_bits),
    .io_value_out_7_1_ready(core_io_value_out_7_1_ready),
    .io_value_out_7_1_valid(core_io_value_out_7_1_valid),
    .io_value_out_7_1_bits(core_io_value_out_7_1_bits),
    .io_value_out_7_2_ready(core_io_value_out_7_2_ready),
    .io_value_out_7_2_valid(core_io_value_out_7_2_valid),
    .io_value_out_7_2_bits(core_io_value_out_7_2_bits),
    .io_value_out_7_3_ready(core_io_value_out_7_3_ready),
    .io_value_out_7_3_valid(core_io_value_out_7_3_valid),
    .io_value_out_7_3_bits(core_io_value_out_7_3_bits),
    .io_value_out_7_4_ready(core_io_value_out_7_4_ready),
    .io_value_out_7_4_valid(core_io_value_out_7_4_valid),
    .io_value_out_7_4_bits(core_io_value_out_7_4_bits),
    .io_value_out_7_5_ready(core_io_value_out_7_5_ready),
    .io_value_out_7_5_valid(core_io_value_out_7_5_valid),
    .io_value_out_7_5_bits(core_io_value_out_7_5_bits),
    .io_value_out_7_6_ready(core_io_value_out_7_6_ready),
    .io_value_out_7_6_valid(core_io_value_out_7_6_valid),
    .io_value_out_7_6_bits(core_io_value_out_7_6_bits),
    .io_value_out_7_7_ready(core_io_value_out_7_7_ready),
    .io_value_out_7_7_valid(core_io_value_out_7_7_valid),
    .io_value_out_7_7_bits(core_io_value_out_7_7_bits),
    .io_value_out_7_8_ready(core_io_value_out_7_8_ready),
    .io_value_out_7_8_valid(core_io_value_out_7_8_valid),
    .io_value_out_7_8_bits(core_io_value_out_7_8_bits),
    .io_value_out_7_9_ready(core_io_value_out_7_9_ready),
    .io_value_out_7_9_valid(core_io_value_out_7_9_valid),
    .io_value_out_7_9_bits(core_io_value_out_7_9_bits),
    .io_value_out_7_10_ready(core_io_value_out_7_10_ready),
    .io_value_out_7_10_valid(core_io_value_out_7_10_valid),
    .io_value_out_7_10_bits(core_io_value_out_7_10_bits),
    .io_value_out_7_11_ready(core_io_value_out_7_11_ready),
    .io_value_out_7_11_valid(core_io_value_out_7_11_valid),
    .io_value_out_7_11_bits(core_io_value_out_7_11_bits),
    .io_value_out_7_12_ready(core_io_value_out_7_12_ready),
    .io_value_out_7_12_valid(core_io_value_out_7_12_valid),
    .io_value_out_7_12_bits(core_io_value_out_7_12_bits),
    .io_value_out_7_13_ready(core_io_value_out_7_13_ready),
    .io_value_out_7_13_valid(core_io_value_out_7_13_valid),
    .io_value_out_7_13_bits(core_io_value_out_7_13_bits),
    .io_value_out_7_14_ready(core_io_value_out_7_14_ready),
    .io_value_out_7_14_valid(core_io_value_out_7_14_valid),
    .io_value_out_7_14_bits(core_io_value_out_7_14_bits),
    .io_value_out_7_15_ready(core_io_value_out_7_15_ready),
    .io_value_out_7_15_valid(core_io_value_out_7_15_valid),
    .io_value_out_7_15_bits(core_io_value_out_7_15_bits),
    .io_value_out_8_0_ready(core_io_value_out_8_0_ready),
    .io_value_out_8_0_valid(core_io_value_out_8_0_valid),
    .io_value_out_8_0_bits(core_io_value_out_8_0_bits),
    .io_value_out_8_1_ready(core_io_value_out_8_1_ready),
    .io_value_out_8_1_valid(core_io_value_out_8_1_valid),
    .io_value_out_8_1_bits(core_io_value_out_8_1_bits),
    .io_value_out_8_2_ready(core_io_value_out_8_2_ready),
    .io_value_out_8_2_valid(core_io_value_out_8_2_valid),
    .io_value_out_8_2_bits(core_io_value_out_8_2_bits),
    .io_value_out_8_3_ready(core_io_value_out_8_3_ready),
    .io_value_out_8_3_valid(core_io_value_out_8_3_valid),
    .io_value_out_8_3_bits(core_io_value_out_8_3_bits),
    .io_value_out_8_4_ready(core_io_value_out_8_4_ready),
    .io_value_out_8_4_valid(core_io_value_out_8_4_valid),
    .io_value_out_8_4_bits(core_io_value_out_8_4_bits),
    .io_value_out_8_5_ready(core_io_value_out_8_5_ready),
    .io_value_out_8_5_valid(core_io_value_out_8_5_valid),
    .io_value_out_8_5_bits(core_io_value_out_8_5_bits),
    .io_value_out_8_6_ready(core_io_value_out_8_6_ready),
    .io_value_out_8_6_valid(core_io_value_out_8_6_valid),
    .io_value_out_8_6_bits(core_io_value_out_8_6_bits),
    .io_value_out_8_7_ready(core_io_value_out_8_7_ready),
    .io_value_out_8_7_valid(core_io_value_out_8_7_valid),
    .io_value_out_8_7_bits(core_io_value_out_8_7_bits),
    .io_value_out_8_8_ready(core_io_value_out_8_8_ready),
    .io_value_out_8_8_valid(core_io_value_out_8_8_valid),
    .io_value_out_8_8_bits(core_io_value_out_8_8_bits),
    .io_value_out_8_9_ready(core_io_value_out_8_9_ready),
    .io_value_out_8_9_valid(core_io_value_out_8_9_valid),
    .io_value_out_8_9_bits(core_io_value_out_8_9_bits),
    .io_value_out_8_10_ready(core_io_value_out_8_10_ready),
    .io_value_out_8_10_valid(core_io_value_out_8_10_valid),
    .io_value_out_8_10_bits(core_io_value_out_8_10_bits),
    .io_value_out_8_11_ready(core_io_value_out_8_11_ready),
    .io_value_out_8_11_valid(core_io_value_out_8_11_valid),
    .io_value_out_8_11_bits(core_io_value_out_8_11_bits),
    .io_value_out_8_12_ready(core_io_value_out_8_12_ready),
    .io_value_out_8_12_valid(core_io_value_out_8_12_valid),
    .io_value_out_8_12_bits(core_io_value_out_8_12_bits),
    .io_value_out_8_13_ready(core_io_value_out_8_13_ready),
    .io_value_out_8_13_valid(core_io_value_out_8_13_valid),
    .io_value_out_8_13_bits(core_io_value_out_8_13_bits),
    .io_value_out_8_14_ready(core_io_value_out_8_14_ready),
    .io_value_out_8_14_valid(core_io_value_out_8_14_valid),
    .io_value_out_8_14_bits(core_io_value_out_8_14_bits),
    .io_value_out_8_15_ready(core_io_value_out_8_15_ready),
    .io_value_out_8_15_valid(core_io_value_out_8_15_valid),
    .io_value_out_8_15_bits(core_io_value_out_8_15_bits),
    .io_value_out_9_0_ready(core_io_value_out_9_0_ready),
    .io_value_out_9_0_valid(core_io_value_out_9_0_valid),
    .io_value_out_9_0_bits(core_io_value_out_9_0_bits),
    .io_value_out_9_1_ready(core_io_value_out_9_1_ready),
    .io_value_out_9_1_valid(core_io_value_out_9_1_valid),
    .io_value_out_9_1_bits(core_io_value_out_9_1_bits),
    .io_value_out_9_2_ready(core_io_value_out_9_2_ready),
    .io_value_out_9_2_valid(core_io_value_out_9_2_valid),
    .io_value_out_9_2_bits(core_io_value_out_9_2_bits),
    .io_value_out_9_3_ready(core_io_value_out_9_3_ready),
    .io_value_out_9_3_valid(core_io_value_out_9_3_valid),
    .io_value_out_9_3_bits(core_io_value_out_9_3_bits),
    .io_value_out_9_4_ready(core_io_value_out_9_4_ready),
    .io_value_out_9_4_valid(core_io_value_out_9_4_valid),
    .io_value_out_9_4_bits(core_io_value_out_9_4_bits),
    .io_value_out_9_5_ready(core_io_value_out_9_5_ready),
    .io_value_out_9_5_valid(core_io_value_out_9_5_valid),
    .io_value_out_9_5_bits(core_io_value_out_9_5_bits),
    .io_value_out_9_6_ready(core_io_value_out_9_6_ready),
    .io_value_out_9_6_valid(core_io_value_out_9_6_valid),
    .io_value_out_9_6_bits(core_io_value_out_9_6_bits),
    .io_value_out_9_7_ready(core_io_value_out_9_7_ready),
    .io_value_out_9_7_valid(core_io_value_out_9_7_valid),
    .io_value_out_9_7_bits(core_io_value_out_9_7_bits),
    .io_value_out_9_8_ready(core_io_value_out_9_8_ready),
    .io_value_out_9_8_valid(core_io_value_out_9_8_valid),
    .io_value_out_9_8_bits(core_io_value_out_9_8_bits),
    .io_value_out_9_9_ready(core_io_value_out_9_9_ready),
    .io_value_out_9_9_valid(core_io_value_out_9_9_valid),
    .io_value_out_9_9_bits(core_io_value_out_9_9_bits),
    .io_value_out_9_10_ready(core_io_value_out_9_10_ready),
    .io_value_out_9_10_valid(core_io_value_out_9_10_valid),
    .io_value_out_9_10_bits(core_io_value_out_9_10_bits),
    .io_value_out_9_11_ready(core_io_value_out_9_11_ready),
    .io_value_out_9_11_valid(core_io_value_out_9_11_valid),
    .io_value_out_9_11_bits(core_io_value_out_9_11_bits),
    .io_value_out_9_12_ready(core_io_value_out_9_12_ready),
    .io_value_out_9_12_valid(core_io_value_out_9_12_valid),
    .io_value_out_9_12_bits(core_io_value_out_9_12_bits),
    .io_value_out_9_13_ready(core_io_value_out_9_13_ready),
    .io_value_out_9_13_valid(core_io_value_out_9_13_valid),
    .io_value_out_9_13_bits(core_io_value_out_9_13_bits),
    .io_value_out_9_14_ready(core_io_value_out_9_14_ready),
    .io_value_out_9_14_valid(core_io_value_out_9_14_valid),
    .io_value_out_9_14_bits(core_io_value_out_9_14_bits),
    .io_value_out_9_15_ready(core_io_value_out_9_15_ready),
    .io_value_out_9_15_valid(core_io_value_out_9_15_valid),
    .io_value_out_9_15_bits(core_io_value_out_9_15_bits),
    .io_value_out_10_0_ready(core_io_value_out_10_0_ready),
    .io_value_out_10_0_valid(core_io_value_out_10_0_valid),
    .io_value_out_10_0_bits(core_io_value_out_10_0_bits),
    .io_value_out_10_1_ready(core_io_value_out_10_1_ready),
    .io_value_out_10_1_valid(core_io_value_out_10_1_valid),
    .io_value_out_10_1_bits(core_io_value_out_10_1_bits),
    .io_value_out_10_2_ready(core_io_value_out_10_2_ready),
    .io_value_out_10_2_valid(core_io_value_out_10_2_valid),
    .io_value_out_10_2_bits(core_io_value_out_10_2_bits),
    .io_value_out_10_3_ready(core_io_value_out_10_3_ready),
    .io_value_out_10_3_valid(core_io_value_out_10_3_valid),
    .io_value_out_10_3_bits(core_io_value_out_10_3_bits),
    .io_value_out_10_4_ready(core_io_value_out_10_4_ready),
    .io_value_out_10_4_valid(core_io_value_out_10_4_valid),
    .io_value_out_10_4_bits(core_io_value_out_10_4_bits),
    .io_value_out_10_5_ready(core_io_value_out_10_5_ready),
    .io_value_out_10_5_valid(core_io_value_out_10_5_valid),
    .io_value_out_10_5_bits(core_io_value_out_10_5_bits),
    .io_value_out_10_6_ready(core_io_value_out_10_6_ready),
    .io_value_out_10_6_valid(core_io_value_out_10_6_valid),
    .io_value_out_10_6_bits(core_io_value_out_10_6_bits),
    .io_value_out_10_7_ready(core_io_value_out_10_7_ready),
    .io_value_out_10_7_valid(core_io_value_out_10_7_valid),
    .io_value_out_10_7_bits(core_io_value_out_10_7_bits),
    .io_value_out_10_8_ready(core_io_value_out_10_8_ready),
    .io_value_out_10_8_valid(core_io_value_out_10_8_valid),
    .io_value_out_10_8_bits(core_io_value_out_10_8_bits),
    .io_value_out_10_9_ready(core_io_value_out_10_9_ready),
    .io_value_out_10_9_valid(core_io_value_out_10_9_valid),
    .io_value_out_10_9_bits(core_io_value_out_10_9_bits),
    .io_value_out_10_10_ready(core_io_value_out_10_10_ready),
    .io_value_out_10_10_valid(core_io_value_out_10_10_valid),
    .io_value_out_10_10_bits(core_io_value_out_10_10_bits),
    .io_value_out_10_11_ready(core_io_value_out_10_11_ready),
    .io_value_out_10_11_valid(core_io_value_out_10_11_valid),
    .io_value_out_10_11_bits(core_io_value_out_10_11_bits),
    .io_value_out_10_12_ready(core_io_value_out_10_12_ready),
    .io_value_out_10_12_valid(core_io_value_out_10_12_valid),
    .io_value_out_10_12_bits(core_io_value_out_10_12_bits),
    .io_value_out_10_13_ready(core_io_value_out_10_13_ready),
    .io_value_out_10_13_valid(core_io_value_out_10_13_valid),
    .io_value_out_10_13_bits(core_io_value_out_10_13_bits),
    .io_value_out_10_14_ready(core_io_value_out_10_14_ready),
    .io_value_out_10_14_valid(core_io_value_out_10_14_valid),
    .io_value_out_10_14_bits(core_io_value_out_10_14_bits),
    .io_value_out_10_15_ready(core_io_value_out_10_15_ready),
    .io_value_out_10_15_valid(core_io_value_out_10_15_valid),
    .io_value_out_10_15_bits(core_io_value_out_10_15_bits),
    .io_value_out_11_0_ready(core_io_value_out_11_0_ready),
    .io_value_out_11_0_valid(core_io_value_out_11_0_valid),
    .io_value_out_11_0_bits(core_io_value_out_11_0_bits),
    .io_value_out_11_1_ready(core_io_value_out_11_1_ready),
    .io_value_out_11_1_valid(core_io_value_out_11_1_valid),
    .io_value_out_11_1_bits(core_io_value_out_11_1_bits),
    .io_value_out_11_2_ready(core_io_value_out_11_2_ready),
    .io_value_out_11_2_valid(core_io_value_out_11_2_valid),
    .io_value_out_11_2_bits(core_io_value_out_11_2_bits),
    .io_value_out_11_3_ready(core_io_value_out_11_3_ready),
    .io_value_out_11_3_valid(core_io_value_out_11_3_valid),
    .io_value_out_11_3_bits(core_io_value_out_11_3_bits),
    .io_value_out_11_4_ready(core_io_value_out_11_4_ready),
    .io_value_out_11_4_valid(core_io_value_out_11_4_valid),
    .io_value_out_11_4_bits(core_io_value_out_11_4_bits),
    .io_value_out_11_5_ready(core_io_value_out_11_5_ready),
    .io_value_out_11_5_valid(core_io_value_out_11_5_valid),
    .io_value_out_11_5_bits(core_io_value_out_11_5_bits),
    .io_value_out_11_6_ready(core_io_value_out_11_6_ready),
    .io_value_out_11_6_valid(core_io_value_out_11_6_valid),
    .io_value_out_11_6_bits(core_io_value_out_11_6_bits),
    .io_value_out_11_7_ready(core_io_value_out_11_7_ready),
    .io_value_out_11_7_valid(core_io_value_out_11_7_valid),
    .io_value_out_11_7_bits(core_io_value_out_11_7_bits),
    .io_value_out_11_8_ready(core_io_value_out_11_8_ready),
    .io_value_out_11_8_valid(core_io_value_out_11_8_valid),
    .io_value_out_11_8_bits(core_io_value_out_11_8_bits),
    .io_value_out_11_9_ready(core_io_value_out_11_9_ready),
    .io_value_out_11_9_valid(core_io_value_out_11_9_valid),
    .io_value_out_11_9_bits(core_io_value_out_11_9_bits),
    .io_value_out_11_10_ready(core_io_value_out_11_10_ready),
    .io_value_out_11_10_valid(core_io_value_out_11_10_valid),
    .io_value_out_11_10_bits(core_io_value_out_11_10_bits),
    .io_value_out_11_11_ready(core_io_value_out_11_11_ready),
    .io_value_out_11_11_valid(core_io_value_out_11_11_valid),
    .io_value_out_11_11_bits(core_io_value_out_11_11_bits),
    .io_value_out_11_12_ready(core_io_value_out_11_12_ready),
    .io_value_out_11_12_valid(core_io_value_out_11_12_valid),
    .io_value_out_11_12_bits(core_io_value_out_11_12_bits),
    .io_value_out_11_13_ready(core_io_value_out_11_13_ready),
    .io_value_out_11_13_valid(core_io_value_out_11_13_valid),
    .io_value_out_11_13_bits(core_io_value_out_11_13_bits),
    .io_value_out_11_14_ready(core_io_value_out_11_14_ready),
    .io_value_out_11_14_valid(core_io_value_out_11_14_valid),
    .io_value_out_11_14_bits(core_io_value_out_11_14_bits),
    .io_value_out_11_15_ready(core_io_value_out_11_15_ready),
    .io_value_out_11_15_valid(core_io_value_out_11_15_valid),
    .io_value_out_11_15_bits(core_io_value_out_11_15_bits),
    .io_value_out_12_0_ready(core_io_value_out_12_0_ready),
    .io_value_out_12_0_valid(core_io_value_out_12_0_valid),
    .io_value_out_12_0_bits(core_io_value_out_12_0_bits),
    .io_value_out_12_1_ready(core_io_value_out_12_1_ready),
    .io_value_out_12_1_valid(core_io_value_out_12_1_valid),
    .io_value_out_12_1_bits(core_io_value_out_12_1_bits),
    .io_value_out_12_2_ready(core_io_value_out_12_2_ready),
    .io_value_out_12_2_valid(core_io_value_out_12_2_valid),
    .io_value_out_12_2_bits(core_io_value_out_12_2_bits),
    .io_value_out_12_3_ready(core_io_value_out_12_3_ready),
    .io_value_out_12_3_valid(core_io_value_out_12_3_valid),
    .io_value_out_12_3_bits(core_io_value_out_12_3_bits),
    .io_value_out_12_4_ready(core_io_value_out_12_4_ready),
    .io_value_out_12_4_valid(core_io_value_out_12_4_valid),
    .io_value_out_12_4_bits(core_io_value_out_12_4_bits),
    .io_value_out_12_5_ready(core_io_value_out_12_5_ready),
    .io_value_out_12_5_valid(core_io_value_out_12_5_valid),
    .io_value_out_12_5_bits(core_io_value_out_12_5_bits),
    .io_value_out_12_6_ready(core_io_value_out_12_6_ready),
    .io_value_out_12_6_valid(core_io_value_out_12_6_valid),
    .io_value_out_12_6_bits(core_io_value_out_12_6_bits),
    .io_value_out_12_7_ready(core_io_value_out_12_7_ready),
    .io_value_out_12_7_valid(core_io_value_out_12_7_valid),
    .io_value_out_12_7_bits(core_io_value_out_12_7_bits),
    .io_value_out_12_8_ready(core_io_value_out_12_8_ready),
    .io_value_out_12_8_valid(core_io_value_out_12_8_valid),
    .io_value_out_12_8_bits(core_io_value_out_12_8_bits),
    .io_value_out_12_9_ready(core_io_value_out_12_9_ready),
    .io_value_out_12_9_valid(core_io_value_out_12_9_valid),
    .io_value_out_12_9_bits(core_io_value_out_12_9_bits),
    .io_value_out_12_10_ready(core_io_value_out_12_10_ready),
    .io_value_out_12_10_valid(core_io_value_out_12_10_valid),
    .io_value_out_12_10_bits(core_io_value_out_12_10_bits),
    .io_value_out_12_11_ready(core_io_value_out_12_11_ready),
    .io_value_out_12_11_valid(core_io_value_out_12_11_valid),
    .io_value_out_12_11_bits(core_io_value_out_12_11_bits),
    .io_value_out_12_12_ready(core_io_value_out_12_12_ready),
    .io_value_out_12_12_valid(core_io_value_out_12_12_valid),
    .io_value_out_12_12_bits(core_io_value_out_12_12_bits),
    .io_value_out_12_13_ready(core_io_value_out_12_13_ready),
    .io_value_out_12_13_valid(core_io_value_out_12_13_valid),
    .io_value_out_12_13_bits(core_io_value_out_12_13_bits),
    .io_value_out_12_14_ready(core_io_value_out_12_14_ready),
    .io_value_out_12_14_valid(core_io_value_out_12_14_valid),
    .io_value_out_12_14_bits(core_io_value_out_12_14_bits),
    .io_value_out_12_15_ready(core_io_value_out_12_15_ready),
    .io_value_out_12_15_valid(core_io_value_out_12_15_valid),
    .io_value_out_12_15_bits(core_io_value_out_12_15_bits),
    .io_value_out_13_0_ready(core_io_value_out_13_0_ready),
    .io_value_out_13_0_valid(core_io_value_out_13_0_valid),
    .io_value_out_13_0_bits(core_io_value_out_13_0_bits),
    .io_value_out_13_1_ready(core_io_value_out_13_1_ready),
    .io_value_out_13_1_valid(core_io_value_out_13_1_valid),
    .io_value_out_13_1_bits(core_io_value_out_13_1_bits),
    .io_value_out_13_2_ready(core_io_value_out_13_2_ready),
    .io_value_out_13_2_valid(core_io_value_out_13_2_valid),
    .io_value_out_13_2_bits(core_io_value_out_13_2_bits),
    .io_value_out_13_3_ready(core_io_value_out_13_3_ready),
    .io_value_out_13_3_valid(core_io_value_out_13_3_valid),
    .io_value_out_13_3_bits(core_io_value_out_13_3_bits),
    .io_value_out_13_4_ready(core_io_value_out_13_4_ready),
    .io_value_out_13_4_valid(core_io_value_out_13_4_valid),
    .io_value_out_13_4_bits(core_io_value_out_13_4_bits),
    .io_value_out_13_5_ready(core_io_value_out_13_5_ready),
    .io_value_out_13_5_valid(core_io_value_out_13_5_valid),
    .io_value_out_13_5_bits(core_io_value_out_13_5_bits),
    .io_value_out_13_6_ready(core_io_value_out_13_6_ready),
    .io_value_out_13_6_valid(core_io_value_out_13_6_valid),
    .io_value_out_13_6_bits(core_io_value_out_13_6_bits),
    .io_value_out_13_7_ready(core_io_value_out_13_7_ready),
    .io_value_out_13_7_valid(core_io_value_out_13_7_valid),
    .io_value_out_13_7_bits(core_io_value_out_13_7_bits),
    .io_value_out_13_8_ready(core_io_value_out_13_8_ready),
    .io_value_out_13_8_valid(core_io_value_out_13_8_valid),
    .io_value_out_13_8_bits(core_io_value_out_13_8_bits),
    .io_value_out_13_9_ready(core_io_value_out_13_9_ready),
    .io_value_out_13_9_valid(core_io_value_out_13_9_valid),
    .io_value_out_13_9_bits(core_io_value_out_13_9_bits),
    .io_value_out_13_10_ready(core_io_value_out_13_10_ready),
    .io_value_out_13_10_valid(core_io_value_out_13_10_valid),
    .io_value_out_13_10_bits(core_io_value_out_13_10_bits),
    .io_value_out_13_11_ready(core_io_value_out_13_11_ready),
    .io_value_out_13_11_valid(core_io_value_out_13_11_valid),
    .io_value_out_13_11_bits(core_io_value_out_13_11_bits),
    .io_value_out_13_12_ready(core_io_value_out_13_12_ready),
    .io_value_out_13_12_valid(core_io_value_out_13_12_valid),
    .io_value_out_13_12_bits(core_io_value_out_13_12_bits),
    .io_value_out_13_13_ready(core_io_value_out_13_13_ready),
    .io_value_out_13_13_valid(core_io_value_out_13_13_valid),
    .io_value_out_13_13_bits(core_io_value_out_13_13_bits),
    .io_value_out_13_14_ready(core_io_value_out_13_14_ready),
    .io_value_out_13_14_valid(core_io_value_out_13_14_valid),
    .io_value_out_13_14_bits(core_io_value_out_13_14_bits),
    .io_value_out_13_15_ready(core_io_value_out_13_15_ready),
    .io_value_out_13_15_valid(core_io_value_out_13_15_valid),
    .io_value_out_13_15_bits(core_io_value_out_13_15_bits),
    .io_value_out_14_0_ready(core_io_value_out_14_0_ready),
    .io_value_out_14_0_valid(core_io_value_out_14_0_valid),
    .io_value_out_14_0_bits(core_io_value_out_14_0_bits),
    .io_value_out_14_1_ready(core_io_value_out_14_1_ready),
    .io_value_out_14_1_valid(core_io_value_out_14_1_valid),
    .io_value_out_14_1_bits(core_io_value_out_14_1_bits),
    .io_value_out_14_2_ready(core_io_value_out_14_2_ready),
    .io_value_out_14_2_valid(core_io_value_out_14_2_valid),
    .io_value_out_14_2_bits(core_io_value_out_14_2_bits),
    .io_value_out_14_3_ready(core_io_value_out_14_3_ready),
    .io_value_out_14_3_valid(core_io_value_out_14_3_valid),
    .io_value_out_14_3_bits(core_io_value_out_14_3_bits),
    .io_value_out_14_4_ready(core_io_value_out_14_4_ready),
    .io_value_out_14_4_valid(core_io_value_out_14_4_valid),
    .io_value_out_14_4_bits(core_io_value_out_14_4_bits),
    .io_value_out_14_5_ready(core_io_value_out_14_5_ready),
    .io_value_out_14_5_valid(core_io_value_out_14_5_valid),
    .io_value_out_14_5_bits(core_io_value_out_14_5_bits),
    .io_value_out_14_6_ready(core_io_value_out_14_6_ready),
    .io_value_out_14_6_valid(core_io_value_out_14_6_valid),
    .io_value_out_14_6_bits(core_io_value_out_14_6_bits),
    .io_value_out_14_7_ready(core_io_value_out_14_7_ready),
    .io_value_out_14_7_valid(core_io_value_out_14_7_valid),
    .io_value_out_14_7_bits(core_io_value_out_14_7_bits),
    .io_value_out_14_8_ready(core_io_value_out_14_8_ready),
    .io_value_out_14_8_valid(core_io_value_out_14_8_valid),
    .io_value_out_14_8_bits(core_io_value_out_14_8_bits),
    .io_value_out_14_9_ready(core_io_value_out_14_9_ready),
    .io_value_out_14_9_valid(core_io_value_out_14_9_valid),
    .io_value_out_14_9_bits(core_io_value_out_14_9_bits),
    .io_value_out_14_10_ready(core_io_value_out_14_10_ready),
    .io_value_out_14_10_valid(core_io_value_out_14_10_valid),
    .io_value_out_14_10_bits(core_io_value_out_14_10_bits),
    .io_value_out_14_11_ready(core_io_value_out_14_11_ready),
    .io_value_out_14_11_valid(core_io_value_out_14_11_valid),
    .io_value_out_14_11_bits(core_io_value_out_14_11_bits),
    .io_value_out_14_12_ready(core_io_value_out_14_12_ready),
    .io_value_out_14_12_valid(core_io_value_out_14_12_valid),
    .io_value_out_14_12_bits(core_io_value_out_14_12_bits),
    .io_value_out_14_13_ready(core_io_value_out_14_13_ready),
    .io_value_out_14_13_valid(core_io_value_out_14_13_valid),
    .io_value_out_14_13_bits(core_io_value_out_14_13_bits),
    .io_value_out_14_14_ready(core_io_value_out_14_14_ready),
    .io_value_out_14_14_valid(core_io_value_out_14_14_valid),
    .io_value_out_14_14_bits(core_io_value_out_14_14_bits),
    .io_value_out_14_15_ready(core_io_value_out_14_15_ready),
    .io_value_out_14_15_valid(core_io_value_out_14_15_valid),
    .io_value_out_14_15_bits(core_io_value_out_14_15_bits),
    .io_value_out_15_0_ready(core_io_value_out_15_0_ready),
    .io_value_out_15_0_valid(core_io_value_out_15_0_valid),
    .io_value_out_15_0_bits(core_io_value_out_15_0_bits),
    .io_value_out_15_1_ready(core_io_value_out_15_1_ready),
    .io_value_out_15_1_valid(core_io_value_out_15_1_valid),
    .io_value_out_15_1_bits(core_io_value_out_15_1_bits),
    .io_value_out_15_2_ready(core_io_value_out_15_2_ready),
    .io_value_out_15_2_valid(core_io_value_out_15_2_valid),
    .io_value_out_15_2_bits(core_io_value_out_15_2_bits),
    .io_value_out_15_3_ready(core_io_value_out_15_3_ready),
    .io_value_out_15_3_valid(core_io_value_out_15_3_valid),
    .io_value_out_15_3_bits(core_io_value_out_15_3_bits),
    .io_value_out_15_4_ready(core_io_value_out_15_4_ready),
    .io_value_out_15_4_valid(core_io_value_out_15_4_valid),
    .io_value_out_15_4_bits(core_io_value_out_15_4_bits),
    .io_value_out_15_5_ready(core_io_value_out_15_5_ready),
    .io_value_out_15_5_valid(core_io_value_out_15_5_valid),
    .io_value_out_15_5_bits(core_io_value_out_15_5_bits),
    .io_value_out_15_6_ready(core_io_value_out_15_6_ready),
    .io_value_out_15_6_valid(core_io_value_out_15_6_valid),
    .io_value_out_15_6_bits(core_io_value_out_15_6_bits),
    .io_value_out_15_7_ready(core_io_value_out_15_7_ready),
    .io_value_out_15_7_valid(core_io_value_out_15_7_valid),
    .io_value_out_15_7_bits(core_io_value_out_15_7_bits),
    .io_value_out_15_8_ready(core_io_value_out_15_8_ready),
    .io_value_out_15_8_valid(core_io_value_out_15_8_valid),
    .io_value_out_15_8_bits(core_io_value_out_15_8_bits),
    .io_value_out_15_9_ready(core_io_value_out_15_9_ready),
    .io_value_out_15_9_valid(core_io_value_out_15_9_valid),
    .io_value_out_15_9_bits(core_io_value_out_15_9_bits),
    .io_value_out_15_10_ready(core_io_value_out_15_10_ready),
    .io_value_out_15_10_valid(core_io_value_out_15_10_valid),
    .io_value_out_15_10_bits(core_io_value_out_15_10_bits),
    .io_value_out_15_11_ready(core_io_value_out_15_11_ready),
    .io_value_out_15_11_valid(core_io_value_out_15_11_valid),
    .io_value_out_15_11_bits(core_io_value_out_15_11_bits),
    .io_value_out_15_12_ready(core_io_value_out_15_12_ready),
    .io_value_out_15_12_valid(core_io_value_out_15_12_valid),
    .io_value_out_15_12_bits(core_io_value_out_15_12_bits),
    .io_value_out_15_13_ready(core_io_value_out_15_13_ready),
    .io_value_out_15_13_valid(core_io_value_out_15_13_valid),
    .io_value_out_15_13_bits(core_io_value_out_15_13_bits),
    .io_value_out_15_14_ready(core_io_value_out_15_14_ready),
    .io_value_out_15_14_valid(core_io_value_out_15_14_valid),
    .io_value_out_15_14_bits(core_io_value_out_15_14_bits),
    .io_value_out_15_15_ready(core_io_value_out_15_15_ready),
    .io_value_out_15_15_valid(core_io_value_out_15_15_valid),
    .io_value_out_15_15_bits(core_io_value_out_15_15_bits)
  );
  StreamTranspose wsplit ( // @[Stab.scala 314:22]
    .clock(wsplit_clock),
    .reset(wsplit_reset),
    .io_stream_in_ready(wsplit_io_stream_in_ready),
    .io_stream_in_valid(wsplit_io_stream_in_valid),
    .io_stream_in_bits(wsplit_io_stream_in_bits),
    .io_stream_out_0_ready(wsplit_io_stream_out_0_ready),
    .io_stream_out_0_valid(wsplit_io_stream_out_0_valid),
    .io_stream_out_0_bits(wsplit_io_stream_out_0_bits),
    .io_stream_out_1_ready(wsplit_io_stream_out_1_ready),
    .io_stream_out_1_valid(wsplit_io_stream_out_1_valid),
    .io_stream_out_1_bits(wsplit_io_stream_out_1_bits),
    .io_stream_out_2_ready(wsplit_io_stream_out_2_ready),
    .io_stream_out_2_valid(wsplit_io_stream_out_2_valid),
    .io_stream_out_2_bits(wsplit_io_stream_out_2_bits),
    .io_stream_out_3_ready(wsplit_io_stream_out_3_ready),
    .io_stream_out_3_valid(wsplit_io_stream_out_3_valid),
    .io_stream_out_3_bits(wsplit_io_stream_out_3_bits),
    .io_stream_out_4_ready(wsplit_io_stream_out_4_ready),
    .io_stream_out_4_valid(wsplit_io_stream_out_4_valid),
    .io_stream_out_4_bits(wsplit_io_stream_out_4_bits),
    .io_stream_out_5_ready(wsplit_io_stream_out_5_ready),
    .io_stream_out_5_valid(wsplit_io_stream_out_5_valid),
    .io_stream_out_5_bits(wsplit_io_stream_out_5_bits),
    .io_stream_out_6_ready(wsplit_io_stream_out_6_ready),
    .io_stream_out_6_valid(wsplit_io_stream_out_6_valid),
    .io_stream_out_6_bits(wsplit_io_stream_out_6_bits),
    .io_stream_out_7_ready(wsplit_io_stream_out_7_ready),
    .io_stream_out_7_valid(wsplit_io_stream_out_7_valid),
    .io_stream_out_7_bits(wsplit_io_stream_out_7_bits),
    .io_stream_out_8_ready(wsplit_io_stream_out_8_ready),
    .io_stream_out_8_valid(wsplit_io_stream_out_8_valid),
    .io_stream_out_8_bits(wsplit_io_stream_out_8_bits),
    .io_stream_out_9_ready(wsplit_io_stream_out_9_ready),
    .io_stream_out_9_valid(wsplit_io_stream_out_9_valid),
    .io_stream_out_9_bits(wsplit_io_stream_out_9_bits),
    .io_stream_out_10_ready(wsplit_io_stream_out_10_ready),
    .io_stream_out_10_valid(wsplit_io_stream_out_10_valid),
    .io_stream_out_10_bits(wsplit_io_stream_out_10_bits),
    .io_stream_out_11_ready(wsplit_io_stream_out_11_ready),
    .io_stream_out_11_valid(wsplit_io_stream_out_11_valid),
    .io_stream_out_11_bits(wsplit_io_stream_out_11_bits),
    .io_stream_out_12_ready(wsplit_io_stream_out_12_ready),
    .io_stream_out_12_valid(wsplit_io_stream_out_12_valid),
    .io_stream_out_12_bits(wsplit_io_stream_out_12_bits),
    .io_stream_out_13_ready(wsplit_io_stream_out_13_ready),
    .io_stream_out_13_valid(wsplit_io_stream_out_13_valid),
    .io_stream_out_13_bits(wsplit_io_stream_out_13_bits),
    .io_stream_out_14_ready(wsplit_io_stream_out_14_ready),
    .io_stream_out_14_valid(wsplit_io_stream_out_14_valid),
    .io_stream_out_14_bits(wsplit_io_stream_out_14_bits),
    .io_stream_out_15_ready(wsplit_io_stream_out_15_ready),
    .io_stream_out_15_valid(wsplit_io_stream_out_15_valid),
    .io_stream_out_15_bits(wsplit_io_stream_out_15_bits)
  );
  StreamTranspose vsplit ( // @[Stab.scala 315:22]
    .clock(vsplit_clock),
    .reset(vsplit_reset),
    .io_stream_in_ready(vsplit_io_stream_in_ready),
    .io_stream_in_valid(vsplit_io_stream_in_valid),
    .io_stream_in_bits(vsplit_io_stream_in_bits),
    .io_stream_out_0_ready(vsplit_io_stream_out_0_ready),
    .io_stream_out_0_valid(vsplit_io_stream_out_0_valid),
    .io_stream_out_0_bits(vsplit_io_stream_out_0_bits),
    .io_stream_out_1_ready(vsplit_io_stream_out_1_ready),
    .io_stream_out_1_valid(vsplit_io_stream_out_1_valid),
    .io_stream_out_1_bits(vsplit_io_stream_out_1_bits),
    .io_stream_out_2_ready(vsplit_io_stream_out_2_ready),
    .io_stream_out_2_valid(vsplit_io_stream_out_2_valid),
    .io_stream_out_2_bits(vsplit_io_stream_out_2_bits),
    .io_stream_out_3_ready(vsplit_io_stream_out_3_ready),
    .io_stream_out_3_valid(vsplit_io_stream_out_3_valid),
    .io_stream_out_3_bits(vsplit_io_stream_out_3_bits),
    .io_stream_out_4_ready(vsplit_io_stream_out_4_ready),
    .io_stream_out_4_valid(vsplit_io_stream_out_4_valid),
    .io_stream_out_4_bits(vsplit_io_stream_out_4_bits),
    .io_stream_out_5_ready(vsplit_io_stream_out_5_ready),
    .io_stream_out_5_valid(vsplit_io_stream_out_5_valid),
    .io_stream_out_5_bits(vsplit_io_stream_out_5_bits),
    .io_stream_out_6_ready(vsplit_io_stream_out_6_ready),
    .io_stream_out_6_valid(vsplit_io_stream_out_6_valid),
    .io_stream_out_6_bits(vsplit_io_stream_out_6_bits),
    .io_stream_out_7_ready(vsplit_io_stream_out_7_ready),
    .io_stream_out_7_valid(vsplit_io_stream_out_7_valid),
    .io_stream_out_7_bits(vsplit_io_stream_out_7_bits),
    .io_stream_out_8_ready(vsplit_io_stream_out_8_ready),
    .io_stream_out_8_valid(vsplit_io_stream_out_8_valid),
    .io_stream_out_8_bits(vsplit_io_stream_out_8_bits),
    .io_stream_out_9_ready(vsplit_io_stream_out_9_ready),
    .io_stream_out_9_valid(vsplit_io_stream_out_9_valid),
    .io_stream_out_9_bits(vsplit_io_stream_out_9_bits),
    .io_stream_out_10_ready(vsplit_io_stream_out_10_ready),
    .io_stream_out_10_valid(vsplit_io_stream_out_10_valid),
    .io_stream_out_10_bits(vsplit_io_stream_out_10_bits),
    .io_stream_out_11_ready(vsplit_io_stream_out_11_ready),
    .io_stream_out_11_valid(vsplit_io_stream_out_11_valid),
    .io_stream_out_11_bits(vsplit_io_stream_out_11_bits),
    .io_stream_out_12_ready(vsplit_io_stream_out_12_ready),
    .io_stream_out_12_valid(vsplit_io_stream_out_12_valid),
    .io_stream_out_12_bits(vsplit_io_stream_out_12_bits),
    .io_stream_out_13_ready(vsplit_io_stream_out_13_ready),
    .io_stream_out_13_valid(vsplit_io_stream_out_13_valid),
    .io_stream_out_13_bits(vsplit_io_stream_out_13_bits),
    .io_stream_out_14_ready(vsplit_io_stream_out_14_ready),
    .io_stream_out_14_valid(vsplit_io_stream_out_14_valid),
    .io_stream_out_14_bits(vsplit_io_stream_out_14_bits),
    .io_stream_out_15_ready(vsplit_io_stream_out_15_ready),
    .io_stream_out_15_valid(vsplit_io_stream_out_15_valid),
    .io_stream_out_15_bits(vsplit_io_stream_out_15_bits)
  );
  StreamAggregator rmerge ( // @[Stab.scala 317:22]
    .clock(rmerge_clock),
    .reset(rmerge_reset),
    .io_stream_in_0_ready(rmerge_io_stream_in_0_ready),
    .io_stream_in_0_valid(rmerge_io_stream_in_0_valid),
    .io_stream_in_0_bits(rmerge_io_stream_in_0_bits),
    .io_stream_in_1_ready(rmerge_io_stream_in_1_ready),
    .io_stream_in_1_valid(rmerge_io_stream_in_1_valid),
    .io_stream_in_1_bits(rmerge_io_stream_in_1_bits),
    .io_stream_in_2_ready(rmerge_io_stream_in_2_ready),
    .io_stream_in_2_valid(rmerge_io_stream_in_2_valid),
    .io_stream_in_2_bits(rmerge_io_stream_in_2_bits),
    .io_stream_in_3_ready(rmerge_io_stream_in_3_ready),
    .io_stream_in_3_valid(rmerge_io_stream_in_3_valid),
    .io_stream_in_3_bits(rmerge_io_stream_in_3_bits),
    .io_stream_in_4_ready(rmerge_io_stream_in_4_ready),
    .io_stream_in_4_valid(rmerge_io_stream_in_4_valid),
    .io_stream_in_4_bits(rmerge_io_stream_in_4_bits),
    .io_stream_in_5_ready(rmerge_io_stream_in_5_ready),
    .io_stream_in_5_valid(rmerge_io_stream_in_5_valid),
    .io_stream_in_5_bits(rmerge_io_stream_in_5_bits),
    .io_stream_in_6_ready(rmerge_io_stream_in_6_ready),
    .io_stream_in_6_valid(rmerge_io_stream_in_6_valid),
    .io_stream_in_6_bits(rmerge_io_stream_in_6_bits),
    .io_stream_in_7_ready(rmerge_io_stream_in_7_ready),
    .io_stream_in_7_valid(rmerge_io_stream_in_7_valid),
    .io_stream_in_7_bits(rmerge_io_stream_in_7_bits),
    .io_stream_in_8_ready(rmerge_io_stream_in_8_ready),
    .io_stream_in_8_valid(rmerge_io_stream_in_8_valid),
    .io_stream_in_8_bits(rmerge_io_stream_in_8_bits),
    .io_stream_in_9_ready(rmerge_io_stream_in_9_ready),
    .io_stream_in_9_valid(rmerge_io_stream_in_9_valid),
    .io_stream_in_9_bits(rmerge_io_stream_in_9_bits),
    .io_stream_in_10_ready(rmerge_io_stream_in_10_ready),
    .io_stream_in_10_valid(rmerge_io_stream_in_10_valid),
    .io_stream_in_10_bits(rmerge_io_stream_in_10_bits),
    .io_stream_in_11_ready(rmerge_io_stream_in_11_ready),
    .io_stream_in_11_valid(rmerge_io_stream_in_11_valid),
    .io_stream_in_11_bits(rmerge_io_stream_in_11_bits),
    .io_stream_in_12_ready(rmerge_io_stream_in_12_ready),
    .io_stream_in_12_valid(rmerge_io_stream_in_12_valid),
    .io_stream_in_12_bits(rmerge_io_stream_in_12_bits),
    .io_stream_in_13_ready(rmerge_io_stream_in_13_ready),
    .io_stream_in_13_valid(rmerge_io_stream_in_13_valid),
    .io_stream_in_13_bits(rmerge_io_stream_in_13_bits),
    .io_stream_in_14_ready(rmerge_io_stream_in_14_ready),
    .io_stream_in_14_valid(rmerge_io_stream_in_14_valid),
    .io_stream_in_14_bits(rmerge_io_stream_in_14_bits),
    .io_stream_in_15_ready(rmerge_io_stream_in_15_ready),
    .io_stream_in_15_valid(rmerge_io_stream_in_15_valid),
    .io_stream_in_15_bits(rmerge_io_stream_in_15_bits),
    .io_stream_in_16_ready(rmerge_io_stream_in_16_ready),
    .io_stream_in_16_valid(rmerge_io_stream_in_16_valid),
    .io_stream_in_16_bits(rmerge_io_stream_in_16_bits),
    .io_stream_in_17_ready(rmerge_io_stream_in_17_ready),
    .io_stream_in_17_valid(rmerge_io_stream_in_17_valid),
    .io_stream_in_17_bits(rmerge_io_stream_in_17_bits),
    .io_stream_in_18_ready(rmerge_io_stream_in_18_ready),
    .io_stream_in_18_valid(rmerge_io_stream_in_18_valid),
    .io_stream_in_18_bits(rmerge_io_stream_in_18_bits),
    .io_stream_in_19_ready(rmerge_io_stream_in_19_ready),
    .io_stream_in_19_valid(rmerge_io_stream_in_19_valid),
    .io_stream_in_19_bits(rmerge_io_stream_in_19_bits),
    .io_stream_in_20_ready(rmerge_io_stream_in_20_ready),
    .io_stream_in_20_valid(rmerge_io_stream_in_20_valid),
    .io_stream_in_20_bits(rmerge_io_stream_in_20_bits),
    .io_stream_in_21_ready(rmerge_io_stream_in_21_ready),
    .io_stream_in_21_valid(rmerge_io_stream_in_21_valid),
    .io_stream_in_21_bits(rmerge_io_stream_in_21_bits),
    .io_stream_in_22_ready(rmerge_io_stream_in_22_ready),
    .io_stream_in_22_valid(rmerge_io_stream_in_22_valid),
    .io_stream_in_22_bits(rmerge_io_stream_in_22_bits),
    .io_stream_in_23_ready(rmerge_io_stream_in_23_ready),
    .io_stream_in_23_valid(rmerge_io_stream_in_23_valid),
    .io_stream_in_23_bits(rmerge_io_stream_in_23_bits),
    .io_stream_in_24_ready(rmerge_io_stream_in_24_ready),
    .io_stream_in_24_valid(rmerge_io_stream_in_24_valid),
    .io_stream_in_24_bits(rmerge_io_stream_in_24_bits),
    .io_stream_in_25_ready(rmerge_io_stream_in_25_ready),
    .io_stream_in_25_valid(rmerge_io_stream_in_25_valid),
    .io_stream_in_25_bits(rmerge_io_stream_in_25_bits),
    .io_stream_in_26_ready(rmerge_io_stream_in_26_ready),
    .io_stream_in_26_valid(rmerge_io_stream_in_26_valid),
    .io_stream_in_26_bits(rmerge_io_stream_in_26_bits),
    .io_stream_in_27_ready(rmerge_io_stream_in_27_ready),
    .io_stream_in_27_valid(rmerge_io_stream_in_27_valid),
    .io_stream_in_27_bits(rmerge_io_stream_in_27_bits),
    .io_stream_in_28_ready(rmerge_io_stream_in_28_ready),
    .io_stream_in_28_valid(rmerge_io_stream_in_28_valid),
    .io_stream_in_28_bits(rmerge_io_stream_in_28_bits),
    .io_stream_in_29_ready(rmerge_io_stream_in_29_ready),
    .io_stream_in_29_valid(rmerge_io_stream_in_29_valid),
    .io_stream_in_29_bits(rmerge_io_stream_in_29_bits),
    .io_stream_in_30_ready(rmerge_io_stream_in_30_ready),
    .io_stream_in_30_valid(rmerge_io_stream_in_30_valid),
    .io_stream_in_30_bits(rmerge_io_stream_in_30_bits),
    .io_stream_in_31_ready(rmerge_io_stream_in_31_ready),
    .io_stream_in_31_valid(rmerge_io_stream_in_31_valid),
    .io_stream_in_31_bits(rmerge_io_stream_in_31_bits),
    .io_stream_in_32_ready(rmerge_io_stream_in_32_ready),
    .io_stream_in_32_valid(rmerge_io_stream_in_32_valid),
    .io_stream_in_32_bits(rmerge_io_stream_in_32_bits),
    .io_stream_in_33_ready(rmerge_io_stream_in_33_ready),
    .io_stream_in_33_valid(rmerge_io_stream_in_33_valid),
    .io_stream_in_33_bits(rmerge_io_stream_in_33_bits),
    .io_stream_in_34_ready(rmerge_io_stream_in_34_ready),
    .io_stream_in_34_valid(rmerge_io_stream_in_34_valid),
    .io_stream_in_34_bits(rmerge_io_stream_in_34_bits),
    .io_stream_in_35_ready(rmerge_io_stream_in_35_ready),
    .io_stream_in_35_valid(rmerge_io_stream_in_35_valid),
    .io_stream_in_35_bits(rmerge_io_stream_in_35_bits),
    .io_stream_in_36_ready(rmerge_io_stream_in_36_ready),
    .io_stream_in_36_valid(rmerge_io_stream_in_36_valid),
    .io_stream_in_36_bits(rmerge_io_stream_in_36_bits),
    .io_stream_in_37_ready(rmerge_io_stream_in_37_ready),
    .io_stream_in_37_valid(rmerge_io_stream_in_37_valid),
    .io_stream_in_37_bits(rmerge_io_stream_in_37_bits),
    .io_stream_in_38_ready(rmerge_io_stream_in_38_ready),
    .io_stream_in_38_valid(rmerge_io_stream_in_38_valid),
    .io_stream_in_38_bits(rmerge_io_stream_in_38_bits),
    .io_stream_in_39_ready(rmerge_io_stream_in_39_ready),
    .io_stream_in_39_valid(rmerge_io_stream_in_39_valid),
    .io_stream_in_39_bits(rmerge_io_stream_in_39_bits),
    .io_stream_in_40_ready(rmerge_io_stream_in_40_ready),
    .io_stream_in_40_valid(rmerge_io_stream_in_40_valid),
    .io_stream_in_40_bits(rmerge_io_stream_in_40_bits),
    .io_stream_in_41_ready(rmerge_io_stream_in_41_ready),
    .io_stream_in_41_valid(rmerge_io_stream_in_41_valid),
    .io_stream_in_41_bits(rmerge_io_stream_in_41_bits),
    .io_stream_in_42_ready(rmerge_io_stream_in_42_ready),
    .io_stream_in_42_valid(rmerge_io_stream_in_42_valid),
    .io_stream_in_42_bits(rmerge_io_stream_in_42_bits),
    .io_stream_in_43_ready(rmerge_io_stream_in_43_ready),
    .io_stream_in_43_valid(rmerge_io_stream_in_43_valid),
    .io_stream_in_43_bits(rmerge_io_stream_in_43_bits),
    .io_stream_in_44_ready(rmerge_io_stream_in_44_ready),
    .io_stream_in_44_valid(rmerge_io_stream_in_44_valid),
    .io_stream_in_44_bits(rmerge_io_stream_in_44_bits),
    .io_stream_in_45_ready(rmerge_io_stream_in_45_ready),
    .io_stream_in_45_valid(rmerge_io_stream_in_45_valid),
    .io_stream_in_45_bits(rmerge_io_stream_in_45_bits),
    .io_stream_in_46_ready(rmerge_io_stream_in_46_ready),
    .io_stream_in_46_valid(rmerge_io_stream_in_46_valid),
    .io_stream_in_46_bits(rmerge_io_stream_in_46_bits),
    .io_stream_in_47_ready(rmerge_io_stream_in_47_ready),
    .io_stream_in_47_valid(rmerge_io_stream_in_47_valid),
    .io_stream_in_47_bits(rmerge_io_stream_in_47_bits),
    .io_stream_in_48_ready(rmerge_io_stream_in_48_ready),
    .io_stream_in_48_valid(rmerge_io_stream_in_48_valid),
    .io_stream_in_48_bits(rmerge_io_stream_in_48_bits),
    .io_stream_in_49_ready(rmerge_io_stream_in_49_ready),
    .io_stream_in_49_valid(rmerge_io_stream_in_49_valid),
    .io_stream_in_49_bits(rmerge_io_stream_in_49_bits),
    .io_stream_in_50_ready(rmerge_io_stream_in_50_ready),
    .io_stream_in_50_valid(rmerge_io_stream_in_50_valid),
    .io_stream_in_50_bits(rmerge_io_stream_in_50_bits),
    .io_stream_in_51_ready(rmerge_io_stream_in_51_ready),
    .io_stream_in_51_valid(rmerge_io_stream_in_51_valid),
    .io_stream_in_51_bits(rmerge_io_stream_in_51_bits),
    .io_stream_in_52_ready(rmerge_io_stream_in_52_ready),
    .io_stream_in_52_valid(rmerge_io_stream_in_52_valid),
    .io_stream_in_52_bits(rmerge_io_stream_in_52_bits),
    .io_stream_in_53_ready(rmerge_io_stream_in_53_ready),
    .io_stream_in_53_valid(rmerge_io_stream_in_53_valid),
    .io_stream_in_53_bits(rmerge_io_stream_in_53_bits),
    .io_stream_in_54_ready(rmerge_io_stream_in_54_ready),
    .io_stream_in_54_valid(rmerge_io_stream_in_54_valid),
    .io_stream_in_54_bits(rmerge_io_stream_in_54_bits),
    .io_stream_in_55_ready(rmerge_io_stream_in_55_ready),
    .io_stream_in_55_valid(rmerge_io_stream_in_55_valid),
    .io_stream_in_55_bits(rmerge_io_stream_in_55_bits),
    .io_stream_in_56_ready(rmerge_io_stream_in_56_ready),
    .io_stream_in_56_valid(rmerge_io_stream_in_56_valid),
    .io_stream_in_56_bits(rmerge_io_stream_in_56_bits),
    .io_stream_in_57_ready(rmerge_io_stream_in_57_ready),
    .io_stream_in_57_valid(rmerge_io_stream_in_57_valid),
    .io_stream_in_57_bits(rmerge_io_stream_in_57_bits),
    .io_stream_in_58_ready(rmerge_io_stream_in_58_ready),
    .io_stream_in_58_valid(rmerge_io_stream_in_58_valid),
    .io_stream_in_58_bits(rmerge_io_stream_in_58_bits),
    .io_stream_in_59_ready(rmerge_io_stream_in_59_ready),
    .io_stream_in_59_valid(rmerge_io_stream_in_59_valid),
    .io_stream_in_59_bits(rmerge_io_stream_in_59_bits),
    .io_stream_in_60_ready(rmerge_io_stream_in_60_ready),
    .io_stream_in_60_valid(rmerge_io_stream_in_60_valid),
    .io_stream_in_60_bits(rmerge_io_stream_in_60_bits),
    .io_stream_in_61_ready(rmerge_io_stream_in_61_ready),
    .io_stream_in_61_valid(rmerge_io_stream_in_61_valid),
    .io_stream_in_61_bits(rmerge_io_stream_in_61_bits),
    .io_stream_in_62_ready(rmerge_io_stream_in_62_ready),
    .io_stream_in_62_valid(rmerge_io_stream_in_62_valid),
    .io_stream_in_62_bits(rmerge_io_stream_in_62_bits),
    .io_stream_in_63_ready(rmerge_io_stream_in_63_ready),
    .io_stream_in_63_valid(rmerge_io_stream_in_63_valid),
    .io_stream_in_63_bits(rmerge_io_stream_in_63_bits),
    .io_stream_in_64_ready(rmerge_io_stream_in_64_ready),
    .io_stream_in_64_valid(rmerge_io_stream_in_64_valid),
    .io_stream_in_64_bits(rmerge_io_stream_in_64_bits),
    .io_stream_in_65_ready(rmerge_io_stream_in_65_ready),
    .io_stream_in_65_valid(rmerge_io_stream_in_65_valid),
    .io_stream_in_65_bits(rmerge_io_stream_in_65_bits),
    .io_stream_in_66_ready(rmerge_io_stream_in_66_ready),
    .io_stream_in_66_valid(rmerge_io_stream_in_66_valid),
    .io_stream_in_66_bits(rmerge_io_stream_in_66_bits),
    .io_stream_in_67_ready(rmerge_io_stream_in_67_ready),
    .io_stream_in_67_valid(rmerge_io_stream_in_67_valid),
    .io_stream_in_67_bits(rmerge_io_stream_in_67_bits),
    .io_stream_in_68_ready(rmerge_io_stream_in_68_ready),
    .io_stream_in_68_valid(rmerge_io_stream_in_68_valid),
    .io_stream_in_68_bits(rmerge_io_stream_in_68_bits),
    .io_stream_in_69_ready(rmerge_io_stream_in_69_ready),
    .io_stream_in_69_valid(rmerge_io_stream_in_69_valid),
    .io_stream_in_69_bits(rmerge_io_stream_in_69_bits),
    .io_stream_in_70_ready(rmerge_io_stream_in_70_ready),
    .io_stream_in_70_valid(rmerge_io_stream_in_70_valid),
    .io_stream_in_70_bits(rmerge_io_stream_in_70_bits),
    .io_stream_in_71_ready(rmerge_io_stream_in_71_ready),
    .io_stream_in_71_valid(rmerge_io_stream_in_71_valid),
    .io_stream_in_71_bits(rmerge_io_stream_in_71_bits),
    .io_stream_in_72_ready(rmerge_io_stream_in_72_ready),
    .io_stream_in_72_valid(rmerge_io_stream_in_72_valid),
    .io_stream_in_72_bits(rmerge_io_stream_in_72_bits),
    .io_stream_in_73_ready(rmerge_io_stream_in_73_ready),
    .io_stream_in_73_valid(rmerge_io_stream_in_73_valid),
    .io_stream_in_73_bits(rmerge_io_stream_in_73_bits),
    .io_stream_in_74_ready(rmerge_io_stream_in_74_ready),
    .io_stream_in_74_valid(rmerge_io_stream_in_74_valid),
    .io_stream_in_74_bits(rmerge_io_stream_in_74_bits),
    .io_stream_in_75_ready(rmerge_io_stream_in_75_ready),
    .io_stream_in_75_valid(rmerge_io_stream_in_75_valid),
    .io_stream_in_75_bits(rmerge_io_stream_in_75_bits),
    .io_stream_in_76_ready(rmerge_io_stream_in_76_ready),
    .io_stream_in_76_valid(rmerge_io_stream_in_76_valid),
    .io_stream_in_76_bits(rmerge_io_stream_in_76_bits),
    .io_stream_in_77_ready(rmerge_io_stream_in_77_ready),
    .io_stream_in_77_valid(rmerge_io_stream_in_77_valid),
    .io_stream_in_77_bits(rmerge_io_stream_in_77_bits),
    .io_stream_in_78_ready(rmerge_io_stream_in_78_ready),
    .io_stream_in_78_valid(rmerge_io_stream_in_78_valid),
    .io_stream_in_78_bits(rmerge_io_stream_in_78_bits),
    .io_stream_in_79_ready(rmerge_io_stream_in_79_ready),
    .io_stream_in_79_valid(rmerge_io_stream_in_79_valid),
    .io_stream_in_79_bits(rmerge_io_stream_in_79_bits),
    .io_stream_in_80_ready(rmerge_io_stream_in_80_ready),
    .io_stream_in_80_valid(rmerge_io_stream_in_80_valid),
    .io_stream_in_80_bits(rmerge_io_stream_in_80_bits),
    .io_stream_in_81_ready(rmerge_io_stream_in_81_ready),
    .io_stream_in_81_valid(rmerge_io_stream_in_81_valid),
    .io_stream_in_81_bits(rmerge_io_stream_in_81_bits),
    .io_stream_in_82_ready(rmerge_io_stream_in_82_ready),
    .io_stream_in_82_valid(rmerge_io_stream_in_82_valid),
    .io_stream_in_82_bits(rmerge_io_stream_in_82_bits),
    .io_stream_in_83_ready(rmerge_io_stream_in_83_ready),
    .io_stream_in_83_valid(rmerge_io_stream_in_83_valid),
    .io_stream_in_83_bits(rmerge_io_stream_in_83_bits),
    .io_stream_in_84_ready(rmerge_io_stream_in_84_ready),
    .io_stream_in_84_valid(rmerge_io_stream_in_84_valid),
    .io_stream_in_84_bits(rmerge_io_stream_in_84_bits),
    .io_stream_in_85_ready(rmerge_io_stream_in_85_ready),
    .io_stream_in_85_valid(rmerge_io_stream_in_85_valid),
    .io_stream_in_85_bits(rmerge_io_stream_in_85_bits),
    .io_stream_in_86_ready(rmerge_io_stream_in_86_ready),
    .io_stream_in_86_valid(rmerge_io_stream_in_86_valid),
    .io_stream_in_86_bits(rmerge_io_stream_in_86_bits),
    .io_stream_in_87_ready(rmerge_io_stream_in_87_ready),
    .io_stream_in_87_valid(rmerge_io_stream_in_87_valid),
    .io_stream_in_87_bits(rmerge_io_stream_in_87_bits),
    .io_stream_in_88_ready(rmerge_io_stream_in_88_ready),
    .io_stream_in_88_valid(rmerge_io_stream_in_88_valid),
    .io_stream_in_88_bits(rmerge_io_stream_in_88_bits),
    .io_stream_in_89_ready(rmerge_io_stream_in_89_ready),
    .io_stream_in_89_valid(rmerge_io_stream_in_89_valid),
    .io_stream_in_89_bits(rmerge_io_stream_in_89_bits),
    .io_stream_in_90_ready(rmerge_io_stream_in_90_ready),
    .io_stream_in_90_valid(rmerge_io_stream_in_90_valid),
    .io_stream_in_90_bits(rmerge_io_stream_in_90_bits),
    .io_stream_in_91_ready(rmerge_io_stream_in_91_ready),
    .io_stream_in_91_valid(rmerge_io_stream_in_91_valid),
    .io_stream_in_91_bits(rmerge_io_stream_in_91_bits),
    .io_stream_in_92_ready(rmerge_io_stream_in_92_ready),
    .io_stream_in_92_valid(rmerge_io_stream_in_92_valid),
    .io_stream_in_92_bits(rmerge_io_stream_in_92_bits),
    .io_stream_in_93_ready(rmerge_io_stream_in_93_ready),
    .io_stream_in_93_valid(rmerge_io_stream_in_93_valid),
    .io_stream_in_93_bits(rmerge_io_stream_in_93_bits),
    .io_stream_in_94_ready(rmerge_io_stream_in_94_ready),
    .io_stream_in_94_valid(rmerge_io_stream_in_94_valid),
    .io_stream_in_94_bits(rmerge_io_stream_in_94_bits),
    .io_stream_in_95_ready(rmerge_io_stream_in_95_ready),
    .io_stream_in_95_valid(rmerge_io_stream_in_95_valid),
    .io_stream_in_95_bits(rmerge_io_stream_in_95_bits),
    .io_stream_in_96_ready(rmerge_io_stream_in_96_ready),
    .io_stream_in_96_valid(rmerge_io_stream_in_96_valid),
    .io_stream_in_96_bits(rmerge_io_stream_in_96_bits),
    .io_stream_in_97_ready(rmerge_io_stream_in_97_ready),
    .io_stream_in_97_valid(rmerge_io_stream_in_97_valid),
    .io_stream_in_97_bits(rmerge_io_stream_in_97_bits),
    .io_stream_in_98_ready(rmerge_io_stream_in_98_ready),
    .io_stream_in_98_valid(rmerge_io_stream_in_98_valid),
    .io_stream_in_98_bits(rmerge_io_stream_in_98_bits),
    .io_stream_in_99_ready(rmerge_io_stream_in_99_ready),
    .io_stream_in_99_valid(rmerge_io_stream_in_99_valid),
    .io_stream_in_99_bits(rmerge_io_stream_in_99_bits),
    .io_stream_in_100_ready(rmerge_io_stream_in_100_ready),
    .io_stream_in_100_valid(rmerge_io_stream_in_100_valid),
    .io_stream_in_100_bits(rmerge_io_stream_in_100_bits),
    .io_stream_in_101_ready(rmerge_io_stream_in_101_ready),
    .io_stream_in_101_valid(rmerge_io_stream_in_101_valid),
    .io_stream_in_101_bits(rmerge_io_stream_in_101_bits),
    .io_stream_in_102_ready(rmerge_io_stream_in_102_ready),
    .io_stream_in_102_valid(rmerge_io_stream_in_102_valid),
    .io_stream_in_102_bits(rmerge_io_stream_in_102_bits),
    .io_stream_in_103_ready(rmerge_io_stream_in_103_ready),
    .io_stream_in_103_valid(rmerge_io_stream_in_103_valid),
    .io_stream_in_103_bits(rmerge_io_stream_in_103_bits),
    .io_stream_in_104_ready(rmerge_io_stream_in_104_ready),
    .io_stream_in_104_valid(rmerge_io_stream_in_104_valid),
    .io_stream_in_104_bits(rmerge_io_stream_in_104_bits),
    .io_stream_in_105_ready(rmerge_io_stream_in_105_ready),
    .io_stream_in_105_valid(rmerge_io_stream_in_105_valid),
    .io_stream_in_105_bits(rmerge_io_stream_in_105_bits),
    .io_stream_in_106_ready(rmerge_io_stream_in_106_ready),
    .io_stream_in_106_valid(rmerge_io_stream_in_106_valid),
    .io_stream_in_106_bits(rmerge_io_stream_in_106_bits),
    .io_stream_in_107_ready(rmerge_io_stream_in_107_ready),
    .io_stream_in_107_valid(rmerge_io_stream_in_107_valid),
    .io_stream_in_107_bits(rmerge_io_stream_in_107_bits),
    .io_stream_in_108_ready(rmerge_io_stream_in_108_ready),
    .io_stream_in_108_valid(rmerge_io_stream_in_108_valid),
    .io_stream_in_108_bits(rmerge_io_stream_in_108_bits),
    .io_stream_in_109_ready(rmerge_io_stream_in_109_ready),
    .io_stream_in_109_valid(rmerge_io_stream_in_109_valid),
    .io_stream_in_109_bits(rmerge_io_stream_in_109_bits),
    .io_stream_in_110_ready(rmerge_io_stream_in_110_ready),
    .io_stream_in_110_valid(rmerge_io_stream_in_110_valid),
    .io_stream_in_110_bits(rmerge_io_stream_in_110_bits),
    .io_stream_in_111_ready(rmerge_io_stream_in_111_ready),
    .io_stream_in_111_valid(rmerge_io_stream_in_111_valid),
    .io_stream_in_111_bits(rmerge_io_stream_in_111_bits),
    .io_stream_in_112_ready(rmerge_io_stream_in_112_ready),
    .io_stream_in_112_valid(rmerge_io_stream_in_112_valid),
    .io_stream_in_112_bits(rmerge_io_stream_in_112_bits),
    .io_stream_in_113_ready(rmerge_io_stream_in_113_ready),
    .io_stream_in_113_valid(rmerge_io_stream_in_113_valid),
    .io_stream_in_113_bits(rmerge_io_stream_in_113_bits),
    .io_stream_in_114_ready(rmerge_io_stream_in_114_ready),
    .io_stream_in_114_valid(rmerge_io_stream_in_114_valid),
    .io_stream_in_114_bits(rmerge_io_stream_in_114_bits),
    .io_stream_in_115_ready(rmerge_io_stream_in_115_ready),
    .io_stream_in_115_valid(rmerge_io_stream_in_115_valid),
    .io_stream_in_115_bits(rmerge_io_stream_in_115_bits),
    .io_stream_in_116_ready(rmerge_io_stream_in_116_ready),
    .io_stream_in_116_valid(rmerge_io_stream_in_116_valid),
    .io_stream_in_116_bits(rmerge_io_stream_in_116_bits),
    .io_stream_in_117_ready(rmerge_io_stream_in_117_ready),
    .io_stream_in_117_valid(rmerge_io_stream_in_117_valid),
    .io_stream_in_117_bits(rmerge_io_stream_in_117_bits),
    .io_stream_in_118_ready(rmerge_io_stream_in_118_ready),
    .io_stream_in_118_valid(rmerge_io_stream_in_118_valid),
    .io_stream_in_118_bits(rmerge_io_stream_in_118_bits),
    .io_stream_in_119_ready(rmerge_io_stream_in_119_ready),
    .io_stream_in_119_valid(rmerge_io_stream_in_119_valid),
    .io_stream_in_119_bits(rmerge_io_stream_in_119_bits),
    .io_stream_in_120_ready(rmerge_io_stream_in_120_ready),
    .io_stream_in_120_valid(rmerge_io_stream_in_120_valid),
    .io_stream_in_120_bits(rmerge_io_stream_in_120_bits),
    .io_stream_in_121_ready(rmerge_io_stream_in_121_ready),
    .io_stream_in_121_valid(rmerge_io_stream_in_121_valid),
    .io_stream_in_121_bits(rmerge_io_stream_in_121_bits),
    .io_stream_in_122_ready(rmerge_io_stream_in_122_ready),
    .io_stream_in_122_valid(rmerge_io_stream_in_122_valid),
    .io_stream_in_122_bits(rmerge_io_stream_in_122_bits),
    .io_stream_in_123_ready(rmerge_io_stream_in_123_ready),
    .io_stream_in_123_valid(rmerge_io_stream_in_123_valid),
    .io_stream_in_123_bits(rmerge_io_stream_in_123_bits),
    .io_stream_in_124_ready(rmerge_io_stream_in_124_ready),
    .io_stream_in_124_valid(rmerge_io_stream_in_124_valid),
    .io_stream_in_124_bits(rmerge_io_stream_in_124_bits),
    .io_stream_in_125_ready(rmerge_io_stream_in_125_ready),
    .io_stream_in_125_valid(rmerge_io_stream_in_125_valid),
    .io_stream_in_125_bits(rmerge_io_stream_in_125_bits),
    .io_stream_in_126_ready(rmerge_io_stream_in_126_ready),
    .io_stream_in_126_valid(rmerge_io_stream_in_126_valid),
    .io_stream_in_126_bits(rmerge_io_stream_in_126_bits),
    .io_stream_in_127_ready(rmerge_io_stream_in_127_ready),
    .io_stream_in_127_valid(rmerge_io_stream_in_127_valid),
    .io_stream_in_127_bits(rmerge_io_stream_in_127_bits),
    .io_stream_in_128_ready(rmerge_io_stream_in_128_ready),
    .io_stream_in_128_valid(rmerge_io_stream_in_128_valid),
    .io_stream_in_128_bits(rmerge_io_stream_in_128_bits),
    .io_stream_in_129_ready(rmerge_io_stream_in_129_ready),
    .io_stream_in_129_valid(rmerge_io_stream_in_129_valid),
    .io_stream_in_129_bits(rmerge_io_stream_in_129_bits),
    .io_stream_in_130_ready(rmerge_io_stream_in_130_ready),
    .io_stream_in_130_valid(rmerge_io_stream_in_130_valid),
    .io_stream_in_130_bits(rmerge_io_stream_in_130_bits),
    .io_stream_in_131_ready(rmerge_io_stream_in_131_ready),
    .io_stream_in_131_valid(rmerge_io_stream_in_131_valid),
    .io_stream_in_131_bits(rmerge_io_stream_in_131_bits),
    .io_stream_in_132_ready(rmerge_io_stream_in_132_ready),
    .io_stream_in_132_valid(rmerge_io_stream_in_132_valid),
    .io_stream_in_132_bits(rmerge_io_stream_in_132_bits),
    .io_stream_in_133_ready(rmerge_io_stream_in_133_ready),
    .io_stream_in_133_valid(rmerge_io_stream_in_133_valid),
    .io_stream_in_133_bits(rmerge_io_stream_in_133_bits),
    .io_stream_in_134_ready(rmerge_io_stream_in_134_ready),
    .io_stream_in_134_valid(rmerge_io_stream_in_134_valid),
    .io_stream_in_134_bits(rmerge_io_stream_in_134_bits),
    .io_stream_in_135_ready(rmerge_io_stream_in_135_ready),
    .io_stream_in_135_valid(rmerge_io_stream_in_135_valid),
    .io_stream_in_135_bits(rmerge_io_stream_in_135_bits),
    .io_stream_in_136_ready(rmerge_io_stream_in_136_ready),
    .io_stream_in_136_valid(rmerge_io_stream_in_136_valid),
    .io_stream_in_136_bits(rmerge_io_stream_in_136_bits),
    .io_stream_in_137_ready(rmerge_io_stream_in_137_ready),
    .io_stream_in_137_valid(rmerge_io_stream_in_137_valid),
    .io_stream_in_137_bits(rmerge_io_stream_in_137_bits),
    .io_stream_in_138_ready(rmerge_io_stream_in_138_ready),
    .io_stream_in_138_valid(rmerge_io_stream_in_138_valid),
    .io_stream_in_138_bits(rmerge_io_stream_in_138_bits),
    .io_stream_in_139_ready(rmerge_io_stream_in_139_ready),
    .io_stream_in_139_valid(rmerge_io_stream_in_139_valid),
    .io_stream_in_139_bits(rmerge_io_stream_in_139_bits),
    .io_stream_in_140_ready(rmerge_io_stream_in_140_ready),
    .io_stream_in_140_valid(rmerge_io_stream_in_140_valid),
    .io_stream_in_140_bits(rmerge_io_stream_in_140_bits),
    .io_stream_in_141_ready(rmerge_io_stream_in_141_ready),
    .io_stream_in_141_valid(rmerge_io_stream_in_141_valid),
    .io_stream_in_141_bits(rmerge_io_stream_in_141_bits),
    .io_stream_in_142_ready(rmerge_io_stream_in_142_ready),
    .io_stream_in_142_valid(rmerge_io_stream_in_142_valid),
    .io_stream_in_142_bits(rmerge_io_stream_in_142_bits),
    .io_stream_in_143_ready(rmerge_io_stream_in_143_ready),
    .io_stream_in_143_valid(rmerge_io_stream_in_143_valid),
    .io_stream_in_143_bits(rmerge_io_stream_in_143_bits),
    .io_stream_in_144_ready(rmerge_io_stream_in_144_ready),
    .io_stream_in_144_valid(rmerge_io_stream_in_144_valid),
    .io_stream_in_144_bits(rmerge_io_stream_in_144_bits),
    .io_stream_in_145_ready(rmerge_io_stream_in_145_ready),
    .io_stream_in_145_valid(rmerge_io_stream_in_145_valid),
    .io_stream_in_145_bits(rmerge_io_stream_in_145_bits),
    .io_stream_in_146_ready(rmerge_io_stream_in_146_ready),
    .io_stream_in_146_valid(rmerge_io_stream_in_146_valid),
    .io_stream_in_146_bits(rmerge_io_stream_in_146_bits),
    .io_stream_in_147_ready(rmerge_io_stream_in_147_ready),
    .io_stream_in_147_valid(rmerge_io_stream_in_147_valid),
    .io_stream_in_147_bits(rmerge_io_stream_in_147_bits),
    .io_stream_in_148_ready(rmerge_io_stream_in_148_ready),
    .io_stream_in_148_valid(rmerge_io_stream_in_148_valid),
    .io_stream_in_148_bits(rmerge_io_stream_in_148_bits),
    .io_stream_in_149_ready(rmerge_io_stream_in_149_ready),
    .io_stream_in_149_valid(rmerge_io_stream_in_149_valid),
    .io_stream_in_149_bits(rmerge_io_stream_in_149_bits),
    .io_stream_in_150_ready(rmerge_io_stream_in_150_ready),
    .io_stream_in_150_valid(rmerge_io_stream_in_150_valid),
    .io_stream_in_150_bits(rmerge_io_stream_in_150_bits),
    .io_stream_in_151_ready(rmerge_io_stream_in_151_ready),
    .io_stream_in_151_valid(rmerge_io_stream_in_151_valid),
    .io_stream_in_151_bits(rmerge_io_stream_in_151_bits),
    .io_stream_in_152_ready(rmerge_io_stream_in_152_ready),
    .io_stream_in_152_valid(rmerge_io_stream_in_152_valid),
    .io_stream_in_152_bits(rmerge_io_stream_in_152_bits),
    .io_stream_in_153_ready(rmerge_io_stream_in_153_ready),
    .io_stream_in_153_valid(rmerge_io_stream_in_153_valid),
    .io_stream_in_153_bits(rmerge_io_stream_in_153_bits),
    .io_stream_in_154_ready(rmerge_io_stream_in_154_ready),
    .io_stream_in_154_valid(rmerge_io_stream_in_154_valid),
    .io_stream_in_154_bits(rmerge_io_stream_in_154_bits),
    .io_stream_in_155_ready(rmerge_io_stream_in_155_ready),
    .io_stream_in_155_valid(rmerge_io_stream_in_155_valid),
    .io_stream_in_155_bits(rmerge_io_stream_in_155_bits),
    .io_stream_in_156_ready(rmerge_io_stream_in_156_ready),
    .io_stream_in_156_valid(rmerge_io_stream_in_156_valid),
    .io_stream_in_156_bits(rmerge_io_stream_in_156_bits),
    .io_stream_in_157_ready(rmerge_io_stream_in_157_ready),
    .io_stream_in_157_valid(rmerge_io_stream_in_157_valid),
    .io_stream_in_157_bits(rmerge_io_stream_in_157_bits),
    .io_stream_in_158_ready(rmerge_io_stream_in_158_ready),
    .io_stream_in_158_valid(rmerge_io_stream_in_158_valid),
    .io_stream_in_158_bits(rmerge_io_stream_in_158_bits),
    .io_stream_in_159_ready(rmerge_io_stream_in_159_ready),
    .io_stream_in_159_valid(rmerge_io_stream_in_159_valid),
    .io_stream_in_159_bits(rmerge_io_stream_in_159_bits),
    .io_stream_in_160_ready(rmerge_io_stream_in_160_ready),
    .io_stream_in_160_valid(rmerge_io_stream_in_160_valid),
    .io_stream_in_160_bits(rmerge_io_stream_in_160_bits),
    .io_stream_in_161_ready(rmerge_io_stream_in_161_ready),
    .io_stream_in_161_valid(rmerge_io_stream_in_161_valid),
    .io_stream_in_161_bits(rmerge_io_stream_in_161_bits),
    .io_stream_in_162_ready(rmerge_io_stream_in_162_ready),
    .io_stream_in_162_valid(rmerge_io_stream_in_162_valid),
    .io_stream_in_162_bits(rmerge_io_stream_in_162_bits),
    .io_stream_in_163_ready(rmerge_io_stream_in_163_ready),
    .io_stream_in_163_valid(rmerge_io_stream_in_163_valid),
    .io_stream_in_163_bits(rmerge_io_stream_in_163_bits),
    .io_stream_in_164_ready(rmerge_io_stream_in_164_ready),
    .io_stream_in_164_valid(rmerge_io_stream_in_164_valid),
    .io_stream_in_164_bits(rmerge_io_stream_in_164_bits),
    .io_stream_in_165_ready(rmerge_io_stream_in_165_ready),
    .io_stream_in_165_valid(rmerge_io_stream_in_165_valid),
    .io_stream_in_165_bits(rmerge_io_stream_in_165_bits),
    .io_stream_in_166_ready(rmerge_io_stream_in_166_ready),
    .io_stream_in_166_valid(rmerge_io_stream_in_166_valid),
    .io_stream_in_166_bits(rmerge_io_stream_in_166_bits),
    .io_stream_in_167_ready(rmerge_io_stream_in_167_ready),
    .io_stream_in_167_valid(rmerge_io_stream_in_167_valid),
    .io_stream_in_167_bits(rmerge_io_stream_in_167_bits),
    .io_stream_in_168_ready(rmerge_io_stream_in_168_ready),
    .io_stream_in_168_valid(rmerge_io_stream_in_168_valid),
    .io_stream_in_168_bits(rmerge_io_stream_in_168_bits),
    .io_stream_in_169_ready(rmerge_io_stream_in_169_ready),
    .io_stream_in_169_valid(rmerge_io_stream_in_169_valid),
    .io_stream_in_169_bits(rmerge_io_stream_in_169_bits),
    .io_stream_in_170_ready(rmerge_io_stream_in_170_ready),
    .io_stream_in_170_valid(rmerge_io_stream_in_170_valid),
    .io_stream_in_170_bits(rmerge_io_stream_in_170_bits),
    .io_stream_in_171_ready(rmerge_io_stream_in_171_ready),
    .io_stream_in_171_valid(rmerge_io_stream_in_171_valid),
    .io_stream_in_171_bits(rmerge_io_stream_in_171_bits),
    .io_stream_in_172_ready(rmerge_io_stream_in_172_ready),
    .io_stream_in_172_valid(rmerge_io_stream_in_172_valid),
    .io_stream_in_172_bits(rmerge_io_stream_in_172_bits),
    .io_stream_in_173_ready(rmerge_io_stream_in_173_ready),
    .io_stream_in_173_valid(rmerge_io_stream_in_173_valid),
    .io_stream_in_173_bits(rmerge_io_stream_in_173_bits),
    .io_stream_in_174_ready(rmerge_io_stream_in_174_ready),
    .io_stream_in_174_valid(rmerge_io_stream_in_174_valid),
    .io_stream_in_174_bits(rmerge_io_stream_in_174_bits),
    .io_stream_in_175_ready(rmerge_io_stream_in_175_ready),
    .io_stream_in_175_valid(rmerge_io_stream_in_175_valid),
    .io_stream_in_175_bits(rmerge_io_stream_in_175_bits),
    .io_stream_in_176_ready(rmerge_io_stream_in_176_ready),
    .io_stream_in_176_valid(rmerge_io_stream_in_176_valid),
    .io_stream_in_176_bits(rmerge_io_stream_in_176_bits),
    .io_stream_in_177_ready(rmerge_io_stream_in_177_ready),
    .io_stream_in_177_valid(rmerge_io_stream_in_177_valid),
    .io_stream_in_177_bits(rmerge_io_stream_in_177_bits),
    .io_stream_in_178_ready(rmerge_io_stream_in_178_ready),
    .io_stream_in_178_valid(rmerge_io_stream_in_178_valid),
    .io_stream_in_178_bits(rmerge_io_stream_in_178_bits),
    .io_stream_in_179_ready(rmerge_io_stream_in_179_ready),
    .io_stream_in_179_valid(rmerge_io_stream_in_179_valid),
    .io_stream_in_179_bits(rmerge_io_stream_in_179_bits),
    .io_stream_in_180_ready(rmerge_io_stream_in_180_ready),
    .io_stream_in_180_valid(rmerge_io_stream_in_180_valid),
    .io_stream_in_180_bits(rmerge_io_stream_in_180_bits),
    .io_stream_in_181_ready(rmerge_io_stream_in_181_ready),
    .io_stream_in_181_valid(rmerge_io_stream_in_181_valid),
    .io_stream_in_181_bits(rmerge_io_stream_in_181_bits),
    .io_stream_in_182_ready(rmerge_io_stream_in_182_ready),
    .io_stream_in_182_valid(rmerge_io_stream_in_182_valid),
    .io_stream_in_182_bits(rmerge_io_stream_in_182_bits),
    .io_stream_in_183_ready(rmerge_io_stream_in_183_ready),
    .io_stream_in_183_valid(rmerge_io_stream_in_183_valid),
    .io_stream_in_183_bits(rmerge_io_stream_in_183_bits),
    .io_stream_in_184_ready(rmerge_io_stream_in_184_ready),
    .io_stream_in_184_valid(rmerge_io_stream_in_184_valid),
    .io_stream_in_184_bits(rmerge_io_stream_in_184_bits),
    .io_stream_in_185_ready(rmerge_io_stream_in_185_ready),
    .io_stream_in_185_valid(rmerge_io_stream_in_185_valid),
    .io_stream_in_185_bits(rmerge_io_stream_in_185_bits),
    .io_stream_in_186_ready(rmerge_io_stream_in_186_ready),
    .io_stream_in_186_valid(rmerge_io_stream_in_186_valid),
    .io_stream_in_186_bits(rmerge_io_stream_in_186_bits),
    .io_stream_in_187_ready(rmerge_io_stream_in_187_ready),
    .io_stream_in_187_valid(rmerge_io_stream_in_187_valid),
    .io_stream_in_187_bits(rmerge_io_stream_in_187_bits),
    .io_stream_in_188_ready(rmerge_io_stream_in_188_ready),
    .io_stream_in_188_valid(rmerge_io_stream_in_188_valid),
    .io_stream_in_188_bits(rmerge_io_stream_in_188_bits),
    .io_stream_in_189_ready(rmerge_io_stream_in_189_ready),
    .io_stream_in_189_valid(rmerge_io_stream_in_189_valid),
    .io_stream_in_189_bits(rmerge_io_stream_in_189_bits),
    .io_stream_in_190_ready(rmerge_io_stream_in_190_ready),
    .io_stream_in_190_valid(rmerge_io_stream_in_190_valid),
    .io_stream_in_190_bits(rmerge_io_stream_in_190_bits),
    .io_stream_in_191_ready(rmerge_io_stream_in_191_ready),
    .io_stream_in_191_valid(rmerge_io_stream_in_191_valid),
    .io_stream_in_191_bits(rmerge_io_stream_in_191_bits),
    .io_stream_in_192_ready(rmerge_io_stream_in_192_ready),
    .io_stream_in_192_valid(rmerge_io_stream_in_192_valid),
    .io_stream_in_192_bits(rmerge_io_stream_in_192_bits),
    .io_stream_in_193_ready(rmerge_io_stream_in_193_ready),
    .io_stream_in_193_valid(rmerge_io_stream_in_193_valid),
    .io_stream_in_193_bits(rmerge_io_stream_in_193_bits),
    .io_stream_in_194_ready(rmerge_io_stream_in_194_ready),
    .io_stream_in_194_valid(rmerge_io_stream_in_194_valid),
    .io_stream_in_194_bits(rmerge_io_stream_in_194_bits),
    .io_stream_in_195_ready(rmerge_io_stream_in_195_ready),
    .io_stream_in_195_valid(rmerge_io_stream_in_195_valid),
    .io_stream_in_195_bits(rmerge_io_stream_in_195_bits),
    .io_stream_in_196_ready(rmerge_io_stream_in_196_ready),
    .io_stream_in_196_valid(rmerge_io_stream_in_196_valid),
    .io_stream_in_196_bits(rmerge_io_stream_in_196_bits),
    .io_stream_in_197_ready(rmerge_io_stream_in_197_ready),
    .io_stream_in_197_valid(rmerge_io_stream_in_197_valid),
    .io_stream_in_197_bits(rmerge_io_stream_in_197_bits),
    .io_stream_in_198_ready(rmerge_io_stream_in_198_ready),
    .io_stream_in_198_valid(rmerge_io_stream_in_198_valid),
    .io_stream_in_198_bits(rmerge_io_stream_in_198_bits),
    .io_stream_in_199_ready(rmerge_io_stream_in_199_ready),
    .io_stream_in_199_valid(rmerge_io_stream_in_199_valid),
    .io_stream_in_199_bits(rmerge_io_stream_in_199_bits),
    .io_stream_in_200_ready(rmerge_io_stream_in_200_ready),
    .io_stream_in_200_valid(rmerge_io_stream_in_200_valid),
    .io_stream_in_200_bits(rmerge_io_stream_in_200_bits),
    .io_stream_in_201_ready(rmerge_io_stream_in_201_ready),
    .io_stream_in_201_valid(rmerge_io_stream_in_201_valid),
    .io_stream_in_201_bits(rmerge_io_stream_in_201_bits),
    .io_stream_in_202_ready(rmerge_io_stream_in_202_ready),
    .io_stream_in_202_valid(rmerge_io_stream_in_202_valid),
    .io_stream_in_202_bits(rmerge_io_stream_in_202_bits),
    .io_stream_in_203_ready(rmerge_io_stream_in_203_ready),
    .io_stream_in_203_valid(rmerge_io_stream_in_203_valid),
    .io_stream_in_203_bits(rmerge_io_stream_in_203_bits),
    .io_stream_in_204_ready(rmerge_io_stream_in_204_ready),
    .io_stream_in_204_valid(rmerge_io_stream_in_204_valid),
    .io_stream_in_204_bits(rmerge_io_stream_in_204_bits),
    .io_stream_in_205_ready(rmerge_io_stream_in_205_ready),
    .io_stream_in_205_valid(rmerge_io_stream_in_205_valid),
    .io_stream_in_205_bits(rmerge_io_stream_in_205_bits),
    .io_stream_in_206_ready(rmerge_io_stream_in_206_ready),
    .io_stream_in_206_valid(rmerge_io_stream_in_206_valid),
    .io_stream_in_206_bits(rmerge_io_stream_in_206_bits),
    .io_stream_in_207_ready(rmerge_io_stream_in_207_ready),
    .io_stream_in_207_valid(rmerge_io_stream_in_207_valid),
    .io_stream_in_207_bits(rmerge_io_stream_in_207_bits),
    .io_stream_in_208_ready(rmerge_io_stream_in_208_ready),
    .io_stream_in_208_valid(rmerge_io_stream_in_208_valid),
    .io_stream_in_208_bits(rmerge_io_stream_in_208_bits),
    .io_stream_in_209_ready(rmerge_io_stream_in_209_ready),
    .io_stream_in_209_valid(rmerge_io_stream_in_209_valid),
    .io_stream_in_209_bits(rmerge_io_stream_in_209_bits),
    .io_stream_in_210_ready(rmerge_io_stream_in_210_ready),
    .io_stream_in_210_valid(rmerge_io_stream_in_210_valid),
    .io_stream_in_210_bits(rmerge_io_stream_in_210_bits),
    .io_stream_in_211_ready(rmerge_io_stream_in_211_ready),
    .io_stream_in_211_valid(rmerge_io_stream_in_211_valid),
    .io_stream_in_211_bits(rmerge_io_stream_in_211_bits),
    .io_stream_in_212_ready(rmerge_io_stream_in_212_ready),
    .io_stream_in_212_valid(rmerge_io_stream_in_212_valid),
    .io_stream_in_212_bits(rmerge_io_stream_in_212_bits),
    .io_stream_in_213_ready(rmerge_io_stream_in_213_ready),
    .io_stream_in_213_valid(rmerge_io_stream_in_213_valid),
    .io_stream_in_213_bits(rmerge_io_stream_in_213_bits),
    .io_stream_in_214_ready(rmerge_io_stream_in_214_ready),
    .io_stream_in_214_valid(rmerge_io_stream_in_214_valid),
    .io_stream_in_214_bits(rmerge_io_stream_in_214_bits),
    .io_stream_in_215_ready(rmerge_io_stream_in_215_ready),
    .io_stream_in_215_valid(rmerge_io_stream_in_215_valid),
    .io_stream_in_215_bits(rmerge_io_stream_in_215_bits),
    .io_stream_in_216_ready(rmerge_io_stream_in_216_ready),
    .io_stream_in_216_valid(rmerge_io_stream_in_216_valid),
    .io_stream_in_216_bits(rmerge_io_stream_in_216_bits),
    .io_stream_in_217_ready(rmerge_io_stream_in_217_ready),
    .io_stream_in_217_valid(rmerge_io_stream_in_217_valid),
    .io_stream_in_217_bits(rmerge_io_stream_in_217_bits),
    .io_stream_in_218_ready(rmerge_io_stream_in_218_ready),
    .io_stream_in_218_valid(rmerge_io_stream_in_218_valid),
    .io_stream_in_218_bits(rmerge_io_stream_in_218_bits),
    .io_stream_in_219_ready(rmerge_io_stream_in_219_ready),
    .io_stream_in_219_valid(rmerge_io_stream_in_219_valid),
    .io_stream_in_219_bits(rmerge_io_stream_in_219_bits),
    .io_stream_in_220_ready(rmerge_io_stream_in_220_ready),
    .io_stream_in_220_valid(rmerge_io_stream_in_220_valid),
    .io_stream_in_220_bits(rmerge_io_stream_in_220_bits),
    .io_stream_in_221_ready(rmerge_io_stream_in_221_ready),
    .io_stream_in_221_valid(rmerge_io_stream_in_221_valid),
    .io_stream_in_221_bits(rmerge_io_stream_in_221_bits),
    .io_stream_in_222_ready(rmerge_io_stream_in_222_ready),
    .io_stream_in_222_valid(rmerge_io_stream_in_222_valid),
    .io_stream_in_222_bits(rmerge_io_stream_in_222_bits),
    .io_stream_in_223_ready(rmerge_io_stream_in_223_ready),
    .io_stream_in_223_valid(rmerge_io_stream_in_223_valid),
    .io_stream_in_223_bits(rmerge_io_stream_in_223_bits),
    .io_stream_in_224_ready(rmerge_io_stream_in_224_ready),
    .io_stream_in_224_valid(rmerge_io_stream_in_224_valid),
    .io_stream_in_224_bits(rmerge_io_stream_in_224_bits),
    .io_stream_in_225_ready(rmerge_io_stream_in_225_ready),
    .io_stream_in_225_valid(rmerge_io_stream_in_225_valid),
    .io_stream_in_225_bits(rmerge_io_stream_in_225_bits),
    .io_stream_in_226_ready(rmerge_io_stream_in_226_ready),
    .io_stream_in_226_valid(rmerge_io_stream_in_226_valid),
    .io_stream_in_226_bits(rmerge_io_stream_in_226_bits),
    .io_stream_in_227_ready(rmerge_io_stream_in_227_ready),
    .io_stream_in_227_valid(rmerge_io_stream_in_227_valid),
    .io_stream_in_227_bits(rmerge_io_stream_in_227_bits),
    .io_stream_in_228_ready(rmerge_io_stream_in_228_ready),
    .io_stream_in_228_valid(rmerge_io_stream_in_228_valid),
    .io_stream_in_228_bits(rmerge_io_stream_in_228_bits),
    .io_stream_in_229_ready(rmerge_io_stream_in_229_ready),
    .io_stream_in_229_valid(rmerge_io_stream_in_229_valid),
    .io_stream_in_229_bits(rmerge_io_stream_in_229_bits),
    .io_stream_in_230_ready(rmerge_io_stream_in_230_ready),
    .io_stream_in_230_valid(rmerge_io_stream_in_230_valid),
    .io_stream_in_230_bits(rmerge_io_stream_in_230_bits),
    .io_stream_in_231_ready(rmerge_io_stream_in_231_ready),
    .io_stream_in_231_valid(rmerge_io_stream_in_231_valid),
    .io_stream_in_231_bits(rmerge_io_stream_in_231_bits),
    .io_stream_in_232_ready(rmerge_io_stream_in_232_ready),
    .io_stream_in_232_valid(rmerge_io_stream_in_232_valid),
    .io_stream_in_232_bits(rmerge_io_stream_in_232_bits),
    .io_stream_in_233_ready(rmerge_io_stream_in_233_ready),
    .io_stream_in_233_valid(rmerge_io_stream_in_233_valid),
    .io_stream_in_233_bits(rmerge_io_stream_in_233_bits),
    .io_stream_in_234_ready(rmerge_io_stream_in_234_ready),
    .io_stream_in_234_valid(rmerge_io_stream_in_234_valid),
    .io_stream_in_234_bits(rmerge_io_stream_in_234_bits),
    .io_stream_in_235_ready(rmerge_io_stream_in_235_ready),
    .io_stream_in_235_valid(rmerge_io_stream_in_235_valid),
    .io_stream_in_235_bits(rmerge_io_stream_in_235_bits),
    .io_stream_in_236_ready(rmerge_io_stream_in_236_ready),
    .io_stream_in_236_valid(rmerge_io_stream_in_236_valid),
    .io_stream_in_236_bits(rmerge_io_stream_in_236_bits),
    .io_stream_in_237_ready(rmerge_io_stream_in_237_ready),
    .io_stream_in_237_valid(rmerge_io_stream_in_237_valid),
    .io_stream_in_237_bits(rmerge_io_stream_in_237_bits),
    .io_stream_in_238_ready(rmerge_io_stream_in_238_ready),
    .io_stream_in_238_valid(rmerge_io_stream_in_238_valid),
    .io_stream_in_238_bits(rmerge_io_stream_in_238_bits),
    .io_stream_in_239_ready(rmerge_io_stream_in_239_ready),
    .io_stream_in_239_valid(rmerge_io_stream_in_239_valid),
    .io_stream_in_239_bits(rmerge_io_stream_in_239_bits),
    .io_stream_in_240_ready(rmerge_io_stream_in_240_ready),
    .io_stream_in_240_valid(rmerge_io_stream_in_240_valid),
    .io_stream_in_240_bits(rmerge_io_stream_in_240_bits),
    .io_stream_in_241_ready(rmerge_io_stream_in_241_ready),
    .io_stream_in_241_valid(rmerge_io_stream_in_241_valid),
    .io_stream_in_241_bits(rmerge_io_stream_in_241_bits),
    .io_stream_in_242_ready(rmerge_io_stream_in_242_ready),
    .io_stream_in_242_valid(rmerge_io_stream_in_242_valid),
    .io_stream_in_242_bits(rmerge_io_stream_in_242_bits),
    .io_stream_in_243_ready(rmerge_io_stream_in_243_ready),
    .io_stream_in_243_valid(rmerge_io_stream_in_243_valid),
    .io_stream_in_243_bits(rmerge_io_stream_in_243_bits),
    .io_stream_in_244_ready(rmerge_io_stream_in_244_ready),
    .io_stream_in_244_valid(rmerge_io_stream_in_244_valid),
    .io_stream_in_244_bits(rmerge_io_stream_in_244_bits),
    .io_stream_in_245_ready(rmerge_io_stream_in_245_ready),
    .io_stream_in_245_valid(rmerge_io_stream_in_245_valid),
    .io_stream_in_245_bits(rmerge_io_stream_in_245_bits),
    .io_stream_in_246_ready(rmerge_io_stream_in_246_ready),
    .io_stream_in_246_valid(rmerge_io_stream_in_246_valid),
    .io_stream_in_246_bits(rmerge_io_stream_in_246_bits),
    .io_stream_in_247_ready(rmerge_io_stream_in_247_ready),
    .io_stream_in_247_valid(rmerge_io_stream_in_247_valid),
    .io_stream_in_247_bits(rmerge_io_stream_in_247_bits),
    .io_stream_in_248_ready(rmerge_io_stream_in_248_ready),
    .io_stream_in_248_valid(rmerge_io_stream_in_248_valid),
    .io_stream_in_248_bits(rmerge_io_stream_in_248_bits),
    .io_stream_in_249_ready(rmerge_io_stream_in_249_ready),
    .io_stream_in_249_valid(rmerge_io_stream_in_249_valid),
    .io_stream_in_249_bits(rmerge_io_stream_in_249_bits),
    .io_stream_in_250_ready(rmerge_io_stream_in_250_ready),
    .io_stream_in_250_valid(rmerge_io_stream_in_250_valid),
    .io_stream_in_250_bits(rmerge_io_stream_in_250_bits),
    .io_stream_in_251_ready(rmerge_io_stream_in_251_ready),
    .io_stream_in_251_valid(rmerge_io_stream_in_251_valid),
    .io_stream_in_251_bits(rmerge_io_stream_in_251_bits),
    .io_stream_in_252_ready(rmerge_io_stream_in_252_ready),
    .io_stream_in_252_valid(rmerge_io_stream_in_252_valid),
    .io_stream_in_252_bits(rmerge_io_stream_in_252_bits),
    .io_stream_in_253_ready(rmerge_io_stream_in_253_ready),
    .io_stream_in_253_valid(rmerge_io_stream_in_253_valid),
    .io_stream_in_253_bits(rmerge_io_stream_in_253_bits),
    .io_stream_in_254_ready(rmerge_io_stream_in_254_ready),
    .io_stream_in_254_valid(rmerge_io_stream_in_254_valid),
    .io_stream_in_254_bits(rmerge_io_stream_in_254_bits),
    .io_stream_in_255_ready(rmerge_io_stream_in_255_ready),
    .io_stream_in_255_valid(rmerge_io_stream_in_255_valid),
    .io_stream_in_255_bits(rmerge_io_stream_in_255_bits),
    .io_stream_out_ready(rmerge_io_stream_out_ready),
    .io_stream_out_valid(rmerge_io_stream_out_valid),
    .io_stream_out_bits(rmerge_io_stream_out_bits)
  );
  assign io_value_in_ready = vsplit_io_stream_in_ready; // @[Stab.scala 319:15]
  assign io_weight_in_ready = wsplit_io_stream_in_ready; // @[Stab.scala 320:16]
  assign io_value_out_valid = rmerge_io_stream_out_valid; // @[Stab.scala 326:16]
  assign io_value_out_bits = rmerge_io_stream_out_bits; // @[Stab.scala 326:16]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_weight_in_0_valid = wsplit_io_stream_out_0_valid; // @[Stab.scala 322:24]
  assign core_io_weight_in_0_bits = wsplit_io_stream_out_0_bits; // @[Stab.scala 322:24]
  assign core_io_weight_in_1_valid = wsplit_io_stream_out_1_valid; // @[Stab.scala 322:24]
  assign core_io_weight_in_1_bits = wsplit_io_stream_out_1_bits; // @[Stab.scala 322:24]
  assign core_io_weight_in_2_valid = wsplit_io_stream_out_2_valid; // @[Stab.scala 322:24]
  assign core_io_weight_in_2_bits = wsplit_io_stream_out_2_bits; // @[Stab.scala 322:24]
  assign core_io_weight_in_3_valid = wsplit_io_stream_out_3_valid; // @[Stab.scala 322:24]
  assign core_io_weight_in_3_bits = wsplit_io_stream_out_3_bits; // @[Stab.scala 322:24]
  assign core_io_weight_in_4_valid = wsplit_io_stream_out_4_valid; // @[Stab.scala 322:24]
  assign core_io_weight_in_4_bits = wsplit_io_stream_out_4_bits; // @[Stab.scala 322:24]
  assign core_io_weight_in_5_valid = wsplit_io_stream_out_5_valid; // @[Stab.scala 322:24]
  assign core_io_weight_in_5_bits = wsplit_io_stream_out_5_bits; // @[Stab.scala 322:24]
  assign core_io_weight_in_6_valid = wsplit_io_stream_out_6_valid; // @[Stab.scala 322:24]
  assign core_io_weight_in_6_bits = wsplit_io_stream_out_6_bits; // @[Stab.scala 322:24]
  assign core_io_weight_in_7_valid = wsplit_io_stream_out_7_valid; // @[Stab.scala 322:24]
  assign core_io_weight_in_7_bits = wsplit_io_stream_out_7_bits; // @[Stab.scala 322:24]
  assign core_io_weight_in_8_valid = wsplit_io_stream_out_8_valid; // @[Stab.scala 322:24]
  assign core_io_weight_in_8_bits = wsplit_io_stream_out_8_bits; // @[Stab.scala 322:24]
  assign core_io_weight_in_9_valid = wsplit_io_stream_out_9_valid; // @[Stab.scala 322:24]
  assign core_io_weight_in_9_bits = wsplit_io_stream_out_9_bits; // @[Stab.scala 322:24]
  assign core_io_weight_in_10_valid = wsplit_io_stream_out_10_valid; // @[Stab.scala 322:24]
  assign core_io_weight_in_10_bits = wsplit_io_stream_out_10_bits; // @[Stab.scala 322:24]
  assign core_io_weight_in_11_valid = wsplit_io_stream_out_11_valid; // @[Stab.scala 322:24]
  assign core_io_weight_in_11_bits = wsplit_io_stream_out_11_bits; // @[Stab.scala 322:24]
  assign core_io_weight_in_12_valid = wsplit_io_stream_out_12_valid; // @[Stab.scala 322:24]
  assign core_io_weight_in_12_bits = wsplit_io_stream_out_12_bits; // @[Stab.scala 322:24]
  assign core_io_weight_in_13_valid = wsplit_io_stream_out_13_valid; // @[Stab.scala 322:24]
  assign core_io_weight_in_13_bits = wsplit_io_stream_out_13_bits; // @[Stab.scala 322:24]
  assign core_io_weight_in_14_valid = wsplit_io_stream_out_14_valid; // @[Stab.scala 322:24]
  assign core_io_weight_in_14_bits = wsplit_io_stream_out_14_bits; // @[Stab.scala 322:24]
  assign core_io_weight_in_15_valid = wsplit_io_stream_out_15_valid; // @[Stab.scala 322:24]
  assign core_io_weight_in_15_bits = wsplit_io_stream_out_15_bits; // @[Stab.scala 322:24]
  assign core_io_value_in_0_valid = vsplit_io_stream_out_0_valid; // @[Stab.scala 321:24]
  assign core_io_value_in_0_bits = vsplit_io_stream_out_0_bits; // @[Stab.scala 321:24]
  assign core_io_value_in_1_valid = vsplit_io_stream_out_1_valid; // @[Stab.scala 321:24]
  assign core_io_value_in_1_bits = vsplit_io_stream_out_1_bits; // @[Stab.scala 321:24]
  assign core_io_value_in_2_valid = vsplit_io_stream_out_2_valid; // @[Stab.scala 321:24]
  assign core_io_value_in_2_bits = vsplit_io_stream_out_2_bits; // @[Stab.scala 321:24]
  assign core_io_value_in_3_valid = vsplit_io_stream_out_3_valid; // @[Stab.scala 321:24]
  assign core_io_value_in_3_bits = vsplit_io_stream_out_3_bits; // @[Stab.scala 321:24]
  assign core_io_value_in_4_valid = vsplit_io_stream_out_4_valid; // @[Stab.scala 321:24]
  assign core_io_value_in_4_bits = vsplit_io_stream_out_4_bits; // @[Stab.scala 321:24]
  assign core_io_value_in_5_valid = vsplit_io_stream_out_5_valid; // @[Stab.scala 321:24]
  assign core_io_value_in_5_bits = vsplit_io_stream_out_5_bits; // @[Stab.scala 321:24]
  assign core_io_value_in_6_valid = vsplit_io_stream_out_6_valid; // @[Stab.scala 321:24]
  assign core_io_value_in_6_bits = vsplit_io_stream_out_6_bits; // @[Stab.scala 321:24]
  assign core_io_value_in_7_valid = vsplit_io_stream_out_7_valid; // @[Stab.scala 321:24]
  assign core_io_value_in_7_bits = vsplit_io_stream_out_7_bits; // @[Stab.scala 321:24]
  assign core_io_value_in_8_valid = vsplit_io_stream_out_8_valid; // @[Stab.scala 321:24]
  assign core_io_value_in_8_bits = vsplit_io_stream_out_8_bits; // @[Stab.scala 321:24]
  assign core_io_value_in_9_valid = vsplit_io_stream_out_9_valid; // @[Stab.scala 321:24]
  assign core_io_value_in_9_bits = vsplit_io_stream_out_9_bits; // @[Stab.scala 321:24]
  assign core_io_value_in_10_valid = vsplit_io_stream_out_10_valid; // @[Stab.scala 321:24]
  assign core_io_value_in_10_bits = vsplit_io_stream_out_10_bits; // @[Stab.scala 321:24]
  assign core_io_value_in_11_valid = vsplit_io_stream_out_11_valid; // @[Stab.scala 321:24]
  assign core_io_value_in_11_bits = vsplit_io_stream_out_11_bits; // @[Stab.scala 321:24]
  assign core_io_value_in_12_valid = vsplit_io_stream_out_12_valid; // @[Stab.scala 321:24]
  assign core_io_value_in_12_bits = vsplit_io_stream_out_12_bits; // @[Stab.scala 321:24]
  assign core_io_value_in_13_valid = vsplit_io_stream_out_13_valid; // @[Stab.scala 321:24]
  assign core_io_value_in_13_bits = vsplit_io_stream_out_13_bits; // @[Stab.scala 321:24]
  assign core_io_value_in_14_valid = vsplit_io_stream_out_14_valid; // @[Stab.scala 321:24]
  assign core_io_value_in_14_bits = vsplit_io_stream_out_14_bits; // @[Stab.scala 321:24]
  assign core_io_value_in_15_valid = vsplit_io_stream_out_15_valid; // @[Stab.scala 321:24]
  assign core_io_value_in_15_bits = vsplit_io_stream_out_15_bits; // @[Stab.scala 321:24]
  assign core_io_value_out_0_0_ready = rmerge_io_stream_in_0_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_0_1_ready = rmerge_io_stream_in_1_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_0_2_ready = rmerge_io_stream_in_2_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_0_3_ready = rmerge_io_stream_in_3_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_0_4_ready = rmerge_io_stream_in_4_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_0_5_ready = rmerge_io_stream_in_5_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_0_6_ready = rmerge_io_stream_in_6_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_0_7_ready = rmerge_io_stream_in_7_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_0_8_ready = rmerge_io_stream_in_8_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_0_9_ready = rmerge_io_stream_in_9_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_0_10_ready = rmerge_io_stream_in_10_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_0_11_ready = rmerge_io_stream_in_11_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_0_12_ready = rmerge_io_stream_in_12_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_0_13_ready = rmerge_io_stream_in_13_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_0_14_ready = rmerge_io_stream_in_14_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_0_15_ready = rmerge_io_stream_in_15_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_1_0_ready = rmerge_io_stream_in_16_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_1_1_ready = rmerge_io_stream_in_17_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_1_2_ready = rmerge_io_stream_in_18_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_1_3_ready = rmerge_io_stream_in_19_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_1_4_ready = rmerge_io_stream_in_20_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_1_5_ready = rmerge_io_stream_in_21_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_1_6_ready = rmerge_io_stream_in_22_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_1_7_ready = rmerge_io_stream_in_23_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_1_8_ready = rmerge_io_stream_in_24_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_1_9_ready = rmerge_io_stream_in_25_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_1_10_ready = rmerge_io_stream_in_26_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_1_11_ready = rmerge_io_stream_in_27_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_1_12_ready = rmerge_io_stream_in_28_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_1_13_ready = rmerge_io_stream_in_29_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_1_14_ready = rmerge_io_stream_in_30_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_1_15_ready = rmerge_io_stream_in_31_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_2_0_ready = rmerge_io_stream_in_32_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_2_1_ready = rmerge_io_stream_in_33_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_2_2_ready = rmerge_io_stream_in_34_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_2_3_ready = rmerge_io_stream_in_35_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_2_4_ready = rmerge_io_stream_in_36_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_2_5_ready = rmerge_io_stream_in_37_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_2_6_ready = rmerge_io_stream_in_38_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_2_7_ready = rmerge_io_stream_in_39_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_2_8_ready = rmerge_io_stream_in_40_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_2_9_ready = rmerge_io_stream_in_41_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_2_10_ready = rmerge_io_stream_in_42_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_2_11_ready = rmerge_io_stream_in_43_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_2_12_ready = rmerge_io_stream_in_44_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_2_13_ready = rmerge_io_stream_in_45_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_2_14_ready = rmerge_io_stream_in_46_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_2_15_ready = rmerge_io_stream_in_47_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_3_0_ready = rmerge_io_stream_in_48_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_3_1_ready = rmerge_io_stream_in_49_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_3_2_ready = rmerge_io_stream_in_50_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_3_3_ready = rmerge_io_stream_in_51_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_3_4_ready = rmerge_io_stream_in_52_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_3_5_ready = rmerge_io_stream_in_53_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_3_6_ready = rmerge_io_stream_in_54_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_3_7_ready = rmerge_io_stream_in_55_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_3_8_ready = rmerge_io_stream_in_56_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_3_9_ready = rmerge_io_stream_in_57_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_3_10_ready = rmerge_io_stream_in_58_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_3_11_ready = rmerge_io_stream_in_59_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_3_12_ready = rmerge_io_stream_in_60_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_3_13_ready = rmerge_io_stream_in_61_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_3_14_ready = rmerge_io_stream_in_62_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_3_15_ready = rmerge_io_stream_in_63_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_4_0_ready = rmerge_io_stream_in_64_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_4_1_ready = rmerge_io_stream_in_65_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_4_2_ready = rmerge_io_stream_in_66_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_4_3_ready = rmerge_io_stream_in_67_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_4_4_ready = rmerge_io_stream_in_68_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_4_5_ready = rmerge_io_stream_in_69_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_4_6_ready = rmerge_io_stream_in_70_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_4_7_ready = rmerge_io_stream_in_71_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_4_8_ready = rmerge_io_stream_in_72_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_4_9_ready = rmerge_io_stream_in_73_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_4_10_ready = rmerge_io_stream_in_74_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_4_11_ready = rmerge_io_stream_in_75_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_4_12_ready = rmerge_io_stream_in_76_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_4_13_ready = rmerge_io_stream_in_77_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_4_14_ready = rmerge_io_stream_in_78_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_4_15_ready = rmerge_io_stream_in_79_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_5_0_ready = rmerge_io_stream_in_80_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_5_1_ready = rmerge_io_stream_in_81_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_5_2_ready = rmerge_io_stream_in_82_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_5_3_ready = rmerge_io_stream_in_83_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_5_4_ready = rmerge_io_stream_in_84_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_5_5_ready = rmerge_io_stream_in_85_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_5_6_ready = rmerge_io_stream_in_86_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_5_7_ready = rmerge_io_stream_in_87_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_5_8_ready = rmerge_io_stream_in_88_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_5_9_ready = rmerge_io_stream_in_89_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_5_10_ready = rmerge_io_stream_in_90_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_5_11_ready = rmerge_io_stream_in_91_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_5_12_ready = rmerge_io_stream_in_92_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_5_13_ready = rmerge_io_stream_in_93_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_5_14_ready = rmerge_io_stream_in_94_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_5_15_ready = rmerge_io_stream_in_95_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_6_0_ready = rmerge_io_stream_in_96_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_6_1_ready = rmerge_io_stream_in_97_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_6_2_ready = rmerge_io_stream_in_98_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_6_3_ready = rmerge_io_stream_in_99_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_6_4_ready = rmerge_io_stream_in_100_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_6_5_ready = rmerge_io_stream_in_101_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_6_6_ready = rmerge_io_stream_in_102_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_6_7_ready = rmerge_io_stream_in_103_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_6_8_ready = rmerge_io_stream_in_104_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_6_9_ready = rmerge_io_stream_in_105_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_6_10_ready = rmerge_io_stream_in_106_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_6_11_ready = rmerge_io_stream_in_107_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_6_12_ready = rmerge_io_stream_in_108_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_6_13_ready = rmerge_io_stream_in_109_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_6_14_ready = rmerge_io_stream_in_110_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_6_15_ready = rmerge_io_stream_in_111_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_7_0_ready = rmerge_io_stream_in_112_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_7_1_ready = rmerge_io_stream_in_113_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_7_2_ready = rmerge_io_stream_in_114_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_7_3_ready = rmerge_io_stream_in_115_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_7_4_ready = rmerge_io_stream_in_116_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_7_5_ready = rmerge_io_stream_in_117_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_7_6_ready = rmerge_io_stream_in_118_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_7_7_ready = rmerge_io_stream_in_119_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_7_8_ready = rmerge_io_stream_in_120_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_7_9_ready = rmerge_io_stream_in_121_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_7_10_ready = rmerge_io_stream_in_122_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_7_11_ready = rmerge_io_stream_in_123_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_7_12_ready = rmerge_io_stream_in_124_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_7_13_ready = rmerge_io_stream_in_125_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_7_14_ready = rmerge_io_stream_in_126_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_7_15_ready = rmerge_io_stream_in_127_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_8_0_ready = rmerge_io_stream_in_128_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_8_1_ready = rmerge_io_stream_in_129_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_8_2_ready = rmerge_io_stream_in_130_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_8_3_ready = rmerge_io_stream_in_131_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_8_4_ready = rmerge_io_stream_in_132_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_8_5_ready = rmerge_io_stream_in_133_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_8_6_ready = rmerge_io_stream_in_134_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_8_7_ready = rmerge_io_stream_in_135_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_8_8_ready = rmerge_io_stream_in_136_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_8_9_ready = rmerge_io_stream_in_137_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_8_10_ready = rmerge_io_stream_in_138_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_8_11_ready = rmerge_io_stream_in_139_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_8_12_ready = rmerge_io_stream_in_140_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_8_13_ready = rmerge_io_stream_in_141_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_8_14_ready = rmerge_io_stream_in_142_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_8_15_ready = rmerge_io_stream_in_143_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_9_0_ready = rmerge_io_stream_in_144_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_9_1_ready = rmerge_io_stream_in_145_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_9_2_ready = rmerge_io_stream_in_146_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_9_3_ready = rmerge_io_stream_in_147_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_9_4_ready = rmerge_io_stream_in_148_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_9_5_ready = rmerge_io_stream_in_149_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_9_6_ready = rmerge_io_stream_in_150_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_9_7_ready = rmerge_io_stream_in_151_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_9_8_ready = rmerge_io_stream_in_152_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_9_9_ready = rmerge_io_stream_in_153_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_9_10_ready = rmerge_io_stream_in_154_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_9_11_ready = rmerge_io_stream_in_155_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_9_12_ready = rmerge_io_stream_in_156_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_9_13_ready = rmerge_io_stream_in_157_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_9_14_ready = rmerge_io_stream_in_158_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_9_15_ready = rmerge_io_stream_in_159_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_10_0_ready = rmerge_io_stream_in_160_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_10_1_ready = rmerge_io_stream_in_161_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_10_2_ready = rmerge_io_stream_in_162_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_10_3_ready = rmerge_io_stream_in_163_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_10_4_ready = rmerge_io_stream_in_164_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_10_5_ready = rmerge_io_stream_in_165_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_10_6_ready = rmerge_io_stream_in_166_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_10_7_ready = rmerge_io_stream_in_167_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_10_8_ready = rmerge_io_stream_in_168_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_10_9_ready = rmerge_io_stream_in_169_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_10_10_ready = rmerge_io_stream_in_170_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_10_11_ready = rmerge_io_stream_in_171_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_10_12_ready = rmerge_io_stream_in_172_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_10_13_ready = rmerge_io_stream_in_173_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_10_14_ready = rmerge_io_stream_in_174_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_10_15_ready = rmerge_io_stream_in_175_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_11_0_ready = rmerge_io_stream_in_176_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_11_1_ready = rmerge_io_stream_in_177_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_11_2_ready = rmerge_io_stream_in_178_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_11_3_ready = rmerge_io_stream_in_179_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_11_4_ready = rmerge_io_stream_in_180_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_11_5_ready = rmerge_io_stream_in_181_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_11_6_ready = rmerge_io_stream_in_182_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_11_7_ready = rmerge_io_stream_in_183_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_11_8_ready = rmerge_io_stream_in_184_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_11_9_ready = rmerge_io_stream_in_185_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_11_10_ready = rmerge_io_stream_in_186_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_11_11_ready = rmerge_io_stream_in_187_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_11_12_ready = rmerge_io_stream_in_188_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_11_13_ready = rmerge_io_stream_in_189_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_11_14_ready = rmerge_io_stream_in_190_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_11_15_ready = rmerge_io_stream_in_191_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_12_0_ready = rmerge_io_stream_in_192_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_12_1_ready = rmerge_io_stream_in_193_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_12_2_ready = rmerge_io_stream_in_194_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_12_3_ready = rmerge_io_stream_in_195_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_12_4_ready = rmerge_io_stream_in_196_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_12_5_ready = rmerge_io_stream_in_197_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_12_6_ready = rmerge_io_stream_in_198_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_12_7_ready = rmerge_io_stream_in_199_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_12_8_ready = rmerge_io_stream_in_200_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_12_9_ready = rmerge_io_stream_in_201_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_12_10_ready = rmerge_io_stream_in_202_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_12_11_ready = rmerge_io_stream_in_203_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_12_12_ready = rmerge_io_stream_in_204_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_12_13_ready = rmerge_io_stream_in_205_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_12_14_ready = rmerge_io_stream_in_206_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_12_15_ready = rmerge_io_stream_in_207_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_13_0_ready = rmerge_io_stream_in_208_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_13_1_ready = rmerge_io_stream_in_209_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_13_2_ready = rmerge_io_stream_in_210_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_13_3_ready = rmerge_io_stream_in_211_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_13_4_ready = rmerge_io_stream_in_212_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_13_5_ready = rmerge_io_stream_in_213_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_13_6_ready = rmerge_io_stream_in_214_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_13_7_ready = rmerge_io_stream_in_215_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_13_8_ready = rmerge_io_stream_in_216_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_13_9_ready = rmerge_io_stream_in_217_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_13_10_ready = rmerge_io_stream_in_218_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_13_11_ready = rmerge_io_stream_in_219_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_13_12_ready = rmerge_io_stream_in_220_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_13_13_ready = rmerge_io_stream_in_221_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_13_14_ready = rmerge_io_stream_in_222_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_13_15_ready = rmerge_io_stream_in_223_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_14_0_ready = rmerge_io_stream_in_224_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_14_1_ready = rmerge_io_stream_in_225_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_14_2_ready = rmerge_io_stream_in_226_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_14_3_ready = rmerge_io_stream_in_227_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_14_4_ready = rmerge_io_stream_in_228_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_14_5_ready = rmerge_io_stream_in_229_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_14_6_ready = rmerge_io_stream_in_230_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_14_7_ready = rmerge_io_stream_in_231_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_14_8_ready = rmerge_io_stream_in_232_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_14_9_ready = rmerge_io_stream_in_233_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_14_10_ready = rmerge_io_stream_in_234_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_14_11_ready = rmerge_io_stream_in_235_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_14_12_ready = rmerge_io_stream_in_236_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_14_13_ready = rmerge_io_stream_in_237_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_14_14_ready = rmerge_io_stream_in_238_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_14_15_ready = rmerge_io_stream_in_239_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_15_0_ready = rmerge_io_stream_in_240_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_15_1_ready = rmerge_io_stream_in_241_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_15_2_ready = rmerge_io_stream_in_242_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_15_3_ready = rmerge_io_stream_in_243_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_15_4_ready = rmerge_io_stream_in_244_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_15_5_ready = rmerge_io_stream_in_245_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_15_6_ready = rmerge_io_stream_in_246_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_15_7_ready = rmerge_io_stream_in_247_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_15_8_ready = rmerge_io_stream_in_248_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_15_9_ready = rmerge_io_stream_in_249_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_15_10_ready = rmerge_io_stream_in_250_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_15_11_ready = rmerge_io_stream_in_251_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_15_12_ready = rmerge_io_stream_in_252_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_15_13_ready = rmerge_io_stream_in_253_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_15_14_ready = rmerge_io_stream_in_254_ready; // @[Stab.scala 324:84]
  assign core_io_value_out_15_15_ready = rmerge_io_stream_in_255_ready; // @[Stab.scala 324:84]
  assign wsplit_clock = clock;
  assign wsplit_reset = reset;
  assign wsplit_io_stream_in_valid = io_weight_in_valid; // @[Stab.scala 320:16]
  assign wsplit_io_stream_in_bits = io_weight_in_bits; // @[Stab.scala 320:16]
  assign wsplit_io_stream_out_0_ready = core_io_weight_in_0_ready; // @[Stab.scala 322:24]
  assign wsplit_io_stream_out_1_ready = core_io_weight_in_1_ready; // @[Stab.scala 322:24]
  assign wsplit_io_stream_out_2_ready = core_io_weight_in_2_ready; // @[Stab.scala 322:24]
  assign wsplit_io_stream_out_3_ready = core_io_weight_in_3_ready; // @[Stab.scala 322:24]
  assign wsplit_io_stream_out_4_ready = core_io_weight_in_4_ready; // @[Stab.scala 322:24]
  assign wsplit_io_stream_out_5_ready = core_io_weight_in_5_ready; // @[Stab.scala 322:24]
  assign wsplit_io_stream_out_6_ready = core_io_weight_in_6_ready; // @[Stab.scala 322:24]
  assign wsplit_io_stream_out_7_ready = core_io_weight_in_7_ready; // @[Stab.scala 322:24]
  assign wsplit_io_stream_out_8_ready = core_io_weight_in_8_ready; // @[Stab.scala 322:24]
  assign wsplit_io_stream_out_9_ready = core_io_weight_in_9_ready; // @[Stab.scala 322:24]
  assign wsplit_io_stream_out_10_ready = core_io_weight_in_10_ready; // @[Stab.scala 322:24]
  assign wsplit_io_stream_out_11_ready = core_io_weight_in_11_ready; // @[Stab.scala 322:24]
  assign wsplit_io_stream_out_12_ready = core_io_weight_in_12_ready; // @[Stab.scala 322:24]
  assign wsplit_io_stream_out_13_ready = core_io_weight_in_13_ready; // @[Stab.scala 322:24]
  assign wsplit_io_stream_out_14_ready = core_io_weight_in_14_ready; // @[Stab.scala 322:24]
  assign wsplit_io_stream_out_15_ready = core_io_weight_in_15_ready; // @[Stab.scala 322:24]
  assign vsplit_clock = clock;
  assign vsplit_reset = reset;
  assign vsplit_io_stream_in_valid = io_value_in_valid; // @[Stab.scala 319:15]
  assign vsplit_io_stream_in_bits = io_value_in_bits; // @[Stab.scala 319:15]
  assign vsplit_io_stream_out_0_ready = core_io_value_in_0_ready; // @[Stab.scala 321:24]
  assign vsplit_io_stream_out_1_ready = core_io_value_in_1_ready; // @[Stab.scala 321:24]
  assign vsplit_io_stream_out_2_ready = core_io_value_in_2_ready; // @[Stab.scala 321:24]
  assign vsplit_io_stream_out_3_ready = core_io_value_in_3_ready; // @[Stab.scala 321:24]
  assign vsplit_io_stream_out_4_ready = core_io_value_in_4_ready; // @[Stab.scala 321:24]
  assign vsplit_io_stream_out_5_ready = core_io_value_in_5_ready; // @[Stab.scala 321:24]
  assign vsplit_io_stream_out_6_ready = core_io_value_in_6_ready; // @[Stab.scala 321:24]
  assign vsplit_io_stream_out_7_ready = core_io_value_in_7_ready; // @[Stab.scala 321:24]
  assign vsplit_io_stream_out_8_ready = core_io_value_in_8_ready; // @[Stab.scala 321:24]
  assign vsplit_io_stream_out_9_ready = core_io_value_in_9_ready; // @[Stab.scala 321:24]
  assign vsplit_io_stream_out_10_ready = core_io_value_in_10_ready; // @[Stab.scala 321:24]
  assign vsplit_io_stream_out_11_ready = core_io_value_in_11_ready; // @[Stab.scala 321:24]
  assign vsplit_io_stream_out_12_ready = core_io_value_in_12_ready; // @[Stab.scala 321:24]
  assign vsplit_io_stream_out_13_ready = core_io_value_in_13_ready; // @[Stab.scala 321:24]
  assign vsplit_io_stream_out_14_ready = core_io_value_in_14_ready; // @[Stab.scala 321:24]
  assign vsplit_io_stream_out_15_ready = core_io_value_in_15_ready; // @[Stab.scala 321:24]
  assign rmerge_clock = clock;
  assign rmerge_reset = reset;
  assign rmerge_io_stream_in_0_valid = core_io_value_out_0_0_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_0_bits = core_io_value_out_0_0_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_1_valid = core_io_value_out_0_1_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_1_bits = core_io_value_out_0_1_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_2_valid = core_io_value_out_0_2_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_2_bits = core_io_value_out_0_2_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_3_valid = core_io_value_out_0_3_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_3_bits = core_io_value_out_0_3_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_4_valid = core_io_value_out_0_4_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_4_bits = core_io_value_out_0_4_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_5_valid = core_io_value_out_0_5_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_5_bits = core_io_value_out_0_5_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_6_valid = core_io_value_out_0_6_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_6_bits = core_io_value_out_0_6_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_7_valid = core_io_value_out_0_7_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_7_bits = core_io_value_out_0_7_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_8_valid = core_io_value_out_0_8_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_8_bits = core_io_value_out_0_8_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_9_valid = core_io_value_out_0_9_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_9_bits = core_io_value_out_0_9_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_10_valid = core_io_value_out_0_10_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_10_bits = core_io_value_out_0_10_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_11_valid = core_io_value_out_0_11_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_11_bits = core_io_value_out_0_11_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_12_valid = core_io_value_out_0_12_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_12_bits = core_io_value_out_0_12_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_13_valid = core_io_value_out_0_13_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_13_bits = core_io_value_out_0_13_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_14_valid = core_io_value_out_0_14_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_14_bits = core_io_value_out_0_14_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_15_valid = core_io_value_out_0_15_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_15_bits = core_io_value_out_0_15_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_16_valid = core_io_value_out_1_0_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_16_bits = core_io_value_out_1_0_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_17_valid = core_io_value_out_1_1_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_17_bits = core_io_value_out_1_1_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_18_valid = core_io_value_out_1_2_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_18_bits = core_io_value_out_1_2_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_19_valid = core_io_value_out_1_3_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_19_bits = core_io_value_out_1_3_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_20_valid = core_io_value_out_1_4_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_20_bits = core_io_value_out_1_4_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_21_valid = core_io_value_out_1_5_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_21_bits = core_io_value_out_1_5_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_22_valid = core_io_value_out_1_6_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_22_bits = core_io_value_out_1_6_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_23_valid = core_io_value_out_1_7_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_23_bits = core_io_value_out_1_7_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_24_valid = core_io_value_out_1_8_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_24_bits = core_io_value_out_1_8_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_25_valid = core_io_value_out_1_9_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_25_bits = core_io_value_out_1_9_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_26_valid = core_io_value_out_1_10_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_26_bits = core_io_value_out_1_10_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_27_valid = core_io_value_out_1_11_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_27_bits = core_io_value_out_1_11_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_28_valid = core_io_value_out_1_12_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_28_bits = core_io_value_out_1_12_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_29_valid = core_io_value_out_1_13_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_29_bits = core_io_value_out_1_13_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_30_valid = core_io_value_out_1_14_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_30_bits = core_io_value_out_1_14_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_31_valid = core_io_value_out_1_15_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_31_bits = core_io_value_out_1_15_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_32_valid = core_io_value_out_2_0_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_32_bits = core_io_value_out_2_0_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_33_valid = core_io_value_out_2_1_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_33_bits = core_io_value_out_2_1_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_34_valid = core_io_value_out_2_2_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_34_bits = core_io_value_out_2_2_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_35_valid = core_io_value_out_2_3_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_35_bits = core_io_value_out_2_3_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_36_valid = core_io_value_out_2_4_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_36_bits = core_io_value_out_2_4_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_37_valid = core_io_value_out_2_5_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_37_bits = core_io_value_out_2_5_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_38_valid = core_io_value_out_2_6_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_38_bits = core_io_value_out_2_6_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_39_valid = core_io_value_out_2_7_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_39_bits = core_io_value_out_2_7_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_40_valid = core_io_value_out_2_8_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_40_bits = core_io_value_out_2_8_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_41_valid = core_io_value_out_2_9_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_41_bits = core_io_value_out_2_9_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_42_valid = core_io_value_out_2_10_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_42_bits = core_io_value_out_2_10_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_43_valid = core_io_value_out_2_11_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_43_bits = core_io_value_out_2_11_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_44_valid = core_io_value_out_2_12_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_44_bits = core_io_value_out_2_12_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_45_valid = core_io_value_out_2_13_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_45_bits = core_io_value_out_2_13_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_46_valid = core_io_value_out_2_14_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_46_bits = core_io_value_out_2_14_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_47_valid = core_io_value_out_2_15_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_47_bits = core_io_value_out_2_15_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_48_valid = core_io_value_out_3_0_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_48_bits = core_io_value_out_3_0_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_49_valid = core_io_value_out_3_1_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_49_bits = core_io_value_out_3_1_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_50_valid = core_io_value_out_3_2_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_50_bits = core_io_value_out_3_2_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_51_valid = core_io_value_out_3_3_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_51_bits = core_io_value_out_3_3_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_52_valid = core_io_value_out_3_4_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_52_bits = core_io_value_out_3_4_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_53_valid = core_io_value_out_3_5_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_53_bits = core_io_value_out_3_5_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_54_valid = core_io_value_out_3_6_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_54_bits = core_io_value_out_3_6_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_55_valid = core_io_value_out_3_7_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_55_bits = core_io_value_out_3_7_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_56_valid = core_io_value_out_3_8_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_56_bits = core_io_value_out_3_8_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_57_valid = core_io_value_out_3_9_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_57_bits = core_io_value_out_3_9_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_58_valid = core_io_value_out_3_10_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_58_bits = core_io_value_out_3_10_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_59_valid = core_io_value_out_3_11_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_59_bits = core_io_value_out_3_11_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_60_valid = core_io_value_out_3_12_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_60_bits = core_io_value_out_3_12_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_61_valid = core_io_value_out_3_13_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_61_bits = core_io_value_out_3_13_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_62_valid = core_io_value_out_3_14_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_62_bits = core_io_value_out_3_14_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_63_valid = core_io_value_out_3_15_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_63_bits = core_io_value_out_3_15_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_64_valid = core_io_value_out_4_0_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_64_bits = core_io_value_out_4_0_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_65_valid = core_io_value_out_4_1_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_65_bits = core_io_value_out_4_1_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_66_valid = core_io_value_out_4_2_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_66_bits = core_io_value_out_4_2_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_67_valid = core_io_value_out_4_3_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_67_bits = core_io_value_out_4_3_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_68_valid = core_io_value_out_4_4_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_68_bits = core_io_value_out_4_4_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_69_valid = core_io_value_out_4_5_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_69_bits = core_io_value_out_4_5_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_70_valid = core_io_value_out_4_6_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_70_bits = core_io_value_out_4_6_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_71_valid = core_io_value_out_4_7_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_71_bits = core_io_value_out_4_7_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_72_valid = core_io_value_out_4_8_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_72_bits = core_io_value_out_4_8_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_73_valid = core_io_value_out_4_9_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_73_bits = core_io_value_out_4_9_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_74_valid = core_io_value_out_4_10_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_74_bits = core_io_value_out_4_10_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_75_valid = core_io_value_out_4_11_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_75_bits = core_io_value_out_4_11_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_76_valid = core_io_value_out_4_12_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_76_bits = core_io_value_out_4_12_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_77_valid = core_io_value_out_4_13_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_77_bits = core_io_value_out_4_13_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_78_valid = core_io_value_out_4_14_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_78_bits = core_io_value_out_4_14_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_79_valid = core_io_value_out_4_15_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_79_bits = core_io_value_out_4_15_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_80_valid = core_io_value_out_5_0_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_80_bits = core_io_value_out_5_0_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_81_valid = core_io_value_out_5_1_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_81_bits = core_io_value_out_5_1_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_82_valid = core_io_value_out_5_2_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_82_bits = core_io_value_out_5_2_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_83_valid = core_io_value_out_5_3_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_83_bits = core_io_value_out_5_3_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_84_valid = core_io_value_out_5_4_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_84_bits = core_io_value_out_5_4_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_85_valid = core_io_value_out_5_5_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_85_bits = core_io_value_out_5_5_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_86_valid = core_io_value_out_5_6_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_86_bits = core_io_value_out_5_6_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_87_valid = core_io_value_out_5_7_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_87_bits = core_io_value_out_5_7_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_88_valid = core_io_value_out_5_8_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_88_bits = core_io_value_out_5_8_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_89_valid = core_io_value_out_5_9_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_89_bits = core_io_value_out_5_9_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_90_valid = core_io_value_out_5_10_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_90_bits = core_io_value_out_5_10_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_91_valid = core_io_value_out_5_11_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_91_bits = core_io_value_out_5_11_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_92_valid = core_io_value_out_5_12_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_92_bits = core_io_value_out_5_12_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_93_valid = core_io_value_out_5_13_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_93_bits = core_io_value_out_5_13_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_94_valid = core_io_value_out_5_14_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_94_bits = core_io_value_out_5_14_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_95_valid = core_io_value_out_5_15_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_95_bits = core_io_value_out_5_15_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_96_valid = core_io_value_out_6_0_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_96_bits = core_io_value_out_6_0_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_97_valid = core_io_value_out_6_1_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_97_bits = core_io_value_out_6_1_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_98_valid = core_io_value_out_6_2_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_98_bits = core_io_value_out_6_2_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_99_valid = core_io_value_out_6_3_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_99_bits = core_io_value_out_6_3_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_100_valid = core_io_value_out_6_4_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_100_bits = core_io_value_out_6_4_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_101_valid = core_io_value_out_6_5_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_101_bits = core_io_value_out_6_5_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_102_valid = core_io_value_out_6_6_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_102_bits = core_io_value_out_6_6_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_103_valid = core_io_value_out_6_7_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_103_bits = core_io_value_out_6_7_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_104_valid = core_io_value_out_6_8_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_104_bits = core_io_value_out_6_8_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_105_valid = core_io_value_out_6_9_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_105_bits = core_io_value_out_6_9_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_106_valid = core_io_value_out_6_10_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_106_bits = core_io_value_out_6_10_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_107_valid = core_io_value_out_6_11_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_107_bits = core_io_value_out_6_11_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_108_valid = core_io_value_out_6_12_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_108_bits = core_io_value_out_6_12_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_109_valid = core_io_value_out_6_13_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_109_bits = core_io_value_out_6_13_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_110_valid = core_io_value_out_6_14_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_110_bits = core_io_value_out_6_14_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_111_valid = core_io_value_out_6_15_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_111_bits = core_io_value_out_6_15_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_112_valid = core_io_value_out_7_0_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_112_bits = core_io_value_out_7_0_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_113_valid = core_io_value_out_7_1_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_113_bits = core_io_value_out_7_1_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_114_valid = core_io_value_out_7_2_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_114_bits = core_io_value_out_7_2_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_115_valid = core_io_value_out_7_3_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_115_bits = core_io_value_out_7_3_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_116_valid = core_io_value_out_7_4_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_116_bits = core_io_value_out_7_4_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_117_valid = core_io_value_out_7_5_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_117_bits = core_io_value_out_7_5_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_118_valid = core_io_value_out_7_6_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_118_bits = core_io_value_out_7_6_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_119_valid = core_io_value_out_7_7_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_119_bits = core_io_value_out_7_7_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_120_valid = core_io_value_out_7_8_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_120_bits = core_io_value_out_7_8_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_121_valid = core_io_value_out_7_9_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_121_bits = core_io_value_out_7_9_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_122_valid = core_io_value_out_7_10_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_122_bits = core_io_value_out_7_10_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_123_valid = core_io_value_out_7_11_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_123_bits = core_io_value_out_7_11_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_124_valid = core_io_value_out_7_12_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_124_bits = core_io_value_out_7_12_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_125_valid = core_io_value_out_7_13_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_125_bits = core_io_value_out_7_13_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_126_valid = core_io_value_out_7_14_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_126_bits = core_io_value_out_7_14_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_127_valid = core_io_value_out_7_15_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_127_bits = core_io_value_out_7_15_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_128_valid = core_io_value_out_8_0_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_128_bits = core_io_value_out_8_0_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_129_valid = core_io_value_out_8_1_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_129_bits = core_io_value_out_8_1_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_130_valid = core_io_value_out_8_2_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_130_bits = core_io_value_out_8_2_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_131_valid = core_io_value_out_8_3_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_131_bits = core_io_value_out_8_3_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_132_valid = core_io_value_out_8_4_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_132_bits = core_io_value_out_8_4_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_133_valid = core_io_value_out_8_5_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_133_bits = core_io_value_out_8_5_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_134_valid = core_io_value_out_8_6_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_134_bits = core_io_value_out_8_6_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_135_valid = core_io_value_out_8_7_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_135_bits = core_io_value_out_8_7_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_136_valid = core_io_value_out_8_8_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_136_bits = core_io_value_out_8_8_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_137_valid = core_io_value_out_8_9_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_137_bits = core_io_value_out_8_9_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_138_valid = core_io_value_out_8_10_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_138_bits = core_io_value_out_8_10_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_139_valid = core_io_value_out_8_11_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_139_bits = core_io_value_out_8_11_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_140_valid = core_io_value_out_8_12_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_140_bits = core_io_value_out_8_12_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_141_valid = core_io_value_out_8_13_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_141_bits = core_io_value_out_8_13_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_142_valid = core_io_value_out_8_14_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_142_bits = core_io_value_out_8_14_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_143_valid = core_io_value_out_8_15_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_143_bits = core_io_value_out_8_15_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_144_valid = core_io_value_out_9_0_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_144_bits = core_io_value_out_9_0_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_145_valid = core_io_value_out_9_1_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_145_bits = core_io_value_out_9_1_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_146_valid = core_io_value_out_9_2_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_146_bits = core_io_value_out_9_2_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_147_valid = core_io_value_out_9_3_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_147_bits = core_io_value_out_9_3_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_148_valid = core_io_value_out_9_4_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_148_bits = core_io_value_out_9_4_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_149_valid = core_io_value_out_9_5_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_149_bits = core_io_value_out_9_5_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_150_valid = core_io_value_out_9_6_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_150_bits = core_io_value_out_9_6_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_151_valid = core_io_value_out_9_7_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_151_bits = core_io_value_out_9_7_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_152_valid = core_io_value_out_9_8_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_152_bits = core_io_value_out_9_8_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_153_valid = core_io_value_out_9_9_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_153_bits = core_io_value_out_9_9_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_154_valid = core_io_value_out_9_10_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_154_bits = core_io_value_out_9_10_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_155_valid = core_io_value_out_9_11_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_155_bits = core_io_value_out_9_11_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_156_valid = core_io_value_out_9_12_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_156_bits = core_io_value_out_9_12_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_157_valid = core_io_value_out_9_13_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_157_bits = core_io_value_out_9_13_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_158_valid = core_io_value_out_9_14_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_158_bits = core_io_value_out_9_14_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_159_valid = core_io_value_out_9_15_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_159_bits = core_io_value_out_9_15_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_160_valid = core_io_value_out_10_0_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_160_bits = core_io_value_out_10_0_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_161_valid = core_io_value_out_10_1_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_161_bits = core_io_value_out_10_1_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_162_valid = core_io_value_out_10_2_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_162_bits = core_io_value_out_10_2_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_163_valid = core_io_value_out_10_3_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_163_bits = core_io_value_out_10_3_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_164_valid = core_io_value_out_10_4_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_164_bits = core_io_value_out_10_4_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_165_valid = core_io_value_out_10_5_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_165_bits = core_io_value_out_10_5_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_166_valid = core_io_value_out_10_6_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_166_bits = core_io_value_out_10_6_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_167_valid = core_io_value_out_10_7_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_167_bits = core_io_value_out_10_7_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_168_valid = core_io_value_out_10_8_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_168_bits = core_io_value_out_10_8_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_169_valid = core_io_value_out_10_9_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_169_bits = core_io_value_out_10_9_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_170_valid = core_io_value_out_10_10_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_170_bits = core_io_value_out_10_10_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_171_valid = core_io_value_out_10_11_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_171_bits = core_io_value_out_10_11_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_172_valid = core_io_value_out_10_12_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_172_bits = core_io_value_out_10_12_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_173_valid = core_io_value_out_10_13_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_173_bits = core_io_value_out_10_13_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_174_valid = core_io_value_out_10_14_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_174_bits = core_io_value_out_10_14_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_175_valid = core_io_value_out_10_15_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_175_bits = core_io_value_out_10_15_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_176_valid = core_io_value_out_11_0_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_176_bits = core_io_value_out_11_0_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_177_valid = core_io_value_out_11_1_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_177_bits = core_io_value_out_11_1_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_178_valid = core_io_value_out_11_2_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_178_bits = core_io_value_out_11_2_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_179_valid = core_io_value_out_11_3_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_179_bits = core_io_value_out_11_3_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_180_valid = core_io_value_out_11_4_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_180_bits = core_io_value_out_11_4_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_181_valid = core_io_value_out_11_5_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_181_bits = core_io_value_out_11_5_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_182_valid = core_io_value_out_11_6_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_182_bits = core_io_value_out_11_6_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_183_valid = core_io_value_out_11_7_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_183_bits = core_io_value_out_11_7_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_184_valid = core_io_value_out_11_8_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_184_bits = core_io_value_out_11_8_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_185_valid = core_io_value_out_11_9_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_185_bits = core_io_value_out_11_9_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_186_valid = core_io_value_out_11_10_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_186_bits = core_io_value_out_11_10_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_187_valid = core_io_value_out_11_11_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_187_bits = core_io_value_out_11_11_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_188_valid = core_io_value_out_11_12_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_188_bits = core_io_value_out_11_12_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_189_valid = core_io_value_out_11_13_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_189_bits = core_io_value_out_11_13_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_190_valid = core_io_value_out_11_14_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_190_bits = core_io_value_out_11_14_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_191_valid = core_io_value_out_11_15_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_191_bits = core_io_value_out_11_15_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_192_valid = core_io_value_out_12_0_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_192_bits = core_io_value_out_12_0_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_193_valid = core_io_value_out_12_1_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_193_bits = core_io_value_out_12_1_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_194_valid = core_io_value_out_12_2_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_194_bits = core_io_value_out_12_2_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_195_valid = core_io_value_out_12_3_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_195_bits = core_io_value_out_12_3_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_196_valid = core_io_value_out_12_4_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_196_bits = core_io_value_out_12_4_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_197_valid = core_io_value_out_12_5_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_197_bits = core_io_value_out_12_5_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_198_valid = core_io_value_out_12_6_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_198_bits = core_io_value_out_12_6_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_199_valid = core_io_value_out_12_7_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_199_bits = core_io_value_out_12_7_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_200_valid = core_io_value_out_12_8_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_200_bits = core_io_value_out_12_8_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_201_valid = core_io_value_out_12_9_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_201_bits = core_io_value_out_12_9_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_202_valid = core_io_value_out_12_10_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_202_bits = core_io_value_out_12_10_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_203_valid = core_io_value_out_12_11_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_203_bits = core_io_value_out_12_11_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_204_valid = core_io_value_out_12_12_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_204_bits = core_io_value_out_12_12_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_205_valid = core_io_value_out_12_13_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_205_bits = core_io_value_out_12_13_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_206_valid = core_io_value_out_12_14_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_206_bits = core_io_value_out_12_14_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_207_valid = core_io_value_out_12_15_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_207_bits = core_io_value_out_12_15_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_208_valid = core_io_value_out_13_0_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_208_bits = core_io_value_out_13_0_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_209_valid = core_io_value_out_13_1_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_209_bits = core_io_value_out_13_1_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_210_valid = core_io_value_out_13_2_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_210_bits = core_io_value_out_13_2_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_211_valid = core_io_value_out_13_3_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_211_bits = core_io_value_out_13_3_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_212_valid = core_io_value_out_13_4_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_212_bits = core_io_value_out_13_4_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_213_valid = core_io_value_out_13_5_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_213_bits = core_io_value_out_13_5_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_214_valid = core_io_value_out_13_6_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_214_bits = core_io_value_out_13_6_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_215_valid = core_io_value_out_13_7_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_215_bits = core_io_value_out_13_7_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_216_valid = core_io_value_out_13_8_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_216_bits = core_io_value_out_13_8_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_217_valid = core_io_value_out_13_9_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_217_bits = core_io_value_out_13_9_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_218_valid = core_io_value_out_13_10_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_218_bits = core_io_value_out_13_10_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_219_valid = core_io_value_out_13_11_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_219_bits = core_io_value_out_13_11_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_220_valid = core_io_value_out_13_12_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_220_bits = core_io_value_out_13_12_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_221_valid = core_io_value_out_13_13_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_221_bits = core_io_value_out_13_13_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_222_valid = core_io_value_out_13_14_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_222_bits = core_io_value_out_13_14_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_223_valid = core_io_value_out_13_15_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_223_bits = core_io_value_out_13_15_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_224_valid = core_io_value_out_14_0_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_224_bits = core_io_value_out_14_0_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_225_valid = core_io_value_out_14_1_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_225_bits = core_io_value_out_14_1_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_226_valid = core_io_value_out_14_2_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_226_bits = core_io_value_out_14_2_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_227_valid = core_io_value_out_14_3_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_227_bits = core_io_value_out_14_3_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_228_valid = core_io_value_out_14_4_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_228_bits = core_io_value_out_14_4_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_229_valid = core_io_value_out_14_5_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_229_bits = core_io_value_out_14_5_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_230_valid = core_io_value_out_14_6_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_230_bits = core_io_value_out_14_6_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_231_valid = core_io_value_out_14_7_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_231_bits = core_io_value_out_14_7_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_232_valid = core_io_value_out_14_8_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_232_bits = core_io_value_out_14_8_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_233_valid = core_io_value_out_14_9_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_233_bits = core_io_value_out_14_9_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_234_valid = core_io_value_out_14_10_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_234_bits = core_io_value_out_14_10_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_235_valid = core_io_value_out_14_11_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_235_bits = core_io_value_out_14_11_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_236_valid = core_io_value_out_14_12_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_236_bits = core_io_value_out_14_12_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_237_valid = core_io_value_out_14_13_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_237_bits = core_io_value_out_14_13_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_238_valid = core_io_value_out_14_14_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_238_bits = core_io_value_out_14_14_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_239_valid = core_io_value_out_14_15_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_239_bits = core_io_value_out_14_15_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_240_valid = core_io_value_out_15_0_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_240_bits = core_io_value_out_15_0_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_241_valid = core_io_value_out_15_1_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_241_bits = core_io_value_out_15_1_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_242_valid = core_io_value_out_15_2_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_242_bits = core_io_value_out_15_2_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_243_valid = core_io_value_out_15_3_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_243_bits = core_io_value_out_15_3_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_244_valid = core_io_value_out_15_4_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_244_bits = core_io_value_out_15_4_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_245_valid = core_io_value_out_15_5_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_245_bits = core_io_value_out_15_5_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_246_valid = core_io_value_out_15_6_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_246_bits = core_io_value_out_15_6_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_247_valid = core_io_value_out_15_7_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_247_bits = core_io_value_out_15_7_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_248_valid = core_io_value_out_15_8_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_248_bits = core_io_value_out_15_8_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_249_valid = core_io_value_out_15_9_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_249_bits = core_io_value_out_15_9_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_250_valid = core_io_value_out_15_10_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_250_bits = core_io_value_out_15_10_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_251_valid = core_io_value_out_15_11_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_251_bits = core_io_value_out_15_11_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_252_valid = core_io_value_out_15_12_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_252_bits = core_io_value_out_15_12_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_253_valid = core_io_value_out_15_13_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_253_bits = core_io_value_out_15_13_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_254_valid = core_io_value_out_15_14_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_254_bits = core_io_value_out_15_14_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_255_valid = core_io_value_out_15_15_valid; // @[Stab.scala 324:84]
  assign rmerge_io_stream_in_255_bits = core_io_value_out_15_15_bits; // @[Stab.scala 324:84]
  assign rmerge_io_stream_out_ready = io_value_out_ready; // @[Stab.scala 326:16]
endmodule
