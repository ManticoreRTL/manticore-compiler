module InstructionDecoder(
  input         clock,
  input         reset,
  output        io_instruction_ready,
  input         io_instruction_valid,
  input  [31:0] io_instruction_bits,
  input         io_decode_ready,
  output        io_decode_valid,
  output [4:0]  io_decode_bits_dest_reg,
  output [3:0]  io_decode_bits_exec_state,
  output        io_decode_bits_rt_as_op1,
  output        io_decode_bits_imm_u_as_op2,
  output        io_decode_bits_imm_s_as_op2,
  output        io_decode_bits_shamt_as_op2,
  output        io_decode_bits_rs_as_op2,
  output [3:0]  io_decode_bits_alu_funct
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[FemtoMips32.scala 131:23]
  reg [5:0] opcode; // @[FemtoMips32.scala 132:19]
  reg [5:0] funct; // @[FemtoMips32.scala 133:19]
  reg [4:0] rd; // @[FemtoMips32.scala 134:19]
  reg [4:0] rt; // @[FemtoMips32.scala 135:19]
  reg  alu_use_funct; // @[FemtoMips32.scala 138:26]
  reg [4:0] decode_result_dest_reg; // @[FemtoMips32.scala 139:26]
  reg [3:0] decode_result_exec_state; // @[FemtoMips32.scala 139:26]
  reg  decode_result_rt_as_op1; // @[FemtoMips32.scala 139:26]
  reg  decode_result_imm_u_as_op2; // @[FemtoMips32.scala 139:26]
  reg  decode_result_imm_s_as_op2; // @[FemtoMips32.scala 139:26]
  reg  decode_result_shamt_as_op2; // @[FemtoMips32.scala 139:26]
  reg  decode_result_rs_as_op2; // @[FemtoMips32.scala 139:26]
  wire  _T_3 = io_instruction_ready & io_instruction_valid; // @[Decoupled.scala 50:35]
  wire  _T_10 = io_decode_ready & io_decode_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _GEN_5 = _T_10 ? 2'h0 : state; // @[FemtoMips32.scala 161:28 162:15 131:23]
  wire  _GEN_9 = 2'h1 == state ? 1'h0 : 2'h2 == state; // @[FemtoMips32.scala 143:17 141:24]
  wire  _T_12 = funct < 6'h4; // @[FemtoMips32.scala 181:16]
  wire  _T_13 = funct < 6'h8; // @[FemtoMips32.scala 185:22]
  wire  _GEN_19 = funct < 6'h4 | _T_13; // @[FemtoMips32.scala 181:23 182:34]
  wire  _GEN_22 = funct < 6'h4 ? 1'h0 : _T_13; // @[FemtoMips32.scala 181:23 170:30]
  wire  _T_15 = opcode == 6'h4; // @[FemtoMips32.scala 194:21]
  wire  _decode_result_imm_u_as_op2_T_2 = funct == 6'h9 | funct == 6'hb; // @[FemtoMips32.scala 198:52]
  wire  _T_19 = opcode == 6'hf; // @[FemtoMips32.scala 201:21]
  wire  _T_21 = opcode == 6'h2b; // @[FemtoMips32.scala 209:21]
  wire [3:0] _GEN_23 = opcode == 6'h2b ? 4'h9 : 4'h4; // @[FemtoMips32.scala 174:28 209:29 210:32]
  wire [3:0] _GEN_25 = opcode == 6'h23 ? 4'h8 : _GEN_23; // @[FemtoMips32.scala 205:29 206:32]
  wire  _GEN_26 = opcode == 6'h23 | _T_21; // @[FemtoMips32.scala 205:29 207:32]
  wire [4:0] _GEN_27 = opcode == 6'h23 ? rt : 5'h0; // @[FemtoMips32.scala 175:28 205:29 208:32]
  wire [3:0] _GEN_28 = opcode == 6'hf ? 4'h4 : _GEN_25; // @[FemtoMips32.scala 201:30 202:32]
  wire [4:0] _GEN_29 = opcode == 6'hf ? rt : _GEN_27; // @[FemtoMips32.scala 201:30 203:32]
  wire  _GEN_30 = opcode == 6'hf | _GEN_26; // @[FemtoMips32.scala 201:30 204:32]
  wire  _GEN_32 = opcode < 6'hf & opcode > 6'h7 & (funct == 6'h9 | funct == 6'hb); // @[FemtoMips32.scala 169:30 196:45 198:32]
  wire  _alu_funct_T = funct == 6'h0; // @[FemtoMips32.scala 214:30]
  wire  _alu_funct_T_1 = funct == 6'h2; // @[FemtoMips32.scala 214:30]
  wire  _alu_funct_T_2 = funct == 6'h6; // @[FemtoMips32.scala 214:30]
  wire  _alu_funct_T_3 = _alu_funct_T_1 | _alu_funct_T_2; // @[FemtoMips32.scala 220:18]
  wire  _alu_funct_T_4 = funct == 6'h3; // @[FemtoMips32.scala 214:30]
  wire  _alu_funct_T_5 = funct == 6'h7; // @[FemtoMips32.scala 214:30]
  wire  _alu_funct_T_6 = _alu_funct_T_4 | _alu_funct_T_5; // @[FemtoMips32.scala 221:18]
  wire  _alu_funct_T_7 = funct == 6'h20; // @[FemtoMips32.scala 214:30]
  wire  _alu_funct_T_8 = funct == 6'h21; // @[FemtoMips32.scala 214:30]
  wire  _alu_funct_T_9 = funct == 6'h22; // @[FemtoMips32.scala 214:30]
  wire  _alu_funct_T_10 = funct == 6'h23; // @[FemtoMips32.scala 214:30]
  wire  _alu_funct_T_11 = funct == 6'h24; // @[FemtoMips32.scala 214:30]
  wire  _alu_funct_T_12 = funct == 6'h25; // @[FemtoMips32.scala 214:30]
  wire  _alu_funct_T_13 = funct == 6'h26; // @[FemtoMips32.scala 214:30]
  wire  _alu_funct_T_14 = funct == 6'h27; // @[FemtoMips32.scala 214:30]
  wire  _alu_funct_T_15 = funct == 6'h2a; // @[FemtoMips32.scala 214:30]
  wire  _alu_funct_T_16 = funct == 6'h2b; // @[FemtoMips32.scala 214:30]
  wire [3:0] _alu_funct_T_17 = _alu_funct_T_16 ? 4'ha : 4'h0; // @[Mux.scala 101:16]
  wire [3:0] _alu_funct_T_18 = _alu_funct_T_15 ? 4'h9 : _alu_funct_T_17; // @[Mux.scala 101:16]
  wire [3:0] _alu_funct_T_19 = _alu_funct_T_14 ? 4'h8 : _alu_funct_T_18; // @[Mux.scala 101:16]
  wire [3:0] _alu_funct_T_20 = _alu_funct_T_13 ? 4'h7 : _alu_funct_T_19; // @[Mux.scala 101:16]
  wire [3:0] _alu_funct_T_21 = _alu_funct_T_12 ? 4'h6 : _alu_funct_T_20; // @[Mux.scala 101:16]
  wire [4:0] _alu_funct_T_22 = _alu_funct_T_11 ? 5'h5 : {{1'd0}, _alu_funct_T_21}; // @[Mux.scala 101:16]
  wire [4:0] _alu_funct_T_23 = _alu_funct_T_10 ? 5'h4 : _alu_funct_T_22; // @[Mux.scala 101:16]
  wire [4:0] _alu_funct_T_24 = _alu_funct_T_9 ? 5'h4 : _alu_funct_T_23; // @[Mux.scala 101:16]
  wire [4:0] _alu_funct_T_25 = _alu_funct_T_8 ? 5'h3 : _alu_funct_T_24; // @[Mux.scala 101:16]
  wire [4:0] _alu_funct_T_26 = _alu_funct_T_7 ? 5'h3 : _alu_funct_T_25; // @[Mux.scala 101:16]
  wire [4:0] _alu_funct_T_27 = _alu_funct_T_6 ? 5'h2 : _alu_funct_T_26; // @[Mux.scala 101:16]
  wire [4:0] _alu_funct_T_28 = _alu_funct_T_3 ? 5'h1 : _alu_funct_T_27; // @[Mux.scala 101:16]
  wire [4:0] alu_funct = _alu_funct_T ? 5'h0 : _alu_funct_T_28; // @[Mux.scala 101:16]
  wire  _alu_opcode_T_1 = opcode == 6'h8; // @[FemtoMips32.scala 215:31]
  wire  _alu_opcode_T_2 = opcode == 6'h9; // @[FemtoMips32.scala 215:31]
  wire  _alu_opcode_T_3 = _alu_opcode_T_1 | _alu_opcode_T_2; // @[FemtoMips32.scala 238:19]
  wire  _alu_opcode_T_4 = opcode == 6'ha; // @[FemtoMips32.scala 215:31]
  wire  _alu_opcode_T_5 = opcode == 6'hb; // @[FemtoMips32.scala 215:31]
  wire  _alu_opcode_T_6 = opcode == 6'hc; // @[FemtoMips32.scala 215:31]
  wire  _alu_opcode_T_7 = opcode == 6'hd; // @[FemtoMips32.scala 215:31]
  wire  _alu_opcode_T_8 = opcode == 6'he; // @[FemtoMips32.scala 215:31]
  wire [3:0] _alu_opcode_T_13 = _GEN_26 ? 4'h3 : 4'h0; // @[Mux.scala 101:16]
  wire [3:0] _alu_opcode_T_14 = _T_19 ? 4'hb : _alu_opcode_T_13; // @[Mux.scala 101:16]
  wire [3:0] _alu_opcode_T_15 = _alu_opcode_T_8 ? 4'h7 : _alu_opcode_T_14; // @[Mux.scala 101:16]
  wire [3:0] _alu_opcode_T_16 = _alu_opcode_T_7 ? 4'h6 : _alu_opcode_T_15; // @[Mux.scala 101:16]
  wire [4:0] _alu_opcode_T_17 = _alu_opcode_T_6 ? 5'h5 : {{1'd0}, _alu_opcode_T_16}; // @[Mux.scala 101:16]
  wire [4:0] _alu_opcode_T_18 = _alu_opcode_T_5 ? 5'ha : _alu_opcode_T_17; // @[Mux.scala 101:16]
  wire [4:0] _alu_opcode_T_19 = _alu_opcode_T_4 ? 5'h9 : _alu_opcode_T_18; // @[Mux.scala 101:16]
  wire [4:0] _alu_opcode_T_20 = _alu_opcode_T_3 ? 5'h3 : _alu_opcode_T_19; // @[Mux.scala 101:16]
  wire [4:0] alu_opcode = _T_15 ? 5'h4 : _alu_opcode_T_20; // @[Mux.scala 101:16]
  wire [4:0] _io_decode_bits_alu_funct_T = alu_use_funct ? alu_funct : alu_opcode; // @[FemtoMips32.scala 249:34]
  assign io_instruction_ready = 2'h0 == state; // @[FemtoMips32.scala 143:17]
  assign io_decode_valid = 2'h0 == state ? 1'h0 : _GEN_9; // @[FemtoMips32.scala 143:17 141:24]
  assign io_decode_bits_dest_reg = decode_result_dest_reg; // @[FemtoMips32.scala 248:28]
  assign io_decode_bits_exec_state = decode_result_exec_state; // @[FemtoMips32.scala 248:28]
  assign io_decode_bits_rt_as_op1 = decode_result_rt_as_op1; // @[FemtoMips32.scala 248:28]
  assign io_decode_bits_imm_u_as_op2 = decode_result_imm_u_as_op2; // @[FemtoMips32.scala 248:28]
  assign io_decode_bits_imm_s_as_op2 = decode_result_imm_s_as_op2; // @[FemtoMips32.scala 248:28]
  assign io_decode_bits_shamt_as_op2 = decode_result_shamt_as_op2; // @[FemtoMips32.scala 248:28]
  assign io_decode_bits_rs_as_op2 = decode_result_rs_as_op2; // @[FemtoMips32.scala 248:28]
  assign io_decode_bits_alu_funct = _io_decode_bits_alu_funct_T[3:0]; // @[FemtoMips32.scala 249:28]
  always @(posedge clock) begin
    if (reset) begin // @[FemtoMips32.scala 131:23]
      state <= 2'h0; // @[FemtoMips32.scala 131:23]
    end else if (2'h0 == state) begin // @[FemtoMips32.scala 143:17]
      state <= {{1'd0}, _T_3};
    end else if (2'h1 == state) begin // @[FemtoMips32.scala 143:17]
      state <= 2'h2; // @[FemtoMips32.scala 157:13]
    end else if (2'h2 == state) begin // @[FemtoMips32.scala 143:17]
      state <= _GEN_5;
    end
    if (2'h0 == state) begin // @[FemtoMips32.scala 143:17]
      if (_T_3) begin // @[FemtoMips32.scala 146:33]
        opcode <= io_instruction_bits[31:26]; // @[FemtoMips32.scala 147:16]
      end
    end
    if (2'h0 == state) begin // @[FemtoMips32.scala 143:17]
      if (_T_3) begin // @[FemtoMips32.scala 146:33]
        funct <= io_instruction_bits[5:0]; // @[FemtoMips32.scala 148:16]
      end
    end
    if (2'h0 == state) begin // @[FemtoMips32.scala 143:17]
      if (_T_3) begin // @[FemtoMips32.scala 146:33]
        rd <= io_instruction_bits[15:11]; // @[FemtoMips32.scala 150:16]
      end
    end
    if (2'h0 == state) begin // @[FemtoMips32.scala 143:17]
      if (_T_3) begin // @[FemtoMips32.scala 146:33]
        rt <= io_instruction_bits[20:16]; // @[FemtoMips32.scala 149:16]
      end
    end
    alu_use_funct <= opcode == 6'h0; // @[FemtoMips32.scala 178:15]
    if (opcode == 6'h0) begin // @[FemtoMips32.scala 178:27]
      decode_result_dest_reg <= rd; // @[FemtoMips32.scala 179:30]
    end else if (opcode == 6'h2) begin // @[FemtoMips32.scala 192:31]
      decode_result_dest_reg <= 5'h0; // @[FemtoMips32.scala 175:28]
    end else if (opcode == 6'h4) begin // @[FemtoMips32.scala 194:30]
      decode_result_dest_reg <= 5'h0; // @[FemtoMips32.scala 175:28]
    end else if (opcode < 6'hf & opcode > 6'h7) begin // @[FemtoMips32.scala 196:45]
      decode_result_dest_reg <= rt; // @[FemtoMips32.scala 200:32]
    end else begin
      decode_result_dest_reg <= _GEN_29;
    end
    if (opcode == 6'h0) begin // @[FemtoMips32.scala 178:27]
      if (funct == 6'hd) begin // @[FemtoMips32.scala 180:36]
        decode_result_exec_state <= 4'hb;
      end else begin
        decode_result_exec_state <= 4'h4;
      end
    end else if (opcode == 6'h2) begin // @[FemtoMips32.scala 192:31]
      decode_result_exec_state <= 4'h6; // @[FemtoMips32.scala 193:30]
    end else if (opcode == 6'h4) begin // @[FemtoMips32.scala 194:30]
      decode_result_exec_state <= 4'h7; // @[FemtoMips32.scala 195:30]
    end else if (opcode < 6'hf & opcode > 6'h7) begin // @[FemtoMips32.scala 196:45]
      decode_result_exec_state <= 4'h4; // @[FemtoMips32.scala 197:32]
    end else begin
      decode_result_exec_state <= _GEN_28;
    end
    decode_result_rt_as_op1 <= opcode == 6'h0 & _GEN_19; // @[FemtoMips32.scala 178:27 172:30]
    if (opcode == 6'h0) begin // @[FemtoMips32.scala 178:27]
      decode_result_imm_u_as_op2 <= 1'h0; // @[FemtoMips32.scala 169:30]
    end else if (opcode == 6'h2) begin // @[FemtoMips32.scala 192:31]
      decode_result_imm_u_as_op2 <= 1'h0; // @[FemtoMips32.scala 169:30]
    end else if (opcode == 6'h4) begin // @[FemtoMips32.scala 194:30]
      decode_result_imm_u_as_op2 <= 1'h0; // @[FemtoMips32.scala 169:30]
    end else begin
      decode_result_imm_u_as_op2 <= _GEN_32;
    end
    if (opcode == 6'h0) begin // @[FemtoMips32.scala 178:27]
      decode_result_imm_s_as_op2 <= 1'h0; // @[FemtoMips32.scala 168:30]
    end else if (opcode == 6'h2) begin // @[FemtoMips32.scala 192:31]
      decode_result_imm_s_as_op2 <= 1'h0; // @[FemtoMips32.scala 168:30]
    end else if (opcode == 6'h4) begin // @[FemtoMips32.scala 194:30]
      decode_result_imm_s_as_op2 <= 1'h0; // @[FemtoMips32.scala 168:30]
    end else if (opcode < 6'hf & opcode > 6'h7) begin // @[FemtoMips32.scala 196:45]
      decode_result_imm_s_as_op2 <= ~_decode_result_imm_u_as_op2_T_2; // @[FemtoMips32.scala 199:32]
    end else begin
      decode_result_imm_s_as_op2 <= _GEN_30;
    end
    decode_result_shamt_as_op2 <= opcode == 6'h0 & _T_12; // @[FemtoMips32.scala 178:27 171:30]
    decode_result_rs_as_op2 <= opcode == 6'h0 & _GEN_22; // @[FemtoMips32.scala 178:27 170:30]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  opcode = _RAND_1[5:0];
  _RAND_2 = {1{`RANDOM}};
  funct = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  rd = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  rt = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  alu_use_funct = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  decode_result_dest_reg = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  decode_result_exec_state = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  decode_result_rt_as_op1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  decode_result_imm_u_as_op2 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  decode_result_imm_s_as_op2 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  decode_result_shamt_as_op2 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  decode_result_rs_as_op2 = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Alu(
  input         clock,
  input  [3:0]  io_funct,
  input  [31:0] io_rs,
  input  [31:0] io_rt,
  output [31:0] io_result
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire [4:0] shamt = io_rt[4:0]; // @[FemtoMips32.scala 101:32]
  wire [62:0] _GEN_2 = {{31'd0}, io_rs}; // @[FemtoMips32.scala 105:26]
  wire [62:0] _result_T = _GEN_2 << shamt; // @[FemtoMips32.scala 105:26]
  wire  _result_T_13 = io_rs == 32'h0; // @[FemtoMips32.scala 113:19]
  wire  _result_T_16 = $signed(io_rs) < $signed(io_rt); // @[FemtoMips32.scala 114:33]
  wire  _result_T_17 = io_rs < io_rt; // @[FemtoMips32.scala 115:26]
  wire [47:0] _GEN_0 = {io_rt, 16'h0}; // @[FemtoMips32.scala 116:26]
  wire [62:0] _result_T_18 = {{15'd0}, _GEN_0}; // @[FemtoMips32.scala 116:26]
  wire  _result_T_19 = io_funct == 4'h0; // @[FemtoMips32.scala 117:38]
  reg [31:0] result_r; // @[FemtoMips32.scala 96:16]
  wire  _result_T_20 = io_funct == 4'h1; // @[FemtoMips32.scala 117:38]
  reg [31:0] result_r_1; // @[FemtoMips32.scala 96:16]
  wire  _result_T_21 = io_funct == 4'h2; // @[FemtoMips32.scala 117:38]
  reg [31:0] result_r_2; // @[FemtoMips32.scala 96:16]
  wire  _result_T_22 = io_funct == 4'h3; // @[FemtoMips32.scala 117:38]
  reg [31:0] result_r_3; // @[FemtoMips32.scala 96:16]
  wire  _result_T_23 = io_funct == 4'h4; // @[FemtoMips32.scala 117:38]
  wire [4:0] _GEN_1 = {{1'd0}, io_funct}; // @[FemtoMips32.scala 117:38]
  wire  _result_T_24 = _GEN_1 == 5'h5; // @[FemtoMips32.scala 117:38]
  reg [31:0] result_r_5; // @[FemtoMips32.scala 96:16]
  wire  _result_T_25 = io_funct == 4'h6; // @[FemtoMips32.scala 117:38]
  reg [31:0] result_r_6; // @[FemtoMips32.scala 96:16]
  wire  _result_T_26 = io_funct == 4'h7; // @[FemtoMips32.scala 117:38]
  wire  _result_T_27 = io_funct == 4'h8; // @[FemtoMips32.scala 117:38]
  reg [31:0] result_r_8; // @[FemtoMips32.scala 96:16]
  wire  _result_T_28 = io_funct == 4'h9; // @[FemtoMips32.scala 117:38]
  reg [31:0] result_r_9; // @[FemtoMips32.scala 96:16]
  wire  _result_T_29 = io_funct == 4'ha; // @[FemtoMips32.scala 117:38]
  reg [31:0] result_r_10; // @[FemtoMips32.scala 96:16]
  wire  _result_T_30 = io_funct == 4'hb; // @[FemtoMips32.scala 117:38]
  reg [31:0] result_r_11; // @[FemtoMips32.scala 96:16]
  wire [31:0] _result_T_31 = _result_T_30 ? result_r_11 : 32'h0; // @[Mux.scala 101:16]
  wire [31:0] _result_T_32 = _result_T_29 ? result_r_10 : _result_T_31; // @[Mux.scala 101:16]
  wire [31:0] _result_T_33 = _result_T_28 ? result_r_9 : _result_T_32; // @[Mux.scala 101:16]
  wire [31:0] _result_T_34 = _result_T_27 ? result_r_8 : _result_T_33; // @[Mux.scala 101:16]
  wire [31:0] _result_T_35 = _result_T_26 ? 32'h0 : _result_T_34; // @[Mux.scala 101:16]
  wire [31:0] _result_T_36 = _result_T_25 ? result_r_6 : _result_T_35; // @[Mux.scala 101:16]
  wire [31:0] _result_T_37 = _result_T_24 ? result_r_5 : _result_T_36; // @[Mux.scala 101:16]
  wire [31:0] _result_T_38 = _result_T_23 ? 32'h0 : _result_T_37; // @[Mux.scala 101:16]
  wire [31:0] _result_T_39 = _result_T_22 ? result_r_3 : _result_T_38; // @[Mux.scala 101:16]
  wire [31:0] _result_T_40 = _result_T_21 ? result_r_2 : _result_T_39; // @[Mux.scala 101:16]
  wire [31:0] _result_T_41 = _result_T_20 ? result_r_1 : _result_T_40; // @[Mux.scala 101:16]
  assign io_result = _result_T_19 ? result_r : _result_T_41; // @[Mux.scala 101:16]
  always @(posedge clock) begin
    result_r <= _result_T[31:0]; // @[FemtoMips32.scala 97:7]
    result_r_1 <= io_rs >> shamt; // @[FemtoMips32.scala 106:26]
    result_r_2 <= $signed(io_rs) >>> shamt; // @[FemtoMips32.scala 107:43]
    result_r_3 <= io_rs + io_rt; // @[FemtoMips32.scala 108:26]
    result_r_5 <= io_rs & io_rt; // @[FemtoMips32.scala 110:26]
    result_r_6 <= io_rs; // @[FemtoMips32.scala 111:26]
    result_r_8 <= {{31'd0}, _result_T_13}; // @[FemtoMips32.scala 97:7]
    result_r_9 <= {{31'd0}, _result_T_16}; // @[FemtoMips32.scala 97:7]
    result_r_10 <= {{31'd0}, _result_T_17}; // @[FemtoMips32.scala 97:7]
    result_r_11 <= _result_T_18[31:0]; // @[FemtoMips32.scala 97:7]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  result_r = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  result_r_1 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  result_r_2 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  result_r_3 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  result_r_5 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  result_r_6 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  result_r_8 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  result_r_9 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  result_r_10 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  result_r_11 = _RAND_9[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FemtoMips32(
  input         clock,
  input         reset,
  input         io_mem_read_req_ready,
  output        io_mem_read_req_valid,
  output [31:0] io_mem_read_req_bits,
  output        io_mem_read_resp_ready,
  input         io_mem_read_resp_valid,
  input  [31:0] io_mem_read_resp_bits,
  input         io_mem_write_req_ready,
  output        io_mem_write_req_valid,
  output [31:0] io_mem_write_req_bits_addr,
  output [31:0] io_mem_write_req_bits_data
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
`endif // RANDOMIZE_REG_INIT
  wire  decode_clock; // @[FemtoMips32.scala 264:29]
  wire  decode_reset; // @[FemtoMips32.scala 264:29]
  wire  decode_io_instruction_ready; // @[FemtoMips32.scala 264:29]
  wire  decode_io_instruction_valid; // @[FemtoMips32.scala 264:29]
  wire [31:0] decode_io_instruction_bits; // @[FemtoMips32.scala 264:29]
  wire  decode_io_decode_ready; // @[FemtoMips32.scala 264:29]
  wire  decode_io_decode_valid; // @[FemtoMips32.scala 264:29]
  wire [4:0] decode_io_decode_bits_dest_reg; // @[FemtoMips32.scala 264:29]
  wire [3:0] decode_io_decode_bits_exec_state; // @[FemtoMips32.scala 264:29]
  wire  decode_io_decode_bits_rt_as_op1; // @[FemtoMips32.scala 264:29]
  wire  decode_io_decode_bits_imm_u_as_op2; // @[FemtoMips32.scala 264:29]
  wire  decode_io_decode_bits_imm_s_as_op2; // @[FemtoMips32.scala 264:29]
  wire  decode_io_decode_bits_shamt_as_op2; // @[FemtoMips32.scala 264:29]
  wire  decode_io_decode_bits_rs_as_op2; // @[FemtoMips32.scala 264:29]
  wire [3:0] decode_io_decode_bits_alu_funct; // @[FemtoMips32.scala 264:29]
  reg [31:0] register_file [0:31]; // @[FemtoMips32.scala 265:26]
  wire  register_file_rs_value_MPORT_en; // @[FemtoMips32.scala 265:26]
  wire [4:0] register_file_rs_value_MPORT_addr; // @[FemtoMips32.scala 265:26]
  wire [31:0] register_file_rs_value_MPORT_data; // @[FemtoMips32.scala 265:26]
  wire  register_file_rt_value_MPORT_en; // @[FemtoMips32.scala 265:26]
  wire [4:0] register_file_rt_value_MPORT_addr; // @[FemtoMips32.scala 265:26]
  wire [31:0] register_file_rt_value_MPORT_data; // @[FemtoMips32.scala 265:26]
  wire [31:0] register_file_MPORT_data; // @[FemtoMips32.scala 265:26]
  wire [4:0] register_file_MPORT_addr; // @[FemtoMips32.scala 265:26]
  wire  register_file_MPORT_mask; // @[FemtoMips32.scala 265:26]
  wire  register_file_MPORT_en; // @[FemtoMips32.scala 265:26]
  wire  alu_clock; // @[FemtoMips32.scala 267:19]
  wire [3:0] alu_io_funct; // @[FemtoMips32.scala 267:19]
  wire [31:0] alu_io_rs; // @[FemtoMips32.scala 267:19]
  wire [31:0] alu_io_rt; // @[FemtoMips32.scala 267:19]
  wire [31:0] alu_io_result; // @[FemtoMips32.scala 267:19]
  reg [3:0] state; // @[FemtoMips32.scala 271:28]
  reg [31:0] pc; // @[FemtoMips32.scala 272:28]
  reg [31:0] instruction; // @[FemtoMips32.scala 273:24]
  wire  imm_sign = instruction[15]; // @[FemtoMips32.scala 276:29]
  wire [31:0] shamt = {27'h0,instruction[10:6]}; // @[Cat.scala 31:58]
  wire [15:0] _imm_sext_T_1 = imm_sign ? 16'hffff : 16'h0; // @[Bitwise.scala 74:12]
  wire [31:0] imm_sext = {_imm_sext_T_1,instruction[15:0]}; // @[Cat.scala 31:58]
  wire [31:0] imm_zext = {16'h0,instruction[15:0]}; // @[Cat.scala 31:58]
  reg [4:0] decode_result_dest_reg; // @[FemtoMips32.scala 281:26]
  reg  decode_result_rt_as_op1; // @[FemtoMips32.scala 281:26]
  reg  decode_result_imm_u_as_op2; // @[FemtoMips32.scala 281:26]
  reg  decode_result_imm_s_as_op2; // @[FemtoMips32.scala 281:26]
  reg  decode_result_shamt_as_op2; // @[FemtoMips32.scala 281:26]
  reg  decode_result_rs_as_op2; // @[FemtoMips32.scala 281:26]
  reg [3:0] decode_result_alu_funct; // @[FemtoMips32.scala 281:26]
  wire  _T_2 = 4'h0 == state; // @[FemtoMips32.scala 327:17]
  wire  _T_21 = 4'h5 == state; // @[FemtoMips32.scala 327:17]
  wire  _T_36 = io_mem_read_resp_ready & io_mem_read_resp_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_39 = 4'h9 == state ? 1'h0 : 4'ha == state & _T_36; // @[FemtoMips32.scala 327:17]
  wire  _GEN_51 = 4'h6 == state ? 1'h0 : _GEN_39; // @[FemtoMips32.scala 327:17]
  wire  _GEN_62 = 4'h7 == state ? 1'h0 : _GEN_51; // @[FemtoMips32.scala 327:17]
  wire  _GEN_68 = 4'h5 == state | _GEN_62; // @[FemtoMips32.scala 327:17 369:17]
  wire  _GEN_80 = 4'h4 == state ? 1'h0 : _GEN_68; // @[FemtoMips32.scala 327:17]
  wire  _GEN_92 = 4'h3 == state ? 1'h0 : _GEN_80; // @[FemtoMips32.scala 327:17]
  wire  _GEN_105 = 4'h2 == state ? 1'h0 : _GEN_92; // @[FemtoMips32.scala 327:17]
  wire  _GEN_120 = 4'h1 == state ? 1'h0 : _GEN_105; // @[FemtoMips32.scala 327:17]
  wire [31:0] rt_value = register_file_rt_value_MPORT_data;
  wire [31:0] rs_value = register_file_rs_value_MPORT_data;
  wire [31:0] _alu_io_rt_T = decode_result_imm_u_as_op2 ? imm_zext : rt_value; // @[FemtoMips32.scala 309:52]
  wire [31:0] _alu_io_rt_T_1 = decode_result_imm_s_as_op2 ? imm_sext : _alu_io_rt_T; // @[FemtoMips32.scala 309:10]
  wire [31:0] _alu_io_rt_T_2 = decode_result_shamt_as_op2 ? shamt : _alu_io_rt_T_1; // @[FemtoMips32.scala 306:8]
  wire  _T_3 = io_mem_read_req_ready & io_mem_read_req_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _GEN_7 = _T_36 ? 2'h2 : 2'h1; // @[FemtoMips32.scala 339:35 341:21 343:15]
  wire  _T_11 = decode_io_instruction_ready & decode_io_instruction_valid; // @[Decoupled.scala 50:35]
  wire [1:0] _GEN_8 = _T_11 ? 2'h3 : 2'h2; // @[FemtoMips32.scala 348:40 349:15 351:15]
  wire  _T_15 = decode_io_decode_ready & decode_io_decode_valid; // @[Decoupled.scala 50:35]
  wire [3:0] _GEN_9 = _T_15 ? decode_io_decode_bits_exec_state : 4'h3; // @[FemtoMips32.scala 357:35 358:15 360:15]
  wire [31:0] _pc_T_1 = pc + 32'h4; // @[FemtoMips32.scala 373:19]
  wire [33:0] _pc_T_4 = {imm_zext, 2'h0}; // @[FemtoMips32.scala 377:36]
  wire [33:0] _GEN_143 = {{2'd0}, _pc_T_1}; // @[FemtoMips32.scala 377:24]
  wire [33:0] _pc_T_6 = _GEN_143 + _pc_T_4; // @[FemtoMips32.scala 377:24]
  wire [33:0] _GEN_10 = rs_value == rt_value ? _pc_T_6 : {{2'd0}, _pc_T_1}; // @[FemtoMips32.scala 376:35 377:12 379:12]
  wire [31:0] _pc_T_11 = {_pc_T_1[31:28],instruction[25:0],2'h0}; // @[Cat.scala 31:58]
  wire [31:0] _io_mem_read_req_bits_T_1 = imm_sext + rs_value; // @[FemtoMips32.scala 389:42]
  wire [3:0] _GEN_11 = _T_3 ? 4'ha : 4'h9; // @[FemtoMips32.scala 391:34 392:15 394:15]
  wire [3:0] _GEN_14 = _T_36 ? 4'h0 : 4'ha; // @[FemtoMips32.scala 399:35 404:15 407:15]
  wire [31:0] _GEN_15 = _T_36 ? _pc_T_1 : pc; // @[FemtoMips32.scala 399:35 405:15 272:28]
  wire  _T_40 = io_mem_write_req_ready & io_mem_write_req_valid; // @[Decoupled.scala 50:35]
  wire [3:0] _GEN_16 = _T_40 ? 4'h0 : 4'h8; // @[FemtoMips32.scala 415:35 416:15 419:15]
  wire [31:0] _GEN_17 = _T_40 ? _pc_T_1 : pc; // @[FemtoMips32.scala 415:35 417:15 272:28]
  wire [3:0] _GEN_19 = 4'hb == state ? 4'hb : state; // @[FemtoMips32.scala 327:17 425:17 271:28]
  wire [3:0] _GEN_23 = 4'h8 == state ? _GEN_16 : _GEN_19; // @[FemtoMips32.scala 327:17]
  wire [31:0] _GEN_24 = 4'h8 == state ? _GEN_17 : pc; // @[FemtoMips32.scala 327:17 272:28]
  wire [3:0] _GEN_29 = 4'ha == state ? _GEN_14 : _GEN_23; // @[FemtoMips32.scala 327:17]
  wire [31:0] _GEN_30 = 4'ha == state ? _GEN_15 : _GEN_24; // @[FemtoMips32.scala 327:17]
  wire  _GEN_31 = 4'ha == state ? 1'h0 : 4'h8 == state; // @[FemtoMips32.scala 327:17 325:25]
  wire [3:0] _GEN_37 = 4'h9 == state ? _GEN_11 : _GEN_29; // @[FemtoMips32.scala 327:17]
  wire  _GEN_38 = 4'h9 == state ? 1'h0 : 4'ha == state; // @[FemtoMips32.scala 327:17 320:26]
  wire [31:0] _GEN_41 = 4'h9 == state ? pc : _GEN_30; // @[FemtoMips32.scala 327:17 272:28]
  wire  _GEN_42 = 4'h9 == state ? 1'h0 : _GEN_31; // @[FemtoMips32.scala 327:17 325:25]
  wire [31:0] _GEN_46 = 4'h6 == state ? _pc_T_11 : _GEN_41; // @[FemtoMips32.scala 327:17 385:13]
  wire [3:0] _GEN_47 = 4'h6 == state ? 4'h0 : _GEN_37; // @[FemtoMips32.scala 327:17 386:13]
  wire  _GEN_49 = 4'h6 == state ? 1'h0 : 4'h9 == state; // @[FemtoMips32.scala 327:17 319:26]
  wire  _GEN_50 = 4'h6 == state ? 1'h0 : _GEN_38; // @[FemtoMips32.scala 327:17 320:26]
  wire  _GEN_53 = 4'h6 == state ? 1'h0 : _GEN_42; // @[FemtoMips32.scala 327:17 325:25]
  wire [33:0] _GEN_57 = 4'h7 == state ? _GEN_10 : {{2'd0}, _GEN_46}; // @[FemtoMips32.scala 327:17]
  wire [3:0] _GEN_58 = 4'h7 == state ? 4'h0 : _GEN_47; // @[FemtoMips32.scala 327:17 381:13]
  wire  _GEN_60 = 4'h7 == state ? 1'h0 : _GEN_49; // @[FemtoMips32.scala 327:17 319:26]
  wire  _GEN_61 = 4'h7 == state ? 1'h0 : _GEN_50; // @[FemtoMips32.scala 327:17 320:26]
  wire  _GEN_64 = 4'h7 == state ? 1'h0 : _GEN_53; // @[FemtoMips32.scala 327:17 325:25]
  wire [3:0] _GEN_70 = 4'h5 == state ? 4'h0 : _GEN_58; // @[FemtoMips32.scala 327:17 372:13]
  wire [33:0] _GEN_71 = 4'h5 == state ? {{2'd0}, _pc_T_1} : _GEN_57; // @[FemtoMips32.scala 327:17 373:13]
  wire  _GEN_73 = 4'h5 == state ? 1'h0 : _GEN_60; // @[FemtoMips32.scala 327:17 319:26]
  wire  _GEN_74 = 4'h5 == state ? 1'h0 : _GEN_61; // @[FemtoMips32.scala 327:17 320:26]
  wire  _GEN_75 = 4'h5 == state ? 1'h0 : _GEN_64; // @[FemtoMips32.scala 327:17 325:25]
  wire [3:0] _GEN_79 = 4'h4 == state ? 4'h5 : _GEN_70; // @[FemtoMips32.scala 327:17 364:13]
  wire [33:0] _GEN_82 = 4'h4 == state ? {{2'd0}, pc} : _GEN_71; // @[FemtoMips32.scala 327:17 272:28]
  wire  _GEN_84 = 4'h4 == state ? 1'h0 : _GEN_73; // @[FemtoMips32.scala 327:17 319:26]
  wire  _GEN_85 = 4'h4 == state ? 1'h0 : _GEN_74; // @[FemtoMips32.scala 327:17 320:26]
  wire  _GEN_86 = 4'h4 == state ? 1'h0 : _GEN_75; // @[FemtoMips32.scala 327:17 325:25]
  wire [3:0] _GEN_91 = 4'h3 == state ? _GEN_9 : _GEN_79; // @[FemtoMips32.scala 327:17]
  wire [33:0] _GEN_94 = 4'h3 == state ? {{2'd0}, pc} : _GEN_82; // @[FemtoMips32.scala 327:17 272:28]
  wire  _GEN_96 = 4'h3 == state ? 1'h0 : _GEN_84; // @[FemtoMips32.scala 327:17 319:26]
  wire  _GEN_97 = 4'h3 == state ? 1'h0 : _GEN_85; // @[FemtoMips32.scala 327:17 320:26]
  wire  _GEN_98 = 4'h3 == state ? 1'h0 : _GEN_86; // @[FemtoMips32.scala 327:17 325:25]
  wire  _GEN_104 = 4'h2 == state ? 1'h0 : 4'h3 == state; // @[FemtoMips32.scala 327:17 316:31]
  wire [33:0] _GEN_107 = 4'h2 == state ? {{2'd0}, pc} : _GEN_94; // @[FemtoMips32.scala 327:17 272:28]
  wire  _GEN_109 = 4'h2 == state ? 1'h0 : _GEN_96; // @[FemtoMips32.scala 327:17 319:26]
  wire  _GEN_110 = 4'h2 == state ? 1'h0 : _GEN_97; // @[FemtoMips32.scala 327:17 320:26]
  wire  _GEN_111 = 4'h2 == state ? 1'h0 : _GEN_98; // @[FemtoMips32.scala 327:17 325:25]
  wire  _GEN_115 = 4'h1 == state | _GEN_110; // @[FemtoMips32.scala 327:17 338:30]
  wire  _GEN_118 = 4'h1 == state ? 1'h0 : 4'h2 == state; // @[FemtoMips32.scala 327:17 314:31]
  wire  _GEN_119 = 4'h1 == state ? 1'h0 : _GEN_104; // @[FemtoMips32.scala 327:17 316:31]
  wire [33:0] _GEN_122 = 4'h1 == state ? {{2'd0}, pc} : _GEN_107; // @[FemtoMips32.scala 327:17 272:28]
  wire  _GEN_124 = 4'h1 == state ? 1'h0 : _GEN_109; // @[FemtoMips32.scala 327:17 319:26]
  wire  _GEN_125 = 4'h1 == state ? 1'h0 : _GEN_111; // @[FemtoMips32.scala 327:17 325:25]
  wire [33:0] _GEN_138 = 4'h0 == state ? {{2'd0}, pc} : _GEN_122; // @[FemtoMips32.scala 327:17 272:28]
  wire [33:0] _GEN_144 = reset ? 34'h0 : _GEN_138; // @[FemtoMips32.scala 272:{28,28}]
  InstructionDecoder decode ( // @[FemtoMips32.scala 264:29]
    .clock(decode_clock),
    .reset(decode_reset),
    .io_instruction_ready(decode_io_instruction_ready),
    .io_instruction_valid(decode_io_instruction_valid),
    .io_instruction_bits(decode_io_instruction_bits),
    .io_decode_ready(decode_io_decode_ready),
    .io_decode_valid(decode_io_decode_valid),
    .io_decode_bits_dest_reg(decode_io_decode_bits_dest_reg),
    .io_decode_bits_exec_state(decode_io_decode_bits_exec_state),
    .io_decode_bits_rt_as_op1(decode_io_decode_bits_rt_as_op1),
    .io_decode_bits_imm_u_as_op2(decode_io_decode_bits_imm_u_as_op2),
    .io_decode_bits_imm_s_as_op2(decode_io_decode_bits_imm_s_as_op2),
    .io_decode_bits_shamt_as_op2(decode_io_decode_bits_shamt_as_op2),
    .io_decode_bits_rs_as_op2(decode_io_decode_bits_rs_as_op2),
    .io_decode_bits_alu_funct(decode_io_decode_bits_alu_funct)
  );
  Alu alu ( // @[FemtoMips32.scala 267:19]
    .clock(alu_clock),
    .io_funct(alu_io_funct),
    .io_rs(alu_io_rs),
    .io_rt(alu_io_rt),
    .io_result(alu_io_result)
  );
  assign register_file_rs_value_MPORT_en = 1'h1;
  assign register_file_rs_value_MPORT_addr = instruction[25:21];
  assign register_file_rs_value_MPORT_data = register_file[register_file_rs_value_MPORT_addr]; // @[FemtoMips32.scala 265:26]
  assign register_file_rt_value_MPORT_en = 1'h1;
  assign register_file_rt_value_MPORT_addr = instruction[20:16];
  assign register_file_rt_value_MPORT_data = register_file[register_file_rt_value_MPORT_addr]; // @[FemtoMips32.scala 265:26]
  assign register_file_MPORT_data = _T_21 ? alu_io_result : io_mem_read_resp_bits;
  assign register_file_MPORT_addr = decode_result_dest_reg;
  assign register_file_MPORT_mask = 1'h1;
  assign register_file_MPORT_en = _T_2 ? 1'h0 : _GEN_120;
  assign io_mem_read_req_valid = 4'h0 == state | _GEN_124; // @[FemtoMips32.scala 327:17 329:29]
  assign io_mem_read_req_bits = 4'h0 == state ? pc : _io_mem_read_req_bits_T_1; // @[FemtoMips32.scala 327:17 330:29]
  assign io_mem_read_resp_ready = 4'h0 == state ? 1'h0 : _GEN_115; // @[FemtoMips32.scala 327:17 320:26]
  assign io_mem_write_req_valid = 4'h0 == state ? 1'h0 : _GEN_125; // @[FemtoMips32.scala 327:17 325:25]
  assign io_mem_write_req_bits_addr = imm_sext + rs_value; // @[FemtoMips32.scala 414:47]
  assign io_mem_write_req_bits_data = register_file_rt_value_MPORT_data; // @[FemtoMips32.scala 327:17 413:34]
  assign decode_clock = clock;
  assign decode_reset = reset;
  assign decode_io_instruction_valid = 4'h0 == state ? 1'h0 : _GEN_118; // @[FemtoMips32.scala 327:17 314:31]
  assign decode_io_instruction_bits = instruction; // @[FemtoMips32.scala 315:31]
  assign decode_io_decode_ready = 4'h0 == state ? 1'h0 : _GEN_119; // @[FemtoMips32.scala 327:17 316:31]
  assign alu_clock = clock;
  assign alu_io_funct = decode_result_alu_funct; // @[FemtoMips32.scala 312:16]
  assign alu_io_rs = decode_result_rt_as_op1 ? rt_value : rs_value; // @[FemtoMips32.scala 297:19]
  assign alu_io_rt = decode_result_rs_as_op2 ? rs_value : _alu_io_rt_T_2; // @[FemtoMips32.scala 303:19]
  always @(posedge clock) begin
    if (register_file_MPORT_en & register_file_MPORT_mask) begin
      register_file[register_file_MPORT_addr] <= register_file_MPORT_data; // @[FemtoMips32.scala 265:26]
    end
    if (reset) begin // @[FemtoMips32.scala 271:28]
      state <= 4'h0; // @[FemtoMips32.scala 271:28]
    end else if (4'h0 == state) begin // @[FemtoMips32.scala 327:17]
      state <= {{3'd0}, _T_3};
    end else if (4'h1 == state) begin // @[FemtoMips32.scala 327:17]
      state <= {{2'd0}, _GEN_7};
    end else if (4'h2 == state) begin // @[FemtoMips32.scala 327:17]
      state <= {{2'd0}, _GEN_8};
    end else begin
      state <= _GEN_91;
    end
    pc <= _GEN_144[31:0]; // @[FemtoMips32.scala 272:{28,28}]
    if (!(4'h0 == state)) begin // @[FemtoMips32.scala 327:17]
      if (4'h1 == state) begin // @[FemtoMips32.scala 327:17]
        if (_T_36) begin // @[FemtoMips32.scala 339:35]
          instruction <= io_mem_read_resp_bits; // @[FemtoMips32.scala 340:21]
        end
      end
    end
    decode_result_dest_reg <= decode_io_decode_bits_dest_reg; // @[FemtoMips32.scala 317:31]
    decode_result_rt_as_op1 <= decode_io_decode_bits_rt_as_op1; // @[FemtoMips32.scala 317:31]
    decode_result_imm_u_as_op2 <= decode_io_decode_bits_imm_u_as_op2; // @[FemtoMips32.scala 317:31]
    decode_result_imm_s_as_op2 <= decode_io_decode_bits_imm_s_as_op2; // @[FemtoMips32.scala 317:31]
    decode_result_shamt_as_op2 <= decode_io_decode_bits_shamt_as_op2; // @[FemtoMips32.scala 317:31]
    decode_result_rs_as_op2 <= decode_io_decode_bits_rs_as_op2; // @[FemtoMips32.scala 317:31]
    decode_result_alu_funct <= decode_io_decode_bits_alu_funct; // @[FemtoMips32.scala 317:31]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    register_file[initvar] = _RAND_0[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  pc = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  instruction = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  decode_result_dest_reg = _RAND_4[4:0];
  _RAND_5 = {1{`RANDOM}};
  decode_result_rt_as_op1 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  decode_result_imm_u_as_op2 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  decode_result_imm_s_as_op2 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  decode_result_shamt_as_op2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  decode_result_rs_as_op2 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  decode_result_alu_funct = _RAND_10[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RouterBuffer(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [31:0] io_enq_bits_address,
  input  [31:0] io_enq_bits_data,
  input         io_enq_bits_wen,
  input  [7:0]  io_enq_bits_id,
  input         io_deq_ready,
  output        io_deq_valid,
  output [31:0] io_deq_bits_address,
  output [31:0] io_deq_bits_data,
  output        io_deq_bits_wen,
  output [7:0]  io_deq_bits_id
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] storage_address; // @[FemtroRing.scala 34:20]
  reg [31:0] storage_data; // @[FemtroRing.scala 34:20]
  reg  storage_wen; // @[FemtroRing.scala 34:20]
  reg [7:0] storage_id; // @[FemtroRing.scala 34:20]
  reg  full; // @[FemtroRing.scala 35:24]
  wire  _T = io_enq_ready & io_enq_valid; // @[Decoupled.scala 50:35]
  wire  _GEN_0 = _T | full; // @[FemtroRing.scala 41:21 42:13 35:24]
  wire  _T_1 = io_deq_ready & io_deq_valid; // @[Decoupled.scala 50:35]
  assign io_enq_ready = ~full; // @[FemtroRing.scala 37:19]
  assign io_deq_valid = full; // @[FemtroRing.scala 38:16]
  assign io_deq_bits_address = storage_address; // @[FemtroRing.scala 39:16]
  assign io_deq_bits_data = storage_data; // @[FemtroRing.scala 39:16]
  assign io_deq_bits_wen = storage_wen; // @[FemtroRing.scala 39:16]
  assign io_deq_bits_id = storage_id; // @[FemtroRing.scala 39:16]
  always @(posedge clock) begin
    if (_T) begin // @[FemtroRing.scala 41:21]
      storage_address <= io_enq_bits_address; // @[FemtroRing.scala 43:13]
    end
    if (_T) begin // @[FemtroRing.scala 41:21]
      storage_data <= io_enq_bits_data; // @[FemtroRing.scala 43:13]
    end
    if (_T) begin // @[FemtroRing.scala 41:21]
      storage_wen <= io_enq_bits_wen; // @[FemtroRing.scala 43:13]
    end
    if (_T) begin // @[FemtroRing.scala 41:21]
      storage_id <= io_enq_bits_id; // @[FemtroRing.scala 43:13]
    end
    if (reset) begin // @[FemtroRing.scala 35:24]
      full <= 1'h0; // @[FemtroRing.scala 35:24]
    end else if (_T_1) begin // @[FemtroRing.scala 46:21]
      full <= 1'h0; // @[FemtroRing.scala 47:10]
    end else begin
      full <= _GEN_0;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  storage_address = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  storage_data = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  storage_wen = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  storage_id = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  full = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Router(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h1 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h1 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h1 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h1; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_1(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h2 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h2 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h2 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_1(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_1 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h2; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_2(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h3 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h3 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h3 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_2(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_2 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h3; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_3(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h4 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h4 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h4 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_3(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_3 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h4; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_4(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h5 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h5 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h5 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_4(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_4 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h5; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_5(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h6 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h6 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h6 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_5(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_5 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h6; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_6(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h7 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h7 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h7 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_6(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_6 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h7; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_7(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h8 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h8 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h8 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_7(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_7 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h8; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_8(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h9 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h9 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h9 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_8(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_8 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h9; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_9(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'ha ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'ha & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'ha ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_9(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_9 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'ha; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_10(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'hb ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'hb & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'hb ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_10(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_10 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'hb; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_11(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'hc ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'hc & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'hc ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_11(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_11 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'hc; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_12(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'hd ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'hd & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'hd ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_12(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_12 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'hd; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_13(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'he ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'he & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'he ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_13(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_13 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'he; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_14(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'hf ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'hf & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'hf ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_14(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_14 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'hf; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_15(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h10 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h10 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h10 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_15(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_15 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h10; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_16(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h11 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h11 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h11 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_16(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_16 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h11; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_17(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h12 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h12 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h12 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_17(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_17 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h12; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_18(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h13 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h13 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h13 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_18(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_18 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h13; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_19(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h14 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h14 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h14 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_19(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_19 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h14; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_20(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h15 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h15 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h15 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_20(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_20 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h15; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_21(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h16 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h16 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h16 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_21(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_21 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h16; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_22(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h17 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h17 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h17 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_22(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_22 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h17; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_23(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h18 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h18 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h18 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_23(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_23 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h18; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_24(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h19 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h19 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h19 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_24(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_24 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h19; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_25(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h1a ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h1a & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h1a ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_25(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_25 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h1a; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_26(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h1b ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h1b & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h1b ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_26(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_26 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h1b; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_27(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h1c ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h1c & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h1c ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_27(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_27 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h1c; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_28(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h1d ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h1d & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h1d ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_28(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_28 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h1d; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_29(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h1e ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h1e & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h1e ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_29(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_29 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h1e; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_30(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h1f ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h1f & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h1f ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_30(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_30 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h1f; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_31(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h20 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h20 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h20 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_31(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_31 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h20; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_32(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h21 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h21 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h21 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_32(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_32 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h21; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_33(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h22 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h22 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h22 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_33(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_33 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h22; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_34(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h23 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h23 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h23 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_34(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_34 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h23; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_35(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h24 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h24 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h24 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_35(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_35 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h24; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_36(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h25 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h25 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h25 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_36(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_36 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h25; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_37(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h26 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h26 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h26 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_37(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_37 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h26; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_38(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h27 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h27 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h27 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_38(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_38 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h27; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_39(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h28 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h28 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h28 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_39(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_39 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h28; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_40(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h29 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h29 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h29 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_40(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_40 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h29; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_41(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h2a ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h2a & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h2a ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_41(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_41 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h2a; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_42(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h2b ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h2b & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h2b ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_42(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_42 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h2b; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_43(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h2c ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h2c & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h2c ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_43(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_43 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h2c; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_44(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h2d ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h2d & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h2d ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_44(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_44 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h2d; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_45(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h2e ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h2e & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h2e ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_45(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_45 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h2e; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_46(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h2f ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h2f & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h2f ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_46(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_46 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h2f; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_47(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h30 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h30 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h30 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_47(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_47 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h30; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_48(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h31 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h31 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h31 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_48(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_48 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h31; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_49(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h32 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h32 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h32 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_49(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_49 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h32; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_50(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h33 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h33 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h33 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_50(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_50 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h33; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_51(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h34 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h34 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h34 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_51(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_51 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h34; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_52(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h35 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h35 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h35 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_52(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_52 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h35; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_53(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h36 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h36 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h36 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_53(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_53 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h36; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_54(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h37 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h37 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h37 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_54(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_54 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h37; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_55(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h38 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h38 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h38 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_55(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_55 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h38; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_56(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h39 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h39 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h39 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_56(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_56 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h39; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_57(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h3a ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h3a & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h3a ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_57(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_57 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h3a; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_58(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h3b ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h3b & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h3b ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_58(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_58 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h3b; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_59(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h3c ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h3c & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h3c ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_59(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_59 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h3c; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_60(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h3d ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h3d & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h3d ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_60(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_60 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h3d; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_61(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h3e ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h3e & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h3e ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_61(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_61 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h3e; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_62(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h3f ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h3f & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h3f ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_62(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_62 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h3f; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_63(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h40 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h40 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h40 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_63(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_63 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h40; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_64(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h41 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h41 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h41 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_64(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_64 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h41; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_65(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h42 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h42 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h42 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_65(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_65 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h42; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_66(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h43 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h43 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h43 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_66(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_66 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h43; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_67(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h44 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h44 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h44 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_67(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_67 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h44; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_68(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h45 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h45 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h45 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_68(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_68 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h45; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_69(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h46 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h46 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h46 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_69(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_69 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h46; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_70(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h47 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h47 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h47 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_70(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_70 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h47; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_71(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h48 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h48 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h48 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_71(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_71 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h48; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_72(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h49 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h49 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h49 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_72(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_72 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h49; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_73(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h4a ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h4a & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h4a ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_73(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_73 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h4a; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_74(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h4b ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h4b & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h4b ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_74(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_74 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h4b; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_75(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h4c ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h4c & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h4c ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_75(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_75 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h4c; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_76(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h4d ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h4d & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h4d ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_76(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_76 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h4d; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_77(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h4e ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h4e & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h4e ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_77(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_77 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h4e; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_78(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h4f ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h4f & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h4f ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_78(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_78 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h4f; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_79(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h50 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h50 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h50 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_79(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_79 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h50; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_80(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h51 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h51 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h51 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_80(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_80 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h51; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_81(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h52 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h52 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h52 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_81(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_81 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h52; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_82(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h53 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h53 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h53 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_82(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_82 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h53; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_83(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h54 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h54 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h54 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_83(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_83 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h54; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_84(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h55 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h55 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h55 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_84(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_84 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h55; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_85(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h56 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h56 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h56 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_85(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_85 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h56; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_86(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h57 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h57 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h57 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_86(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_86 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h57; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_87(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h58 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h58 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h58 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_87(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_87 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h58; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_88(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h59 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h59 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h59 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_88(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_88 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h59; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_89(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h5a ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h5a & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h5a ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_89(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_89 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h5a; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_90(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h5b ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h5b & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h5b ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_90(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_90 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h5b; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_91(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h5c ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h5c & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h5c ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_91(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_91 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h5c; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_92(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h5d ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h5d & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h5d ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_92(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_92 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h5d; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_93(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h5e ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h5e & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h5e ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_93(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_93 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h5e; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_94(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h5f ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h5f & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h5f ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_94(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_94 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h5f; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_95(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h60 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h60 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h60 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_95(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_95 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h60; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_96(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h61 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h61 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h61 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_96(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_96 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h61; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_97(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h62 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h62 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h62 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_97(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_97 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h62; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_98(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h63 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h63 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h63 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_98(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_98 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h63; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_99(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h64 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h64 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h64 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_99(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_99 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h64; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_100(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h65 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h65 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h65 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_100(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_100 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h65; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_101(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h66 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h66 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h66 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_101(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_101 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h66; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_102(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h67 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h67 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h67 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_102(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_102 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h67; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_103(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h68 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h68 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h68 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_103(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_103 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h68; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_104(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h69 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h69 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h69 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_104(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_104 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h69; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_105(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h6a ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h6a & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h6a ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_105(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_105 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h6a; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_106(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h6b ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h6b & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h6b ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_106(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_106 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h6b; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_107(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h6c ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h6c & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h6c ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_107(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_107 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h6c; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_108(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h6d ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h6d & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h6d ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_108(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_108 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h6d; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_109(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h6e ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h6e & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h6e ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_109(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_109 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h6e; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_110(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h6f ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h6f & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h6f ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_110(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_110 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h6f; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_111(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h70 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h70 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h70 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_111(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_111 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h70; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_112(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h71 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h71 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h71 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_112(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_112 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h71; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_113(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h72 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h72 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h72 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_113(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_113 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h72; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_114(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h73 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h73 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h73 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_114(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_114 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h73; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_115(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h74 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h74 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h74 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_115(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_115 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h74; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_116(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h75 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h75 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h75 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_116(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_116 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h75; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_117(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h76 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h76 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h76 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_117(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_117 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h76; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_118(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h77 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h77 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h77 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_118(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_118 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h77; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_119(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h78 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h78 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h78 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_119(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_119 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h78; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_120(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h79 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h79 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h79 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_120(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_120 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h79; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_121(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h7a ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h7a & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h7a ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_121(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_121 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h7a; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_122(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h7b ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h7b & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h7b ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_122(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_122 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h7b; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_123(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h7c ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h7c & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h7c ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_123(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_123 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h7c; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_124(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h7d ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h7d & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h7d ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_124(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_124 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h7d; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_125(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h7e ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h7e & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h7e ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_125(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_125 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h7e; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_126(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h7f ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h7f & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h7f ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_126(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_126 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h7f; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module Router_127(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_coreReq_ready,
  input         io_coreReq_valid,
  input  [31:0] io_coreReq_bits_address,
  input  [31:0] io_coreReq_bits_data,
  input         io_coreReq_bits_wen,
  input         io_coreResp_ready,
  output        io_coreResp_valid,
  output [31:0] io_coreResp_bits_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  packet_clock; // @[FemtroRing.scala 54:26]
  wire  packet_reset; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_enq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_enq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_enq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_ready; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_valid; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_address; // @[FemtroRing.scala 54:26]
  wire [31:0] packet_io_deq_bits_data; // @[FemtroRing.scala 54:26]
  wire  packet_io_deq_bits_wen; // @[FemtroRing.scala 54:26]
  wire [7:0] packet_io_deq_bits_id; // @[FemtroRing.scala 54:26]
  wire  packetCore_clock; // @[FemtroRing.scala 55:26]
  wire  packetCore_reset; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_enq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_enq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_enq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_ready; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_valid; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_address; // @[FemtroRing.scala 55:26]
  wire [31:0] packetCore_io_deq_bits_data; // @[FemtroRing.scala 55:26]
  wire  packetCore_io_deq_bits_wen; // @[FemtroRing.scala 55:26]
  wire [7:0] packetCore_io_deq_bits_id; // @[FemtroRing.scala 55:26]
  wire  packetNext_clock; // @[FemtroRing.scala 56:26]
  wire  packetNext_reset; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_enq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_enq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_enq_bits_id; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_ready; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_valid; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_address; // @[FemtroRing.scala 56:26]
  wire [31:0] packetNext_io_deq_bits_data; // @[FemtroRing.scala 56:26]
  wire  packetNext_io_deq_bits_wen; // @[FemtroRing.scala 56:26]
  wire [7:0] packetNext_io_deq_bits_id; // @[FemtroRing.scala 56:26]
  reg  input_turn; // @[FemtroRing.scala 77:27]
  RouterBuffer packet ( // @[FemtroRing.scala 54:26]
    .clock(packet_clock),
    .reset(packet_reset),
    .io_enq_ready(packet_io_enq_ready),
    .io_enq_valid(packet_io_enq_valid),
    .io_enq_bits_address(packet_io_enq_bits_address),
    .io_enq_bits_data(packet_io_enq_bits_data),
    .io_enq_bits_wen(packet_io_enq_bits_wen),
    .io_enq_bits_id(packet_io_enq_bits_id),
    .io_deq_ready(packet_io_deq_ready),
    .io_deq_valid(packet_io_deq_valid),
    .io_deq_bits_address(packet_io_deq_bits_address),
    .io_deq_bits_data(packet_io_deq_bits_data),
    .io_deq_bits_wen(packet_io_deq_bits_wen),
    .io_deq_bits_id(packet_io_deq_bits_id)
  );
  RouterBuffer packetCore ( // @[FemtroRing.scala 55:26]
    .clock(packetCore_clock),
    .reset(packetCore_reset),
    .io_enq_ready(packetCore_io_enq_ready),
    .io_enq_valid(packetCore_io_enq_valid),
    .io_enq_bits_address(packetCore_io_enq_bits_address),
    .io_enq_bits_data(packetCore_io_enq_bits_data),
    .io_enq_bits_wen(packetCore_io_enq_bits_wen),
    .io_enq_bits_id(packetCore_io_enq_bits_id),
    .io_deq_ready(packetCore_io_deq_ready),
    .io_deq_valid(packetCore_io_deq_valid),
    .io_deq_bits_address(packetCore_io_deq_bits_address),
    .io_deq_bits_data(packetCore_io_deq_bits_data),
    .io_deq_bits_wen(packetCore_io_deq_bits_wen),
    .io_deq_bits_id(packetCore_io_deq_bits_id)
  );
  RouterBuffer packetNext ( // @[FemtroRing.scala 56:26]
    .clock(packetNext_clock),
    .reset(packetNext_reset),
    .io_enq_ready(packetNext_io_enq_ready),
    .io_enq_valid(packetNext_io_enq_valid),
    .io_enq_bits_address(packetNext_io_enq_bits_address),
    .io_enq_bits_data(packetNext_io_enq_bits_data),
    .io_enq_bits_wen(packetNext_io_enq_bits_wen),
    .io_enq_bits_id(packetNext_io_enq_bits_id),
    .io_deq_ready(packetNext_io_deq_ready),
    .io_deq_valid(packetNext_io_deq_valid),
    .io_deq_bits_address(packetNext_io_deq_bits_address),
    .io_deq_bits_data(packetNext_io_deq_bits_data),
    .io_deq_bits_wen(packetNext_io_deq_bits_wen),
    .io_deq_bits_id(packetNext_io_deq_bits_id)
  );
  assign io_prev_ready = input_turn & packet_io_enq_ready; // @[FemtroRing.scala 85:20 86:19 80:26]
  assign io_next_valid = packetNext_io_deq_valid; // @[FemtroRing.scala 58:11]
  assign io_next_bits_address = packetNext_io_deq_bits_address; // @[FemtroRing.scala 58:11]
  assign io_next_bits_data = packetNext_io_deq_bits_data; // @[FemtroRing.scala 58:11]
  assign io_next_bits_wen = packetNext_io_deq_bits_wen; // @[FemtroRing.scala 58:11]
  assign io_next_bits_id = packetNext_io_deq_bits_id; // @[FemtroRing.scala 58:11]
  assign io_coreReq_ready = input_turn ? 1'h0 : packet_io_enq_ready; // @[FemtroRing.scala 85:20 81:26 88:19]
  assign io_coreResp_valid = packetCore_io_deq_valid; // @[FemtroRing.scala 59:15]
  assign io_coreResp_bits_data = packetCore_io_deq_bits_data; // @[FemtroRing.scala 59:15]
  assign packet_clock = clock;
  assign packet_reset = reset;
  assign packet_io_enq_valid = input_turn ? io_prev_valid : io_coreReq_valid; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_address = input_turn ? io_prev_bits_address : io_coreReq_bits_address; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_data = input_turn ? io_prev_bits_data : io_coreReq_bits_data; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_wen = input_turn ? io_prev_bits_wen : io_coreReq_bits_wen; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_enq_bits_id = input_turn ? io_prev_bits_id : 8'h0; // @[FemtroRing.scala 85:20 86:19 88:19]
  assign packet_io_deq_ready = packet_io_deq_bits_id == 8'h80 ? packetCore_io_enq_ready : packetNext_io_enq_ready; // @[FemtroRing.scala 69:41 70:23 73:23]
  assign packetCore_clock = clock;
  assign packetCore_reset = reset;
  assign packetCore_io_enq_valid = packet_io_deq_bits_id == 8'h80 & packet_io_deq_valid; // @[FemtroRing.scala 69:41 70:23 65:27]
  assign packetCore_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetCore_io_deq_ready = io_coreResp_ready; // @[FemtroRing.scala 59:15]
  assign packetNext_clock = clock;
  assign packetNext_reset = reset;
  assign packetNext_io_enq_valid = packet_io_deq_bits_id == 8'h80 ? 1'h0 : packet_io_deq_valid; // @[FemtroRing.scala 63:27 69:41 73:23]
  assign packetNext_io_enq_bits_address = packet_io_deq_bits_address; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_data = packet_io_deq_bits_data; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_wen = packet_io_deq_bits_wen; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_enq_bits_id = packet_io_deq_bits_id; // @[FemtroRing.scala 69:41 70:23 66:27]
  assign packetNext_io_deq_ready = io_next_ready; // @[FemtroRing.scala 58:11]
  always @(posedge clock) begin
    if (reset) begin // @[FemtroRing.scala 77:27]
      input_turn <= 1'h0; // @[FemtroRing.scala 77:27]
    end else begin
      input_turn <= ~input_turn; // @[FemtroRing.scala 78:14]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  input_turn = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module RingCore_127(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id
);
  wire  core_clock; // @[FemtoMips32.scala 442:22]
  wire  core_reset; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_req_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_read_resp_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_read_resp_bits; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_ready; // @[FemtoMips32.scala 442:22]
  wire  core_io_mem_write_req_valid; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_addr; // @[FemtoMips32.scala 442:22]
  wire [31:0] core_io_mem_write_req_bits_data; // @[FemtoMips32.scala 442:22]
  wire  router_clock; // @[FemtoMips32.scala 443:22]
  wire  router_reset; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_prev_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_prev_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_prev_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_next_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_next_bits_wen; // @[FemtoMips32.scala 443:22]
  wire [7:0] router_io_next_bits_id; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_address; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreReq_bits_data; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreReq_bits_wen; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_ready; // @[FemtoMips32.scala 443:22]
  wire  router_io_coreResp_valid; // @[FemtoMips32.scala 443:22]
  wire [31:0] router_io_coreResp_bits_data; // @[FemtoMips32.scala 443:22]
  FemtoMips32 core ( // @[FemtoMips32.scala 442:22]
    .clock(core_clock),
    .reset(core_reset),
    .io_mem_read_req_ready(core_io_mem_read_req_ready),
    .io_mem_read_req_valid(core_io_mem_read_req_valid),
    .io_mem_read_req_bits(core_io_mem_read_req_bits),
    .io_mem_read_resp_ready(core_io_mem_read_resp_ready),
    .io_mem_read_resp_valid(core_io_mem_read_resp_valid),
    .io_mem_read_resp_bits(core_io_mem_read_resp_bits),
    .io_mem_write_req_ready(core_io_mem_write_req_ready),
    .io_mem_write_req_valid(core_io_mem_write_req_valid),
    .io_mem_write_req_bits_addr(core_io_mem_write_req_bits_addr),
    .io_mem_write_req_bits_data(core_io_mem_write_req_bits_data)
  );
  Router_127 router ( // @[FemtoMips32.scala 443:22]
    .clock(router_clock),
    .reset(router_reset),
    .io_prev_ready(router_io_prev_ready),
    .io_prev_valid(router_io_prev_valid),
    .io_prev_bits_address(router_io_prev_bits_address),
    .io_prev_bits_data(router_io_prev_bits_data),
    .io_prev_bits_wen(router_io_prev_bits_wen),
    .io_prev_bits_id(router_io_prev_bits_id),
    .io_next_ready(router_io_next_ready),
    .io_next_valid(router_io_next_valid),
    .io_next_bits_address(router_io_next_bits_address),
    .io_next_bits_data(router_io_next_bits_data),
    .io_next_bits_wen(router_io_next_bits_wen),
    .io_next_bits_id(router_io_next_bits_id),
    .io_coreReq_ready(router_io_coreReq_ready),
    .io_coreReq_valid(router_io_coreReq_valid),
    .io_coreReq_bits_address(router_io_coreReq_bits_address),
    .io_coreReq_bits_data(router_io_coreReq_bits_data),
    .io_coreReq_bits_wen(router_io_coreReq_bits_wen),
    .io_coreResp_ready(router_io_coreResp_ready),
    .io_coreResp_valid(router_io_coreResp_valid),
    .io_coreResp_bits_data(router_io_coreResp_bits_data)
  );
  assign io_prev_ready = router_io_prev_ready; // @[FemtoMips32.scala 463:11]
  assign io_next_valid = router_io_next_valid; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_address = router_io_next_bits_address; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_data = router_io_next_bits_data; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_wen = router_io_next_bits_wen; // @[FemtoMips32.scala 464:11]
  assign io_next_bits_id = router_io_next_bits_id; // @[FemtoMips32.scala 464:11]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_mem_read_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 446:30]
  assign core_io_mem_read_resp_valid = router_io_coreResp_valid; // @[FemtoMips32.scala 458:31]
  assign core_io_mem_read_resp_bits = router_io_coreResp_bits_data; // @[FemtoMips32.scala 459:31]
  assign core_io_mem_write_req_ready = router_io_coreReq_ready; // @[FemtoMips32.scala 461:31]
  assign router_clock = clock;
  assign router_reset = reset;
  assign router_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 463:11]
  assign router_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 463:11]
  assign router_io_next_ready = io_next_ready; // @[FemtoMips32.scala 464:11]
  assign router_io_coreReq_valid = core_io_mem_write_req_valid ? core_io_mem_write_req_valid :
    core_io_mem_read_req_valid; // @[FemtoMips32.scala 447:33]
  assign router_io_coreReq_bits_address = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_addr :
    core_io_mem_read_req_bits; // @[FemtoMips32.scala 448:40]
  assign router_io_coreReq_bits_data = core_io_mem_write_req_valid ? core_io_mem_write_req_bits_data : 32'h80; // @[FemtoMips32.scala 455:37]
  assign router_io_coreReq_bits_wen = core_io_mem_write_req_valid; // @[FemtoMips32.scala 453:31]
  assign router_io_coreResp_ready = core_io_mem_read_resp_ready; // @[FemtoMips32.scala 457:31]
endmodule
module MulticoreRing(
  input         clock,
  input         reset,
  output        io_prev_ready,
  input         io_prev_valid,
  input  [31:0] io_prev_bits_address,
  input  [31:0] io_prev_bits_data,
  input         io_prev_bits_wen,
  input  [7:0]  io_prev_bits_id,
  input         io_next_ready,
  output        io_next_valid,
  output [31:0] io_next_bits_address,
  output [31:0] io_next_bits_data,
  output        io_next_bits_wen,
  output [7:0]  io_next_bits_id,
  output        io_halted
);
  wire  cores_0_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_0_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_0_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_0_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_0_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_0_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_0_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_0_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_0_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_0_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_0_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_0_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_0_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_0_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_1_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_1_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_1_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_1_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_1_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_1_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_1_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_1_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_1_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_1_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_1_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_1_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_1_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_1_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_2_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_2_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_2_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_2_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_2_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_2_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_2_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_2_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_2_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_2_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_2_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_2_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_2_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_2_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_3_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_3_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_3_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_3_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_3_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_3_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_3_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_3_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_3_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_3_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_3_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_3_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_3_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_3_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_4_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_4_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_4_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_4_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_4_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_4_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_4_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_4_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_4_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_4_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_4_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_4_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_4_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_4_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_5_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_5_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_5_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_5_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_5_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_5_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_5_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_5_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_5_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_5_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_5_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_5_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_5_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_5_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_6_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_6_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_6_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_6_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_6_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_6_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_6_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_6_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_6_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_6_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_6_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_6_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_6_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_6_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_7_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_7_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_7_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_7_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_7_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_7_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_7_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_7_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_7_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_7_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_7_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_7_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_7_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_7_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_8_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_8_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_8_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_8_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_8_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_8_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_8_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_8_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_8_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_8_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_8_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_8_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_8_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_8_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_9_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_9_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_9_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_9_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_9_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_9_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_9_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_9_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_9_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_9_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_9_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_9_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_9_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_9_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_10_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_10_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_10_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_10_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_10_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_10_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_10_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_10_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_10_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_10_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_10_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_10_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_10_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_10_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_11_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_11_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_11_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_11_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_11_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_11_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_11_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_11_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_11_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_11_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_11_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_11_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_11_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_11_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_12_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_12_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_12_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_12_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_12_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_12_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_12_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_12_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_12_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_12_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_12_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_12_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_12_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_12_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_13_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_13_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_13_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_13_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_13_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_13_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_13_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_13_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_13_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_13_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_13_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_13_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_13_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_13_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_14_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_14_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_14_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_14_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_14_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_14_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_14_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_14_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_14_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_14_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_14_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_14_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_14_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_14_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_15_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_15_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_15_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_15_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_15_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_15_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_15_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_15_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_15_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_15_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_15_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_15_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_15_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_15_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_16_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_16_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_16_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_16_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_16_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_16_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_16_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_16_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_16_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_16_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_16_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_16_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_16_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_16_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_17_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_17_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_17_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_17_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_17_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_17_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_17_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_17_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_17_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_17_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_17_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_17_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_17_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_17_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_18_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_18_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_18_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_18_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_18_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_18_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_18_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_18_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_18_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_18_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_18_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_18_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_18_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_18_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_19_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_19_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_19_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_19_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_19_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_19_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_19_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_19_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_19_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_19_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_19_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_19_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_19_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_19_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_20_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_20_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_20_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_20_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_20_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_20_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_20_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_20_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_20_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_20_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_20_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_20_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_20_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_20_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_21_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_21_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_21_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_21_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_21_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_21_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_21_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_21_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_21_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_21_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_21_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_21_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_21_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_21_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_22_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_22_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_22_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_22_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_22_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_22_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_22_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_22_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_22_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_22_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_22_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_22_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_22_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_22_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_23_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_23_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_23_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_23_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_23_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_23_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_23_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_23_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_23_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_23_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_23_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_23_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_23_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_23_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_24_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_24_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_24_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_24_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_24_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_24_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_24_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_24_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_24_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_24_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_24_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_24_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_24_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_24_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_25_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_25_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_25_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_25_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_25_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_25_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_25_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_25_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_25_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_25_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_25_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_25_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_25_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_25_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_26_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_26_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_26_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_26_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_26_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_26_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_26_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_26_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_26_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_26_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_26_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_26_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_26_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_26_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_27_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_27_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_27_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_27_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_27_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_27_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_27_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_27_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_27_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_27_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_27_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_27_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_27_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_27_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_28_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_28_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_28_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_28_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_28_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_28_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_28_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_28_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_28_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_28_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_28_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_28_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_28_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_28_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_29_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_29_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_29_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_29_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_29_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_29_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_29_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_29_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_29_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_29_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_29_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_29_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_29_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_29_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_30_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_30_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_30_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_30_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_30_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_30_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_30_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_30_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_30_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_30_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_30_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_30_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_30_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_30_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_31_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_31_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_31_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_31_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_31_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_31_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_31_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_31_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_31_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_31_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_31_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_31_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_31_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_31_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_32_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_32_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_32_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_32_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_32_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_32_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_32_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_32_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_32_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_32_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_32_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_32_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_32_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_32_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_33_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_33_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_33_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_33_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_33_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_33_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_33_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_33_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_33_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_33_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_33_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_33_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_33_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_33_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_34_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_34_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_34_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_34_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_34_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_34_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_34_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_34_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_34_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_34_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_34_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_34_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_34_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_34_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_35_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_35_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_35_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_35_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_35_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_35_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_35_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_35_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_35_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_35_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_35_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_35_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_35_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_35_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_36_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_36_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_36_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_36_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_36_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_36_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_36_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_36_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_36_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_36_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_36_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_36_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_36_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_36_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_37_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_37_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_37_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_37_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_37_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_37_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_37_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_37_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_37_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_37_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_37_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_37_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_37_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_37_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_38_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_38_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_38_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_38_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_38_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_38_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_38_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_38_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_38_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_38_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_38_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_38_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_38_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_38_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_39_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_39_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_39_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_39_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_39_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_39_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_39_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_39_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_39_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_39_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_39_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_39_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_39_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_39_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_40_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_40_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_40_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_40_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_40_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_40_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_40_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_40_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_40_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_40_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_40_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_40_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_40_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_40_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_41_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_41_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_41_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_41_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_41_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_41_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_41_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_41_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_41_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_41_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_41_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_41_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_41_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_41_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_42_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_42_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_42_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_42_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_42_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_42_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_42_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_42_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_42_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_42_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_42_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_42_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_42_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_42_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_43_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_43_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_43_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_43_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_43_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_43_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_43_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_43_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_43_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_43_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_43_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_43_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_43_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_43_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_44_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_44_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_44_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_44_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_44_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_44_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_44_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_44_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_44_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_44_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_44_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_44_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_44_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_44_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_45_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_45_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_45_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_45_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_45_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_45_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_45_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_45_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_45_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_45_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_45_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_45_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_45_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_45_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_46_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_46_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_46_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_46_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_46_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_46_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_46_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_46_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_46_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_46_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_46_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_46_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_46_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_46_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_47_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_47_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_47_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_47_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_47_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_47_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_47_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_47_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_47_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_47_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_47_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_47_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_47_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_47_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_48_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_48_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_48_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_48_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_48_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_48_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_48_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_48_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_48_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_48_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_48_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_48_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_48_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_48_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_49_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_49_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_49_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_49_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_49_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_49_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_49_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_49_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_49_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_49_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_49_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_49_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_49_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_49_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_50_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_50_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_50_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_50_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_50_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_50_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_50_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_50_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_50_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_50_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_50_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_50_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_50_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_50_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_51_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_51_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_51_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_51_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_51_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_51_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_51_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_51_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_51_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_51_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_51_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_51_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_51_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_51_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_52_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_52_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_52_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_52_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_52_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_52_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_52_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_52_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_52_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_52_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_52_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_52_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_52_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_52_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_53_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_53_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_53_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_53_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_53_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_53_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_53_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_53_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_53_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_53_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_53_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_53_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_53_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_53_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_54_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_54_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_54_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_54_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_54_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_54_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_54_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_54_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_54_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_54_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_54_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_54_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_54_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_54_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_55_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_55_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_55_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_55_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_55_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_55_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_55_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_55_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_55_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_55_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_55_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_55_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_55_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_55_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_56_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_56_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_56_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_56_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_56_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_56_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_56_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_56_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_56_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_56_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_56_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_56_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_56_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_56_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_57_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_57_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_57_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_57_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_57_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_57_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_57_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_57_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_57_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_57_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_57_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_57_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_57_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_57_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_58_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_58_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_58_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_58_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_58_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_58_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_58_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_58_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_58_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_58_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_58_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_58_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_58_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_58_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_59_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_59_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_59_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_59_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_59_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_59_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_59_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_59_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_59_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_59_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_59_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_59_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_59_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_59_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_60_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_60_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_60_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_60_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_60_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_60_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_60_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_60_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_60_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_60_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_60_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_60_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_60_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_60_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_61_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_61_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_61_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_61_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_61_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_61_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_61_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_61_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_61_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_61_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_61_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_61_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_61_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_61_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_62_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_62_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_62_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_62_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_62_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_62_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_62_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_62_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_62_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_62_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_62_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_62_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_62_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_62_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_63_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_63_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_63_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_63_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_63_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_63_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_63_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_63_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_63_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_63_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_63_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_63_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_63_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_63_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_64_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_64_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_64_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_64_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_64_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_64_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_64_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_64_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_64_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_64_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_64_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_64_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_64_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_64_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_65_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_65_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_65_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_65_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_65_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_65_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_65_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_65_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_65_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_65_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_65_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_65_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_65_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_65_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_66_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_66_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_66_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_66_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_66_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_66_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_66_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_66_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_66_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_66_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_66_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_66_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_66_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_66_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_67_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_67_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_67_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_67_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_67_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_67_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_67_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_67_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_67_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_67_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_67_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_67_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_67_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_67_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_68_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_68_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_68_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_68_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_68_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_68_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_68_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_68_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_68_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_68_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_68_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_68_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_68_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_68_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_69_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_69_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_69_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_69_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_69_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_69_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_69_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_69_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_69_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_69_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_69_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_69_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_69_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_69_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_70_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_70_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_70_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_70_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_70_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_70_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_70_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_70_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_70_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_70_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_70_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_70_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_70_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_70_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_71_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_71_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_71_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_71_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_71_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_71_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_71_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_71_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_71_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_71_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_71_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_71_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_71_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_71_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_72_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_72_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_72_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_72_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_72_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_72_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_72_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_72_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_72_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_72_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_72_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_72_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_72_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_72_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_73_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_73_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_73_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_73_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_73_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_73_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_73_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_73_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_73_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_73_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_73_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_73_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_73_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_73_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_74_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_74_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_74_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_74_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_74_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_74_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_74_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_74_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_74_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_74_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_74_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_74_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_74_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_74_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_75_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_75_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_75_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_75_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_75_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_75_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_75_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_75_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_75_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_75_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_75_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_75_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_75_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_75_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_76_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_76_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_76_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_76_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_76_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_76_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_76_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_76_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_76_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_76_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_76_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_76_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_76_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_76_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_77_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_77_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_77_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_77_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_77_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_77_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_77_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_77_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_77_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_77_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_77_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_77_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_77_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_77_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_78_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_78_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_78_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_78_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_78_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_78_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_78_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_78_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_78_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_78_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_78_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_78_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_78_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_78_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_79_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_79_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_79_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_79_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_79_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_79_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_79_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_79_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_79_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_79_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_79_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_79_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_79_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_79_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_80_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_80_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_80_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_80_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_80_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_80_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_80_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_80_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_80_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_80_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_80_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_80_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_80_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_80_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_81_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_81_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_81_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_81_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_81_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_81_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_81_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_81_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_81_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_81_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_81_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_81_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_81_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_81_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_82_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_82_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_82_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_82_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_82_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_82_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_82_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_82_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_82_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_82_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_82_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_82_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_82_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_82_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_83_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_83_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_83_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_83_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_83_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_83_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_83_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_83_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_83_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_83_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_83_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_83_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_83_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_83_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_84_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_84_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_84_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_84_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_84_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_84_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_84_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_84_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_84_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_84_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_84_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_84_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_84_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_84_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_85_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_85_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_85_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_85_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_85_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_85_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_85_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_85_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_85_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_85_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_85_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_85_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_85_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_85_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_86_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_86_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_86_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_86_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_86_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_86_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_86_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_86_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_86_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_86_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_86_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_86_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_86_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_86_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_87_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_87_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_87_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_87_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_87_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_87_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_87_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_87_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_87_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_87_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_87_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_87_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_87_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_87_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_88_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_88_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_88_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_88_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_88_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_88_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_88_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_88_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_88_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_88_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_88_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_88_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_88_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_88_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_89_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_89_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_89_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_89_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_89_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_89_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_89_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_89_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_89_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_89_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_89_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_89_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_89_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_89_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_90_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_90_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_90_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_90_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_90_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_90_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_90_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_90_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_90_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_90_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_90_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_90_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_90_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_90_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_91_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_91_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_91_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_91_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_91_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_91_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_91_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_91_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_91_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_91_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_91_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_91_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_91_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_91_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_92_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_92_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_92_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_92_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_92_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_92_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_92_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_92_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_92_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_92_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_92_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_92_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_92_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_92_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_93_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_93_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_93_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_93_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_93_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_93_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_93_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_93_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_93_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_93_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_93_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_93_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_93_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_93_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_94_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_94_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_94_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_94_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_94_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_94_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_94_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_94_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_94_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_94_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_94_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_94_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_94_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_94_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_95_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_95_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_95_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_95_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_95_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_95_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_95_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_95_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_95_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_95_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_95_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_95_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_95_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_95_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_96_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_96_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_96_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_96_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_96_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_96_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_96_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_96_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_96_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_96_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_96_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_96_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_96_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_96_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_97_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_97_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_97_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_97_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_97_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_97_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_97_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_97_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_97_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_97_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_97_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_97_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_97_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_97_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_98_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_98_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_98_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_98_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_98_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_98_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_98_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_98_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_98_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_98_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_98_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_98_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_98_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_98_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_99_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_99_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_99_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_99_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_99_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_99_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_99_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_99_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_99_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_99_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_99_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_99_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_99_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_99_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_100_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_100_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_100_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_100_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_100_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_100_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_100_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_100_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_100_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_100_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_100_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_100_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_100_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_100_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_101_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_101_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_101_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_101_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_101_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_101_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_101_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_101_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_101_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_101_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_101_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_101_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_101_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_101_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_102_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_102_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_102_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_102_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_102_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_102_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_102_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_102_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_102_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_102_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_102_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_102_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_102_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_102_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_103_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_103_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_103_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_103_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_103_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_103_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_103_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_103_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_103_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_103_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_103_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_103_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_103_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_103_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_104_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_104_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_104_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_104_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_104_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_104_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_104_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_104_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_104_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_104_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_104_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_104_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_104_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_104_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_105_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_105_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_105_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_105_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_105_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_105_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_105_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_105_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_105_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_105_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_105_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_105_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_105_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_105_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_106_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_106_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_106_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_106_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_106_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_106_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_106_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_106_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_106_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_106_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_106_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_106_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_106_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_106_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_107_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_107_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_107_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_107_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_107_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_107_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_107_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_107_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_107_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_107_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_107_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_107_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_107_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_107_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_108_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_108_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_108_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_108_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_108_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_108_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_108_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_108_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_108_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_108_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_108_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_108_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_108_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_108_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_109_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_109_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_109_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_109_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_109_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_109_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_109_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_109_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_109_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_109_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_109_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_109_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_109_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_109_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_110_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_110_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_110_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_110_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_110_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_110_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_110_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_110_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_110_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_110_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_110_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_110_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_110_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_110_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_111_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_111_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_111_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_111_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_111_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_111_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_111_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_111_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_111_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_111_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_111_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_111_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_111_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_111_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_112_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_112_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_112_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_112_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_112_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_112_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_112_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_112_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_112_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_112_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_112_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_112_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_112_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_112_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_113_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_113_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_113_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_113_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_113_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_113_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_113_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_113_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_113_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_113_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_113_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_113_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_113_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_113_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_114_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_114_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_114_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_114_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_114_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_114_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_114_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_114_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_114_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_114_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_114_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_114_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_114_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_114_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_115_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_115_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_115_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_115_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_115_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_115_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_115_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_115_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_115_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_115_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_115_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_115_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_115_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_115_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_116_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_116_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_116_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_116_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_116_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_116_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_116_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_116_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_116_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_116_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_116_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_116_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_116_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_116_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_117_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_117_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_117_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_117_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_117_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_117_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_117_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_117_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_117_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_117_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_117_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_117_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_117_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_117_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_118_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_118_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_118_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_118_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_118_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_118_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_118_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_118_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_118_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_118_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_118_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_118_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_118_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_118_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_119_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_119_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_119_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_119_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_119_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_119_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_119_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_119_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_119_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_119_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_119_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_119_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_119_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_119_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_120_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_120_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_120_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_120_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_120_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_120_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_120_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_120_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_120_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_120_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_120_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_120_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_120_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_120_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_121_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_121_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_121_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_121_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_121_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_121_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_121_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_121_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_121_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_121_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_121_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_121_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_121_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_121_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_122_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_122_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_122_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_122_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_122_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_122_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_122_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_122_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_122_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_122_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_122_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_122_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_122_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_122_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_123_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_123_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_123_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_123_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_123_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_123_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_123_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_123_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_123_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_123_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_123_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_123_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_123_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_123_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_124_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_124_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_124_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_124_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_124_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_124_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_124_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_124_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_124_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_124_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_124_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_124_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_124_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_124_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_125_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_125_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_125_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_125_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_125_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_125_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_125_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_125_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_125_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_125_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_125_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_125_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_125_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_125_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_126_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_126_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_126_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_126_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_126_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_126_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_126_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_126_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_126_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_126_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_126_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_126_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_126_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_126_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_127_clock; // @[FemtoMips32.scala 470:51]
  wire  cores_127_reset; // @[FemtoMips32.scala 470:51]
  wire  cores_127_io_prev_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_127_io_prev_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_127_io_prev_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_127_io_prev_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_127_io_prev_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_127_io_prev_bits_id; // @[FemtoMips32.scala 470:51]
  wire  cores_127_io_next_ready; // @[FemtoMips32.scala 470:51]
  wire  cores_127_io_next_valid; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_127_io_next_bits_address; // @[FemtoMips32.scala 470:51]
  wire [31:0] cores_127_io_next_bits_data; // @[FemtoMips32.scala 470:51]
  wire  cores_127_io_next_bits_wen; // @[FemtoMips32.scala 470:51]
  wire [7:0] cores_127_io_next_bits_id; // @[FemtoMips32.scala 470:51]
  RingCore cores_0 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_0_clock),
    .reset(cores_0_reset),
    .io_prev_ready(cores_0_io_prev_ready),
    .io_prev_valid(cores_0_io_prev_valid),
    .io_prev_bits_address(cores_0_io_prev_bits_address),
    .io_prev_bits_data(cores_0_io_prev_bits_data),
    .io_prev_bits_wen(cores_0_io_prev_bits_wen),
    .io_prev_bits_id(cores_0_io_prev_bits_id),
    .io_next_ready(cores_0_io_next_ready),
    .io_next_valid(cores_0_io_next_valid),
    .io_next_bits_address(cores_0_io_next_bits_address),
    .io_next_bits_data(cores_0_io_next_bits_data),
    .io_next_bits_wen(cores_0_io_next_bits_wen),
    .io_next_bits_id(cores_0_io_next_bits_id)
  );
  RingCore_1 cores_1 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_1_clock),
    .reset(cores_1_reset),
    .io_prev_ready(cores_1_io_prev_ready),
    .io_prev_valid(cores_1_io_prev_valid),
    .io_prev_bits_address(cores_1_io_prev_bits_address),
    .io_prev_bits_data(cores_1_io_prev_bits_data),
    .io_prev_bits_wen(cores_1_io_prev_bits_wen),
    .io_prev_bits_id(cores_1_io_prev_bits_id),
    .io_next_ready(cores_1_io_next_ready),
    .io_next_valid(cores_1_io_next_valid),
    .io_next_bits_address(cores_1_io_next_bits_address),
    .io_next_bits_data(cores_1_io_next_bits_data),
    .io_next_bits_wen(cores_1_io_next_bits_wen),
    .io_next_bits_id(cores_1_io_next_bits_id)
  );
  RingCore_2 cores_2 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_2_clock),
    .reset(cores_2_reset),
    .io_prev_ready(cores_2_io_prev_ready),
    .io_prev_valid(cores_2_io_prev_valid),
    .io_prev_bits_address(cores_2_io_prev_bits_address),
    .io_prev_bits_data(cores_2_io_prev_bits_data),
    .io_prev_bits_wen(cores_2_io_prev_bits_wen),
    .io_prev_bits_id(cores_2_io_prev_bits_id),
    .io_next_ready(cores_2_io_next_ready),
    .io_next_valid(cores_2_io_next_valid),
    .io_next_bits_address(cores_2_io_next_bits_address),
    .io_next_bits_data(cores_2_io_next_bits_data),
    .io_next_bits_wen(cores_2_io_next_bits_wen),
    .io_next_bits_id(cores_2_io_next_bits_id)
  );
  RingCore_3 cores_3 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_3_clock),
    .reset(cores_3_reset),
    .io_prev_ready(cores_3_io_prev_ready),
    .io_prev_valid(cores_3_io_prev_valid),
    .io_prev_bits_address(cores_3_io_prev_bits_address),
    .io_prev_bits_data(cores_3_io_prev_bits_data),
    .io_prev_bits_wen(cores_3_io_prev_bits_wen),
    .io_prev_bits_id(cores_3_io_prev_bits_id),
    .io_next_ready(cores_3_io_next_ready),
    .io_next_valid(cores_3_io_next_valid),
    .io_next_bits_address(cores_3_io_next_bits_address),
    .io_next_bits_data(cores_3_io_next_bits_data),
    .io_next_bits_wen(cores_3_io_next_bits_wen),
    .io_next_bits_id(cores_3_io_next_bits_id)
  );
  RingCore_4 cores_4 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_4_clock),
    .reset(cores_4_reset),
    .io_prev_ready(cores_4_io_prev_ready),
    .io_prev_valid(cores_4_io_prev_valid),
    .io_prev_bits_address(cores_4_io_prev_bits_address),
    .io_prev_bits_data(cores_4_io_prev_bits_data),
    .io_prev_bits_wen(cores_4_io_prev_bits_wen),
    .io_prev_bits_id(cores_4_io_prev_bits_id),
    .io_next_ready(cores_4_io_next_ready),
    .io_next_valid(cores_4_io_next_valid),
    .io_next_bits_address(cores_4_io_next_bits_address),
    .io_next_bits_data(cores_4_io_next_bits_data),
    .io_next_bits_wen(cores_4_io_next_bits_wen),
    .io_next_bits_id(cores_4_io_next_bits_id)
  );
  RingCore_5 cores_5 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_5_clock),
    .reset(cores_5_reset),
    .io_prev_ready(cores_5_io_prev_ready),
    .io_prev_valid(cores_5_io_prev_valid),
    .io_prev_bits_address(cores_5_io_prev_bits_address),
    .io_prev_bits_data(cores_5_io_prev_bits_data),
    .io_prev_bits_wen(cores_5_io_prev_bits_wen),
    .io_prev_bits_id(cores_5_io_prev_bits_id),
    .io_next_ready(cores_5_io_next_ready),
    .io_next_valid(cores_5_io_next_valid),
    .io_next_bits_address(cores_5_io_next_bits_address),
    .io_next_bits_data(cores_5_io_next_bits_data),
    .io_next_bits_wen(cores_5_io_next_bits_wen),
    .io_next_bits_id(cores_5_io_next_bits_id)
  );
  RingCore_6 cores_6 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_6_clock),
    .reset(cores_6_reset),
    .io_prev_ready(cores_6_io_prev_ready),
    .io_prev_valid(cores_6_io_prev_valid),
    .io_prev_bits_address(cores_6_io_prev_bits_address),
    .io_prev_bits_data(cores_6_io_prev_bits_data),
    .io_prev_bits_wen(cores_6_io_prev_bits_wen),
    .io_prev_bits_id(cores_6_io_prev_bits_id),
    .io_next_ready(cores_6_io_next_ready),
    .io_next_valid(cores_6_io_next_valid),
    .io_next_bits_address(cores_6_io_next_bits_address),
    .io_next_bits_data(cores_6_io_next_bits_data),
    .io_next_bits_wen(cores_6_io_next_bits_wen),
    .io_next_bits_id(cores_6_io_next_bits_id)
  );
  RingCore_7 cores_7 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_7_clock),
    .reset(cores_7_reset),
    .io_prev_ready(cores_7_io_prev_ready),
    .io_prev_valid(cores_7_io_prev_valid),
    .io_prev_bits_address(cores_7_io_prev_bits_address),
    .io_prev_bits_data(cores_7_io_prev_bits_data),
    .io_prev_bits_wen(cores_7_io_prev_bits_wen),
    .io_prev_bits_id(cores_7_io_prev_bits_id),
    .io_next_ready(cores_7_io_next_ready),
    .io_next_valid(cores_7_io_next_valid),
    .io_next_bits_address(cores_7_io_next_bits_address),
    .io_next_bits_data(cores_7_io_next_bits_data),
    .io_next_bits_wen(cores_7_io_next_bits_wen),
    .io_next_bits_id(cores_7_io_next_bits_id)
  );
  RingCore_8 cores_8 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_8_clock),
    .reset(cores_8_reset),
    .io_prev_ready(cores_8_io_prev_ready),
    .io_prev_valid(cores_8_io_prev_valid),
    .io_prev_bits_address(cores_8_io_prev_bits_address),
    .io_prev_bits_data(cores_8_io_prev_bits_data),
    .io_prev_bits_wen(cores_8_io_prev_bits_wen),
    .io_prev_bits_id(cores_8_io_prev_bits_id),
    .io_next_ready(cores_8_io_next_ready),
    .io_next_valid(cores_8_io_next_valid),
    .io_next_bits_address(cores_8_io_next_bits_address),
    .io_next_bits_data(cores_8_io_next_bits_data),
    .io_next_bits_wen(cores_8_io_next_bits_wen),
    .io_next_bits_id(cores_8_io_next_bits_id)
  );
  RingCore_9 cores_9 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_9_clock),
    .reset(cores_9_reset),
    .io_prev_ready(cores_9_io_prev_ready),
    .io_prev_valid(cores_9_io_prev_valid),
    .io_prev_bits_address(cores_9_io_prev_bits_address),
    .io_prev_bits_data(cores_9_io_prev_bits_data),
    .io_prev_bits_wen(cores_9_io_prev_bits_wen),
    .io_prev_bits_id(cores_9_io_prev_bits_id),
    .io_next_ready(cores_9_io_next_ready),
    .io_next_valid(cores_9_io_next_valid),
    .io_next_bits_address(cores_9_io_next_bits_address),
    .io_next_bits_data(cores_9_io_next_bits_data),
    .io_next_bits_wen(cores_9_io_next_bits_wen),
    .io_next_bits_id(cores_9_io_next_bits_id)
  );
  RingCore_10 cores_10 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_10_clock),
    .reset(cores_10_reset),
    .io_prev_ready(cores_10_io_prev_ready),
    .io_prev_valid(cores_10_io_prev_valid),
    .io_prev_bits_address(cores_10_io_prev_bits_address),
    .io_prev_bits_data(cores_10_io_prev_bits_data),
    .io_prev_bits_wen(cores_10_io_prev_bits_wen),
    .io_prev_bits_id(cores_10_io_prev_bits_id),
    .io_next_ready(cores_10_io_next_ready),
    .io_next_valid(cores_10_io_next_valid),
    .io_next_bits_address(cores_10_io_next_bits_address),
    .io_next_bits_data(cores_10_io_next_bits_data),
    .io_next_bits_wen(cores_10_io_next_bits_wen),
    .io_next_bits_id(cores_10_io_next_bits_id)
  );
  RingCore_11 cores_11 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_11_clock),
    .reset(cores_11_reset),
    .io_prev_ready(cores_11_io_prev_ready),
    .io_prev_valid(cores_11_io_prev_valid),
    .io_prev_bits_address(cores_11_io_prev_bits_address),
    .io_prev_bits_data(cores_11_io_prev_bits_data),
    .io_prev_bits_wen(cores_11_io_prev_bits_wen),
    .io_prev_bits_id(cores_11_io_prev_bits_id),
    .io_next_ready(cores_11_io_next_ready),
    .io_next_valid(cores_11_io_next_valid),
    .io_next_bits_address(cores_11_io_next_bits_address),
    .io_next_bits_data(cores_11_io_next_bits_data),
    .io_next_bits_wen(cores_11_io_next_bits_wen),
    .io_next_bits_id(cores_11_io_next_bits_id)
  );
  RingCore_12 cores_12 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_12_clock),
    .reset(cores_12_reset),
    .io_prev_ready(cores_12_io_prev_ready),
    .io_prev_valid(cores_12_io_prev_valid),
    .io_prev_bits_address(cores_12_io_prev_bits_address),
    .io_prev_bits_data(cores_12_io_prev_bits_data),
    .io_prev_bits_wen(cores_12_io_prev_bits_wen),
    .io_prev_bits_id(cores_12_io_prev_bits_id),
    .io_next_ready(cores_12_io_next_ready),
    .io_next_valid(cores_12_io_next_valid),
    .io_next_bits_address(cores_12_io_next_bits_address),
    .io_next_bits_data(cores_12_io_next_bits_data),
    .io_next_bits_wen(cores_12_io_next_bits_wen),
    .io_next_bits_id(cores_12_io_next_bits_id)
  );
  RingCore_13 cores_13 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_13_clock),
    .reset(cores_13_reset),
    .io_prev_ready(cores_13_io_prev_ready),
    .io_prev_valid(cores_13_io_prev_valid),
    .io_prev_bits_address(cores_13_io_prev_bits_address),
    .io_prev_bits_data(cores_13_io_prev_bits_data),
    .io_prev_bits_wen(cores_13_io_prev_bits_wen),
    .io_prev_bits_id(cores_13_io_prev_bits_id),
    .io_next_ready(cores_13_io_next_ready),
    .io_next_valid(cores_13_io_next_valid),
    .io_next_bits_address(cores_13_io_next_bits_address),
    .io_next_bits_data(cores_13_io_next_bits_data),
    .io_next_bits_wen(cores_13_io_next_bits_wen),
    .io_next_bits_id(cores_13_io_next_bits_id)
  );
  RingCore_14 cores_14 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_14_clock),
    .reset(cores_14_reset),
    .io_prev_ready(cores_14_io_prev_ready),
    .io_prev_valid(cores_14_io_prev_valid),
    .io_prev_bits_address(cores_14_io_prev_bits_address),
    .io_prev_bits_data(cores_14_io_prev_bits_data),
    .io_prev_bits_wen(cores_14_io_prev_bits_wen),
    .io_prev_bits_id(cores_14_io_prev_bits_id),
    .io_next_ready(cores_14_io_next_ready),
    .io_next_valid(cores_14_io_next_valid),
    .io_next_bits_address(cores_14_io_next_bits_address),
    .io_next_bits_data(cores_14_io_next_bits_data),
    .io_next_bits_wen(cores_14_io_next_bits_wen),
    .io_next_bits_id(cores_14_io_next_bits_id)
  );
  RingCore_15 cores_15 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_15_clock),
    .reset(cores_15_reset),
    .io_prev_ready(cores_15_io_prev_ready),
    .io_prev_valid(cores_15_io_prev_valid),
    .io_prev_bits_address(cores_15_io_prev_bits_address),
    .io_prev_bits_data(cores_15_io_prev_bits_data),
    .io_prev_bits_wen(cores_15_io_prev_bits_wen),
    .io_prev_bits_id(cores_15_io_prev_bits_id),
    .io_next_ready(cores_15_io_next_ready),
    .io_next_valid(cores_15_io_next_valid),
    .io_next_bits_address(cores_15_io_next_bits_address),
    .io_next_bits_data(cores_15_io_next_bits_data),
    .io_next_bits_wen(cores_15_io_next_bits_wen),
    .io_next_bits_id(cores_15_io_next_bits_id)
  );
  RingCore_16 cores_16 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_16_clock),
    .reset(cores_16_reset),
    .io_prev_ready(cores_16_io_prev_ready),
    .io_prev_valid(cores_16_io_prev_valid),
    .io_prev_bits_address(cores_16_io_prev_bits_address),
    .io_prev_bits_data(cores_16_io_prev_bits_data),
    .io_prev_bits_wen(cores_16_io_prev_bits_wen),
    .io_prev_bits_id(cores_16_io_prev_bits_id),
    .io_next_ready(cores_16_io_next_ready),
    .io_next_valid(cores_16_io_next_valid),
    .io_next_bits_address(cores_16_io_next_bits_address),
    .io_next_bits_data(cores_16_io_next_bits_data),
    .io_next_bits_wen(cores_16_io_next_bits_wen),
    .io_next_bits_id(cores_16_io_next_bits_id)
  );
  RingCore_17 cores_17 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_17_clock),
    .reset(cores_17_reset),
    .io_prev_ready(cores_17_io_prev_ready),
    .io_prev_valid(cores_17_io_prev_valid),
    .io_prev_bits_address(cores_17_io_prev_bits_address),
    .io_prev_bits_data(cores_17_io_prev_bits_data),
    .io_prev_bits_wen(cores_17_io_prev_bits_wen),
    .io_prev_bits_id(cores_17_io_prev_bits_id),
    .io_next_ready(cores_17_io_next_ready),
    .io_next_valid(cores_17_io_next_valid),
    .io_next_bits_address(cores_17_io_next_bits_address),
    .io_next_bits_data(cores_17_io_next_bits_data),
    .io_next_bits_wen(cores_17_io_next_bits_wen),
    .io_next_bits_id(cores_17_io_next_bits_id)
  );
  RingCore_18 cores_18 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_18_clock),
    .reset(cores_18_reset),
    .io_prev_ready(cores_18_io_prev_ready),
    .io_prev_valid(cores_18_io_prev_valid),
    .io_prev_bits_address(cores_18_io_prev_bits_address),
    .io_prev_bits_data(cores_18_io_prev_bits_data),
    .io_prev_bits_wen(cores_18_io_prev_bits_wen),
    .io_prev_bits_id(cores_18_io_prev_bits_id),
    .io_next_ready(cores_18_io_next_ready),
    .io_next_valid(cores_18_io_next_valid),
    .io_next_bits_address(cores_18_io_next_bits_address),
    .io_next_bits_data(cores_18_io_next_bits_data),
    .io_next_bits_wen(cores_18_io_next_bits_wen),
    .io_next_bits_id(cores_18_io_next_bits_id)
  );
  RingCore_19 cores_19 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_19_clock),
    .reset(cores_19_reset),
    .io_prev_ready(cores_19_io_prev_ready),
    .io_prev_valid(cores_19_io_prev_valid),
    .io_prev_bits_address(cores_19_io_prev_bits_address),
    .io_prev_bits_data(cores_19_io_prev_bits_data),
    .io_prev_bits_wen(cores_19_io_prev_bits_wen),
    .io_prev_bits_id(cores_19_io_prev_bits_id),
    .io_next_ready(cores_19_io_next_ready),
    .io_next_valid(cores_19_io_next_valid),
    .io_next_bits_address(cores_19_io_next_bits_address),
    .io_next_bits_data(cores_19_io_next_bits_data),
    .io_next_bits_wen(cores_19_io_next_bits_wen),
    .io_next_bits_id(cores_19_io_next_bits_id)
  );
  RingCore_20 cores_20 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_20_clock),
    .reset(cores_20_reset),
    .io_prev_ready(cores_20_io_prev_ready),
    .io_prev_valid(cores_20_io_prev_valid),
    .io_prev_bits_address(cores_20_io_prev_bits_address),
    .io_prev_bits_data(cores_20_io_prev_bits_data),
    .io_prev_bits_wen(cores_20_io_prev_bits_wen),
    .io_prev_bits_id(cores_20_io_prev_bits_id),
    .io_next_ready(cores_20_io_next_ready),
    .io_next_valid(cores_20_io_next_valid),
    .io_next_bits_address(cores_20_io_next_bits_address),
    .io_next_bits_data(cores_20_io_next_bits_data),
    .io_next_bits_wen(cores_20_io_next_bits_wen),
    .io_next_bits_id(cores_20_io_next_bits_id)
  );
  RingCore_21 cores_21 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_21_clock),
    .reset(cores_21_reset),
    .io_prev_ready(cores_21_io_prev_ready),
    .io_prev_valid(cores_21_io_prev_valid),
    .io_prev_bits_address(cores_21_io_prev_bits_address),
    .io_prev_bits_data(cores_21_io_prev_bits_data),
    .io_prev_bits_wen(cores_21_io_prev_bits_wen),
    .io_prev_bits_id(cores_21_io_prev_bits_id),
    .io_next_ready(cores_21_io_next_ready),
    .io_next_valid(cores_21_io_next_valid),
    .io_next_bits_address(cores_21_io_next_bits_address),
    .io_next_bits_data(cores_21_io_next_bits_data),
    .io_next_bits_wen(cores_21_io_next_bits_wen),
    .io_next_bits_id(cores_21_io_next_bits_id)
  );
  RingCore_22 cores_22 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_22_clock),
    .reset(cores_22_reset),
    .io_prev_ready(cores_22_io_prev_ready),
    .io_prev_valid(cores_22_io_prev_valid),
    .io_prev_bits_address(cores_22_io_prev_bits_address),
    .io_prev_bits_data(cores_22_io_prev_bits_data),
    .io_prev_bits_wen(cores_22_io_prev_bits_wen),
    .io_prev_bits_id(cores_22_io_prev_bits_id),
    .io_next_ready(cores_22_io_next_ready),
    .io_next_valid(cores_22_io_next_valid),
    .io_next_bits_address(cores_22_io_next_bits_address),
    .io_next_bits_data(cores_22_io_next_bits_data),
    .io_next_bits_wen(cores_22_io_next_bits_wen),
    .io_next_bits_id(cores_22_io_next_bits_id)
  );
  RingCore_23 cores_23 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_23_clock),
    .reset(cores_23_reset),
    .io_prev_ready(cores_23_io_prev_ready),
    .io_prev_valid(cores_23_io_prev_valid),
    .io_prev_bits_address(cores_23_io_prev_bits_address),
    .io_prev_bits_data(cores_23_io_prev_bits_data),
    .io_prev_bits_wen(cores_23_io_prev_bits_wen),
    .io_prev_bits_id(cores_23_io_prev_bits_id),
    .io_next_ready(cores_23_io_next_ready),
    .io_next_valid(cores_23_io_next_valid),
    .io_next_bits_address(cores_23_io_next_bits_address),
    .io_next_bits_data(cores_23_io_next_bits_data),
    .io_next_bits_wen(cores_23_io_next_bits_wen),
    .io_next_bits_id(cores_23_io_next_bits_id)
  );
  RingCore_24 cores_24 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_24_clock),
    .reset(cores_24_reset),
    .io_prev_ready(cores_24_io_prev_ready),
    .io_prev_valid(cores_24_io_prev_valid),
    .io_prev_bits_address(cores_24_io_prev_bits_address),
    .io_prev_bits_data(cores_24_io_prev_bits_data),
    .io_prev_bits_wen(cores_24_io_prev_bits_wen),
    .io_prev_bits_id(cores_24_io_prev_bits_id),
    .io_next_ready(cores_24_io_next_ready),
    .io_next_valid(cores_24_io_next_valid),
    .io_next_bits_address(cores_24_io_next_bits_address),
    .io_next_bits_data(cores_24_io_next_bits_data),
    .io_next_bits_wen(cores_24_io_next_bits_wen),
    .io_next_bits_id(cores_24_io_next_bits_id)
  );
  RingCore_25 cores_25 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_25_clock),
    .reset(cores_25_reset),
    .io_prev_ready(cores_25_io_prev_ready),
    .io_prev_valid(cores_25_io_prev_valid),
    .io_prev_bits_address(cores_25_io_prev_bits_address),
    .io_prev_bits_data(cores_25_io_prev_bits_data),
    .io_prev_bits_wen(cores_25_io_prev_bits_wen),
    .io_prev_bits_id(cores_25_io_prev_bits_id),
    .io_next_ready(cores_25_io_next_ready),
    .io_next_valid(cores_25_io_next_valid),
    .io_next_bits_address(cores_25_io_next_bits_address),
    .io_next_bits_data(cores_25_io_next_bits_data),
    .io_next_bits_wen(cores_25_io_next_bits_wen),
    .io_next_bits_id(cores_25_io_next_bits_id)
  );
  RingCore_26 cores_26 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_26_clock),
    .reset(cores_26_reset),
    .io_prev_ready(cores_26_io_prev_ready),
    .io_prev_valid(cores_26_io_prev_valid),
    .io_prev_bits_address(cores_26_io_prev_bits_address),
    .io_prev_bits_data(cores_26_io_prev_bits_data),
    .io_prev_bits_wen(cores_26_io_prev_bits_wen),
    .io_prev_bits_id(cores_26_io_prev_bits_id),
    .io_next_ready(cores_26_io_next_ready),
    .io_next_valid(cores_26_io_next_valid),
    .io_next_bits_address(cores_26_io_next_bits_address),
    .io_next_bits_data(cores_26_io_next_bits_data),
    .io_next_bits_wen(cores_26_io_next_bits_wen),
    .io_next_bits_id(cores_26_io_next_bits_id)
  );
  RingCore_27 cores_27 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_27_clock),
    .reset(cores_27_reset),
    .io_prev_ready(cores_27_io_prev_ready),
    .io_prev_valid(cores_27_io_prev_valid),
    .io_prev_bits_address(cores_27_io_prev_bits_address),
    .io_prev_bits_data(cores_27_io_prev_bits_data),
    .io_prev_bits_wen(cores_27_io_prev_bits_wen),
    .io_prev_bits_id(cores_27_io_prev_bits_id),
    .io_next_ready(cores_27_io_next_ready),
    .io_next_valid(cores_27_io_next_valid),
    .io_next_bits_address(cores_27_io_next_bits_address),
    .io_next_bits_data(cores_27_io_next_bits_data),
    .io_next_bits_wen(cores_27_io_next_bits_wen),
    .io_next_bits_id(cores_27_io_next_bits_id)
  );
  RingCore_28 cores_28 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_28_clock),
    .reset(cores_28_reset),
    .io_prev_ready(cores_28_io_prev_ready),
    .io_prev_valid(cores_28_io_prev_valid),
    .io_prev_bits_address(cores_28_io_prev_bits_address),
    .io_prev_bits_data(cores_28_io_prev_bits_data),
    .io_prev_bits_wen(cores_28_io_prev_bits_wen),
    .io_prev_bits_id(cores_28_io_prev_bits_id),
    .io_next_ready(cores_28_io_next_ready),
    .io_next_valid(cores_28_io_next_valid),
    .io_next_bits_address(cores_28_io_next_bits_address),
    .io_next_bits_data(cores_28_io_next_bits_data),
    .io_next_bits_wen(cores_28_io_next_bits_wen),
    .io_next_bits_id(cores_28_io_next_bits_id)
  );
  RingCore_29 cores_29 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_29_clock),
    .reset(cores_29_reset),
    .io_prev_ready(cores_29_io_prev_ready),
    .io_prev_valid(cores_29_io_prev_valid),
    .io_prev_bits_address(cores_29_io_prev_bits_address),
    .io_prev_bits_data(cores_29_io_prev_bits_data),
    .io_prev_bits_wen(cores_29_io_prev_bits_wen),
    .io_prev_bits_id(cores_29_io_prev_bits_id),
    .io_next_ready(cores_29_io_next_ready),
    .io_next_valid(cores_29_io_next_valid),
    .io_next_bits_address(cores_29_io_next_bits_address),
    .io_next_bits_data(cores_29_io_next_bits_data),
    .io_next_bits_wen(cores_29_io_next_bits_wen),
    .io_next_bits_id(cores_29_io_next_bits_id)
  );
  RingCore_30 cores_30 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_30_clock),
    .reset(cores_30_reset),
    .io_prev_ready(cores_30_io_prev_ready),
    .io_prev_valid(cores_30_io_prev_valid),
    .io_prev_bits_address(cores_30_io_prev_bits_address),
    .io_prev_bits_data(cores_30_io_prev_bits_data),
    .io_prev_bits_wen(cores_30_io_prev_bits_wen),
    .io_prev_bits_id(cores_30_io_prev_bits_id),
    .io_next_ready(cores_30_io_next_ready),
    .io_next_valid(cores_30_io_next_valid),
    .io_next_bits_address(cores_30_io_next_bits_address),
    .io_next_bits_data(cores_30_io_next_bits_data),
    .io_next_bits_wen(cores_30_io_next_bits_wen),
    .io_next_bits_id(cores_30_io_next_bits_id)
  );
  RingCore_31 cores_31 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_31_clock),
    .reset(cores_31_reset),
    .io_prev_ready(cores_31_io_prev_ready),
    .io_prev_valid(cores_31_io_prev_valid),
    .io_prev_bits_address(cores_31_io_prev_bits_address),
    .io_prev_bits_data(cores_31_io_prev_bits_data),
    .io_prev_bits_wen(cores_31_io_prev_bits_wen),
    .io_prev_bits_id(cores_31_io_prev_bits_id),
    .io_next_ready(cores_31_io_next_ready),
    .io_next_valid(cores_31_io_next_valid),
    .io_next_bits_address(cores_31_io_next_bits_address),
    .io_next_bits_data(cores_31_io_next_bits_data),
    .io_next_bits_wen(cores_31_io_next_bits_wen),
    .io_next_bits_id(cores_31_io_next_bits_id)
  );
  RingCore_32 cores_32 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_32_clock),
    .reset(cores_32_reset),
    .io_prev_ready(cores_32_io_prev_ready),
    .io_prev_valid(cores_32_io_prev_valid),
    .io_prev_bits_address(cores_32_io_prev_bits_address),
    .io_prev_bits_data(cores_32_io_prev_bits_data),
    .io_prev_bits_wen(cores_32_io_prev_bits_wen),
    .io_prev_bits_id(cores_32_io_prev_bits_id),
    .io_next_ready(cores_32_io_next_ready),
    .io_next_valid(cores_32_io_next_valid),
    .io_next_bits_address(cores_32_io_next_bits_address),
    .io_next_bits_data(cores_32_io_next_bits_data),
    .io_next_bits_wen(cores_32_io_next_bits_wen),
    .io_next_bits_id(cores_32_io_next_bits_id)
  );
  RingCore_33 cores_33 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_33_clock),
    .reset(cores_33_reset),
    .io_prev_ready(cores_33_io_prev_ready),
    .io_prev_valid(cores_33_io_prev_valid),
    .io_prev_bits_address(cores_33_io_prev_bits_address),
    .io_prev_bits_data(cores_33_io_prev_bits_data),
    .io_prev_bits_wen(cores_33_io_prev_bits_wen),
    .io_prev_bits_id(cores_33_io_prev_bits_id),
    .io_next_ready(cores_33_io_next_ready),
    .io_next_valid(cores_33_io_next_valid),
    .io_next_bits_address(cores_33_io_next_bits_address),
    .io_next_bits_data(cores_33_io_next_bits_data),
    .io_next_bits_wen(cores_33_io_next_bits_wen),
    .io_next_bits_id(cores_33_io_next_bits_id)
  );
  RingCore_34 cores_34 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_34_clock),
    .reset(cores_34_reset),
    .io_prev_ready(cores_34_io_prev_ready),
    .io_prev_valid(cores_34_io_prev_valid),
    .io_prev_bits_address(cores_34_io_prev_bits_address),
    .io_prev_bits_data(cores_34_io_prev_bits_data),
    .io_prev_bits_wen(cores_34_io_prev_bits_wen),
    .io_prev_bits_id(cores_34_io_prev_bits_id),
    .io_next_ready(cores_34_io_next_ready),
    .io_next_valid(cores_34_io_next_valid),
    .io_next_bits_address(cores_34_io_next_bits_address),
    .io_next_bits_data(cores_34_io_next_bits_data),
    .io_next_bits_wen(cores_34_io_next_bits_wen),
    .io_next_bits_id(cores_34_io_next_bits_id)
  );
  RingCore_35 cores_35 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_35_clock),
    .reset(cores_35_reset),
    .io_prev_ready(cores_35_io_prev_ready),
    .io_prev_valid(cores_35_io_prev_valid),
    .io_prev_bits_address(cores_35_io_prev_bits_address),
    .io_prev_bits_data(cores_35_io_prev_bits_data),
    .io_prev_bits_wen(cores_35_io_prev_bits_wen),
    .io_prev_bits_id(cores_35_io_prev_bits_id),
    .io_next_ready(cores_35_io_next_ready),
    .io_next_valid(cores_35_io_next_valid),
    .io_next_bits_address(cores_35_io_next_bits_address),
    .io_next_bits_data(cores_35_io_next_bits_data),
    .io_next_bits_wen(cores_35_io_next_bits_wen),
    .io_next_bits_id(cores_35_io_next_bits_id)
  );
  RingCore_36 cores_36 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_36_clock),
    .reset(cores_36_reset),
    .io_prev_ready(cores_36_io_prev_ready),
    .io_prev_valid(cores_36_io_prev_valid),
    .io_prev_bits_address(cores_36_io_prev_bits_address),
    .io_prev_bits_data(cores_36_io_prev_bits_data),
    .io_prev_bits_wen(cores_36_io_prev_bits_wen),
    .io_prev_bits_id(cores_36_io_prev_bits_id),
    .io_next_ready(cores_36_io_next_ready),
    .io_next_valid(cores_36_io_next_valid),
    .io_next_bits_address(cores_36_io_next_bits_address),
    .io_next_bits_data(cores_36_io_next_bits_data),
    .io_next_bits_wen(cores_36_io_next_bits_wen),
    .io_next_bits_id(cores_36_io_next_bits_id)
  );
  RingCore_37 cores_37 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_37_clock),
    .reset(cores_37_reset),
    .io_prev_ready(cores_37_io_prev_ready),
    .io_prev_valid(cores_37_io_prev_valid),
    .io_prev_bits_address(cores_37_io_prev_bits_address),
    .io_prev_bits_data(cores_37_io_prev_bits_data),
    .io_prev_bits_wen(cores_37_io_prev_bits_wen),
    .io_prev_bits_id(cores_37_io_prev_bits_id),
    .io_next_ready(cores_37_io_next_ready),
    .io_next_valid(cores_37_io_next_valid),
    .io_next_bits_address(cores_37_io_next_bits_address),
    .io_next_bits_data(cores_37_io_next_bits_data),
    .io_next_bits_wen(cores_37_io_next_bits_wen),
    .io_next_bits_id(cores_37_io_next_bits_id)
  );
  RingCore_38 cores_38 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_38_clock),
    .reset(cores_38_reset),
    .io_prev_ready(cores_38_io_prev_ready),
    .io_prev_valid(cores_38_io_prev_valid),
    .io_prev_bits_address(cores_38_io_prev_bits_address),
    .io_prev_bits_data(cores_38_io_prev_bits_data),
    .io_prev_bits_wen(cores_38_io_prev_bits_wen),
    .io_prev_bits_id(cores_38_io_prev_bits_id),
    .io_next_ready(cores_38_io_next_ready),
    .io_next_valid(cores_38_io_next_valid),
    .io_next_bits_address(cores_38_io_next_bits_address),
    .io_next_bits_data(cores_38_io_next_bits_data),
    .io_next_bits_wen(cores_38_io_next_bits_wen),
    .io_next_bits_id(cores_38_io_next_bits_id)
  );
  RingCore_39 cores_39 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_39_clock),
    .reset(cores_39_reset),
    .io_prev_ready(cores_39_io_prev_ready),
    .io_prev_valid(cores_39_io_prev_valid),
    .io_prev_bits_address(cores_39_io_prev_bits_address),
    .io_prev_bits_data(cores_39_io_prev_bits_data),
    .io_prev_bits_wen(cores_39_io_prev_bits_wen),
    .io_prev_bits_id(cores_39_io_prev_bits_id),
    .io_next_ready(cores_39_io_next_ready),
    .io_next_valid(cores_39_io_next_valid),
    .io_next_bits_address(cores_39_io_next_bits_address),
    .io_next_bits_data(cores_39_io_next_bits_data),
    .io_next_bits_wen(cores_39_io_next_bits_wen),
    .io_next_bits_id(cores_39_io_next_bits_id)
  );
  RingCore_40 cores_40 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_40_clock),
    .reset(cores_40_reset),
    .io_prev_ready(cores_40_io_prev_ready),
    .io_prev_valid(cores_40_io_prev_valid),
    .io_prev_bits_address(cores_40_io_prev_bits_address),
    .io_prev_bits_data(cores_40_io_prev_bits_data),
    .io_prev_bits_wen(cores_40_io_prev_bits_wen),
    .io_prev_bits_id(cores_40_io_prev_bits_id),
    .io_next_ready(cores_40_io_next_ready),
    .io_next_valid(cores_40_io_next_valid),
    .io_next_bits_address(cores_40_io_next_bits_address),
    .io_next_bits_data(cores_40_io_next_bits_data),
    .io_next_bits_wen(cores_40_io_next_bits_wen),
    .io_next_bits_id(cores_40_io_next_bits_id)
  );
  RingCore_41 cores_41 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_41_clock),
    .reset(cores_41_reset),
    .io_prev_ready(cores_41_io_prev_ready),
    .io_prev_valid(cores_41_io_prev_valid),
    .io_prev_bits_address(cores_41_io_prev_bits_address),
    .io_prev_bits_data(cores_41_io_prev_bits_data),
    .io_prev_bits_wen(cores_41_io_prev_bits_wen),
    .io_prev_bits_id(cores_41_io_prev_bits_id),
    .io_next_ready(cores_41_io_next_ready),
    .io_next_valid(cores_41_io_next_valid),
    .io_next_bits_address(cores_41_io_next_bits_address),
    .io_next_bits_data(cores_41_io_next_bits_data),
    .io_next_bits_wen(cores_41_io_next_bits_wen),
    .io_next_bits_id(cores_41_io_next_bits_id)
  );
  RingCore_42 cores_42 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_42_clock),
    .reset(cores_42_reset),
    .io_prev_ready(cores_42_io_prev_ready),
    .io_prev_valid(cores_42_io_prev_valid),
    .io_prev_bits_address(cores_42_io_prev_bits_address),
    .io_prev_bits_data(cores_42_io_prev_bits_data),
    .io_prev_bits_wen(cores_42_io_prev_bits_wen),
    .io_prev_bits_id(cores_42_io_prev_bits_id),
    .io_next_ready(cores_42_io_next_ready),
    .io_next_valid(cores_42_io_next_valid),
    .io_next_bits_address(cores_42_io_next_bits_address),
    .io_next_bits_data(cores_42_io_next_bits_data),
    .io_next_bits_wen(cores_42_io_next_bits_wen),
    .io_next_bits_id(cores_42_io_next_bits_id)
  );
  RingCore_43 cores_43 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_43_clock),
    .reset(cores_43_reset),
    .io_prev_ready(cores_43_io_prev_ready),
    .io_prev_valid(cores_43_io_prev_valid),
    .io_prev_bits_address(cores_43_io_prev_bits_address),
    .io_prev_bits_data(cores_43_io_prev_bits_data),
    .io_prev_bits_wen(cores_43_io_prev_bits_wen),
    .io_prev_bits_id(cores_43_io_prev_bits_id),
    .io_next_ready(cores_43_io_next_ready),
    .io_next_valid(cores_43_io_next_valid),
    .io_next_bits_address(cores_43_io_next_bits_address),
    .io_next_bits_data(cores_43_io_next_bits_data),
    .io_next_bits_wen(cores_43_io_next_bits_wen),
    .io_next_bits_id(cores_43_io_next_bits_id)
  );
  RingCore_44 cores_44 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_44_clock),
    .reset(cores_44_reset),
    .io_prev_ready(cores_44_io_prev_ready),
    .io_prev_valid(cores_44_io_prev_valid),
    .io_prev_bits_address(cores_44_io_prev_bits_address),
    .io_prev_bits_data(cores_44_io_prev_bits_data),
    .io_prev_bits_wen(cores_44_io_prev_bits_wen),
    .io_prev_bits_id(cores_44_io_prev_bits_id),
    .io_next_ready(cores_44_io_next_ready),
    .io_next_valid(cores_44_io_next_valid),
    .io_next_bits_address(cores_44_io_next_bits_address),
    .io_next_bits_data(cores_44_io_next_bits_data),
    .io_next_bits_wen(cores_44_io_next_bits_wen),
    .io_next_bits_id(cores_44_io_next_bits_id)
  );
  RingCore_45 cores_45 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_45_clock),
    .reset(cores_45_reset),
    .io_prev_ready(cores_45_io_prev_ready),
    .io_prev_valid(cores_45_io_prev_valid),
    .io_prev_bits_address(cores_45_io_prev_bits_address),
    .io_prev_bits_data(cores_45_io_prev_bits_data),
    .io_prev_bits_wen(cores_45_io_prev_bits_wen),
    .io_prev_bits_id(cores_45_io_prev_bits_id),
    .io_next_ready(cores_45_io_next_ready),
    .io_next_valid(cores_45_io_next_valid),
    .io_next_bits_address(cores_45_io_next_bits_address),
    .io_next_bits_data(cores_45_io_next_bits_data),
    .io_next_bits_wen(cores_45_io_next_bits_wen),
    .io_next_bits_id(cores_45_io_next_bits_id)
  );
  RingCore_46 cores_46 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_46_clock),
    .reset(cores_46_reset),
    .io_prev_ready(cores_46_io_prev_ready),
    .io_prev_valid(cores_46_io_prev_valid),
    .io_prev_bits_address(cores_46_io_prev_bits_address),
    .io_prev_bits_data(cores_46_io_prev_bits_data),
    .io_prev_bits_wen(cores_46_io_prev_bits_wen),
    .io_prev_bits_id(cores_46_io_prev_bits_id),
    .io_next_ready(cores_46_io_next_ready),
    .io_next_valid(cores_46_io_next_valid),
    .io_next_bits_address(cores_46_io_next_bits_address),
    .io_next_bits_data(cores_46_io_next_bits_data),
    .io_next_bits_wen(cores_46_io_next_bits_wen),
    .io_next_bits_id(cores_46_io_next_bits_id)
  );
  RingCore_47 cores_47 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_47_clock),
    .reset(cores_47_reset),
    .io_prev_ready(cores_47_io_prev_ready),
    .io_prev_valid(cores_47_io_prev_valid),
    .io_prev_bits_address(cores_47_io_prev_bits_address),
    .io_prev_bits_data(cores_47_io_prev_bits_data),
    .io_prev_bits_wen(cores_47_io_prev_bits_wen),
    .io_prev_bits_id(cores_47_io_prev_bits_id),
    .io_next_ready(cores_47_io_next_ready),
    .io_next_valid(cores_47_io_next_valid),
    .io_next_bits_address(cores_47_io_next_bits_address),
    .io_next_bits_data(cores_47_io_next_bits_data),
    .io_next_bits_wen(cores_47_io_next_bits_wen),
    .io_next_bits_id(cores_47_io_next_bits_id)
  );
  RingCore_48 cores_48 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_48_clock),
    .reset(cores_48_reset),
    .io_prev_ready(cores_48_io_prev_ready),
    .io_prev_valid(cores_48_io_prev_valid),
    .io_prev_bits_address(cores_48_io_prev_bits_address),
    .io_prev_bits_data(cores_48_io_prev_bits_data),
    .io_prev_bits_wen(cores_48_io_prev_bits_wen),
    .io_prev_bits_id(cores_48_io_prev_bits_id),
    .io_next_ready(cores_48_io_next_ready),
    .io_next_valid(cores_48_io_next_valid),
    .io_next_bits_address(cores_48_io_next_bits_address),
    .io_next_bits_data(cores_48_io_next_bits_data),
    .io_next_bits_wen(cores_48_io_next_bits_wen),
    .io_next_bits_id(cores_48_io_next_bits_id)
  );
  RingCore_49 cores_49 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_49_clock),
    .reset(cores_49_reset),
    .io_prev_ready(cores_49_io_prev_ready),
    .io_prev_valid(cores_49_io_prev_valid),
    .io_prev_bits_address(cores_49_io_prev_bits_address),
    .io_prev_bits_data(cores_49_io_prev_bits_data),
    .io_prev_bits_wen(cores_49_io_prev_bits_wen),
    .io_prev_bits_id(cores_49_io_prev_bits_id),
    .io_next_ready(cores_49_io_next_ready),
    .io_next_valid(cores_49_io_next_valid),
    .io_next_bits_address(cores_49_io_next_bits_address),
    .io_next_bits_data(cores_49_io_next_bits_data),
    .io_next_bits_wen(cores_49_io_next_bits_wen),
    .io_next_bits_id(cores_49_io_next_bits_id)
  );
  RingCore_50 cores_50 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_50_clock),
    .reset(cores_50_reset),
    .io_prev_ready(cores_50_io_prev_ready),
    .io_prev_valid(cores_50_io_prev_valid),
    .io_prev_bits_address(cores_50_io_prev_bits_address),
    .io_prev_bits_data(cores_50_io_prev_bits_data),
    .io_prev_bits_wen(cores_50_io_prev_bits_wen),
    .io_prev_bits_id(cores_50_io_prev_bits_id),
    .io_next_ready(cores_50_io_next_ready),
    .io_next_valid(cores_50_io_next_valid),
    .io_next_bits_address(cores_50_io_next_bits_address),
    .io_next_bits_data(cores_50_io_next_bits_data),
    .io_next_bits_wen(cores_50_io_next_bits_wen),
    .io_next_bits_id(cores_50_io_next_bits_id)
  );
  RingCore_51 cores_51 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_51_clock),
    .reset(cores_51_reset),
    .io_prev_ready(cores_51_io_prev_ready),
    .io_prev_valid(cores_51_io_prev_valid),
    .io_prev_bits_address(cores_51_io_prev_bits_address),
    .io_prev_bits_data(cores_51_io_prev_bits_data),
    .io_prev_bits_wen(cores_51_io_prev_bits_wen),
    .io_prev_bits_id(cores_51_io_prev_bits_id),
    .io_next_ready(cores_51_io_next_ready),
    .io_next_valid(cores_51_io_next_valid),
    .io_next_bits_address(cores_51_io_next_bits_address),
    .io_next_bits_data(cores_51_io_next_bits_data),
    .io_next_bits_wen(cores_51_io_next_bits_wen),
    .io_next_bits_id(cores_51_io_next_bits_id)
  );
  RingCore_52 cores_52 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_52_clock),
    .reset(cores_52_reset),
    .io_prev_ready(cores_52_io_prev_ready),
    .io_prev_valid(cores_52_io_prev_valid),
    .io_prev_bits_address(cores_52_io_prev_bits_address),
    .io_prev_bits_data(cores_52_io_prev_bits_data),
    .io_prev_bits_wen(cores_52_io_prev_bits_wen),
    .io_prev_bits_id(cores_52_io_prev_bits_id),
    .io_next_ready(cores_52_io_next_ready),
    .io_next_valid(cores_52_io_next_valid),
    .io_next_bits_address(cores_52_io_next_bits_address),
    .io_next_bits_data(cores_52_io_next_bits_data),
    .io_next_bits_wen(cores_52_io_next_bits_wen),
    .io_next_bits_id(cores_52_io_next_bits_id)
  );
  RingCore_53 cores_53 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_53_clock),
    .reset(cores_53_reset),
    .io_prev_ready(cores_53_io_prev_ready),
    .io_prev_valid(cores_53_io_prev_valid),
    .io_prev_bits_address(cores_53_io_prev_bits_address),
    .io_prev_bits_data(cores_53_io_prev_bits_data),
    .io_prev_bits_wen(cores_53_io_prev_bits_wen),
    .io_prev_bits_id(cores_53_io_prev_bits_id),
    .io_next_ready(cores_53_io_next_ready),
    .io_next_valid(cores_53_io_next_valid),
    .io_next_bits_address(cores_53_io_next_bits_address),
    .io_next_bits_data(cores_53_io_next_bits_data),
    .io_next_bits_wen(cores_53_io_next_bits_wen),
    .io_next_bits_id(cores_53_io_next_bits_id)
  );
  RingCore_54 cores_54 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_54_clock),
    .reset(cores_54_reset),
    .io_prev_ready(cores_54_io_prev_ready),
    .io_prev_valid(cores_54_io_prev_valid),
    .io_prev_bits_address(cores_54_io_prev_bits_address),
    .io_prev_bits_data(cores_54_io_prev_bits_data),
    .io_prev_bits_wen(cores_54_io_prev_bits_wen),
    .io_prev_bits_id(cores_54_io_prev_bits_id),
    .io_next_ready(cores_54_io_next_ready),
    .io_next_valid(cores_54_io_next_valid),
    .io_next_bits_address(cores_54_io_next_bits_address),
    .io_next_bits_data(cores_54_io_next_bits_data),
    .io_next_bits_wen(cores_54_io_next_bits_wen),
    .io_next_bits_id(cores_54_io_next_bits_id)
  );
  RingCore_55 cores_55 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_55_clock),
    .reset(cores_55_reset),
    .io_prev_ready(cores_55_io_prev_ready),
    .io_prev_valid(cores_55_io_prev_valid),
    .io_prev_bits_address(cores_55_io_prev_bits_address),
    .io_prev_bits_data(cores_55_io_prev_bits_data),
    .io_prev_bits_wen(cores_55_io_prev_bits_wen),
    .io_prev_bits_id(cores_55_io_prev_bits_id),
    .io_next_ready(cores_55_io_next_ready),
    .io_next_valid(cores_55_io_next_valid),
    .io_next_bits_address(cores_55_io_next_bits_address),
    .io_next_bits_data(cores_55_io_next_bits_data),
    .io_next_bits_wen(cores_55_io_next_bits_wen),
    .io_next_bits_id(cores_55_io_next_bits_id)
  );
  RingCore_56 cores_56 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_56_clock),
    .reset(cores_56_reset),
    .io_prev_ready(cores_56_io_prev_ready),
    .io_prev_valid(cores_56_io_prev_valid),
    .io_prev_bits_address(cores_56_io_prev_bits_address),
    .io_prev_bits_data(cores_56_io_prev_bits_data),
    .io_prev_bits_wen(cores_56_io_prev_bits_wen),
    .io_prev_bits_id(cores_56_io_prev_bits_id),
    .io_next_ready(cores_56_io_next_ready),
    .io_next_valid(cores_56_io_next_valid),
    .io_next_bits_address(cores_56_io_next_bits_address),
    .io_next_bits_data(cores_56_io_next_bits_data),
    .io_next_bits_wen(cores_56_io_next_bits_wen),
    .io_next_bits_id(cores_56_io_next_bits_id)
  );
  RingCore_57 cores_57 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_57_clock),
    .reset(cores_57_reset),
    .io_prev_ready(cores_57_io_prev_ready),
    .io_prev_valid(cores_57_io_prev_valid),
    .io_prev_bits_address(cores_57_io_prev_bits_address),
    .io_prev_bits_data(cores_57_io_prev_bits_data),
    .io_prev_bits_wen(cores_57_io_prev_bits_wen),
    .io_prev_bits_id(cores_57_io_prev_bits_id),
    .io_next_ready(cores_57_io_next_ready),
    .io_next_valid(cores_57_io_next_valid),
    .io_next_bits_address(cores_57_io_next_bits_address),
    .io_next_bits_data(cores_57_io_next_bits_data),
    .io_next_bits_wen(cores_57_io_next_bits_wen),
    .io_next_bits_id(cores_57_io_next_bits_id)
  );
  RingCore_58 cores_58 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_58_clock),
    .reset(cores_58_reset),
    .io_prev_ready(cores_58_io_prev_ready),
    .io_prev_valid(cores_58_io_prev_valid),
    .io_prev_bits_address(cores_58_io_prev_bits_address),
    .io_prev_bits_data(cores_58_io_prev_bits_data),
    .io_prev_bits_wen(cores_58_io_prev_bits_wen),
    .io_prev_bits_id(cores_58_io_prev_bits_id),
    .io_next_ready(cores_58_io_next_ready),
    .io_next_valid(cores_58_io_next_valid),
    .io_next_bits_address(cores_58_io_next_bits_address),
    .io_next_bits_data(cores_58_io_next_bits_data),
    .io_next_bits_wen(cores_58_io_next_bits_wen),
    .io_next_bits_id(cores_58_io_next_bits_id)
  );
  RingCore_59 cores_59 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_59_clock),
    .reset(cores_59_reset),
    .io_prev_ready(cores_59_io_prev_ready),
    .io_prev_valid(cores_59_io_prev_valid),
    .io_prev_bits_address(cores_59_io_prev_bits_address),
    .io_prev_bits_data(cores_59_io_prev_bits_data),
    .io_prev_bits_wen(cores_59_io_prev_bits_wen),
    .io_prev_bits_id(cores_59_io_prev_bits_id),
    .io_next_ready(cores_59_io_next_ready),
    .io_next_valid(cores_59_io_next_valid),
    .io_next_bits_address(cores_59_io_next_bits_address),
    .io_next_bits_data(cores_59_io_next_bits_data),
    .io_next_bits_wen(cores_59_io_next_bits_wen),
    .io_next_bits_id(cores_59_io_next_bits_id)
  );
  RingCore_60 cores_60 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_60_clock),
    .reset(cores_60_reset),
    .io_prev_ready(cores_60_io_prev_ready),
    .io_prev_valid(cores_60_io_prev_valid),
    .io_prev_bits_address(cores_60_io_prev_bits_address),
    .io_prev_bits_data(cores_60_io_prev_bits_data),
    .io_prev_bits_wen(cores_60_io_prev_bits_wen),
    .io_prev_bits_id(cores_60_io_prev_bits_id),
    .io_next_ready(cores_60_io_next_ready),
    .io_next_valid(cores_60_io_next_valid),
    .io_next_bits_address(cores_60_io_next_bits_address),
    .io_next_bits_data(cores_60_io_next_bits_data),
    .io_next_bits_wen(cores_60_io_next_bits_wen),
    .io_next_bits_id(cores_60_io_next_bits_id)
  );
  RingCore_61 cores_61 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_61_clock),
    .reset(cores_61_reset),
    .io_prev_ready(cores_61_io_prev_ready),
    .io_prev_valid(cores_61_io_prev_valid),
    .io_prev_bits_address(cores_61_io_prev_bits_address),
    .io_prev_bits_data(cores_61_io_prev_bits_data),
    .io_prev_bits_wen(cores_61_io_prev_bits_wen),
    .io_prev_bits_id(cores_61_io_prev_bits_id),
    .io_next_ready(cores_61_io_next_ready),
    .io_next_valid(cores_61_io_next_valid),
    .io_next_bits_address(cores_61_io_next_bits_address),
    .io_next_bits_data(cores_61_io_next_bits_data),
    .io_next_bits_wen(cores_61_io_next_bits_wen),
    .io_next_bits_id(cores_61_io_next_bits_id)
  );
  RingCore_62 cores_62 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_62_clock),
    .reset(cores_62_reset),
    .io_prev_ready(cores_62_io_prev_ready),
    .io_prev_valid(cores_62_io_prev_valid),
    .io_prev_bits_address(cores_62_io_prev_bits_address),
    .io_prev_bits_data(cores_62_io_prev_bits_data),
    .io_prev_bits_wen(cores_62_io_prev_bits_wen),
    .io_prev_bits_id(cores_62_io_prev_bits_id),
    .io_next_ready(cores_62_io_next_ready),
    .io_next_valid(cores_62_io_next_valid),
    .io_next_bits_address(cores_62_io_next_bits_address),
    .io_next_bits_data(cores_62_io_next_bits_data),
    .io_next_bits_wen(cores_62_io_next_bits_wen),
    .io_next_bits_id(cores_62_io_next_bits_id)
  );
  RingCore_63 cores_63 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_63_clock),
    .reset(cores_63_reset),
    .io_prev_ready(cores_63_io_prev_ready),
    .io_prev_valid(cores_63_io_prev_valid),
    .io_prev_bits_address(cores_63_io_prev_bits_address),
    .io_prev_bits_data(cores_63_io_prev_bits_data),
    .io_prev_bits_wen(cores_63_io_prev_bits_wen),
    .io_prev_bits_id(cores_63_io_prev_bits_id),
    .io_next_ready(cores_63_io_next_ready),
    .io_next_valid(cores_63_io_next_valid),
    .io_next_bits_address(cores_63_io_next_bits_address),
    .io_next_bits_data(cores_63_io_next_bits_data),
    .io_next_bits_wen(cores_63_io_next_bits_wen),
    .io_next_bits_id(cores_63_io_next_bits_id)
  );
  RingCore_64 cores_64 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_64_clock),
    .reset(cores_64_reset),
    .io_prev_ready(cores_64_io_prev_ready),
    .io_prev_valid(cores_64_io_prev_valid),
    .io_prev_bits_address(cores_64_io_prev_bits_address),
    .io_prev_bits_data(cores_64_io_prev_bits_data),
    .io_prev_bits_wen(cores_64_io_prev_bits_wen),
    .io_prev_bits_id(cores_64_io_prev_bits_id),
    .io_next_ready(cores_64_io_next_ready),
    .io_next_valid(cores_64_io_next_valid),
    .io_next_bits_address(cores_64_io_next_bits_address),
    .io_next_bits_data(cores_64_io_next_bits_data),
    .io_next_bits_wen(cores_64_io_next_bits_wen),
    .io_next_bits_id(cores_64_io_next_bits_id)
  );
  RingCore_65 cores_65 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_65_clock),
    .reset(cores_65_reset),
    .io_prev_ready(cores_65_io_prev_ready),
    .io_prev_valid(cores_65_io_prev_valid),
    .io_prev_bits_address(cores_65_io_prev_bits_address),
    .io_prev_bits_data(cores_65_io_prev_bits_data),
    .io_prev_bits_wen(cores_65_io_prev_bits_wen),
    .io_prev_bits_id(cores_65_io_prev_bits_id),
    .io_next_ready(cores_65_io_next_ready),
    .io_next_valid(cores_65_io_next_valid),
    .io_next_bits_address(cores_65_io_next_bits_address),
    .io_next_bits_data(cores_65_io_next_bits_data),
    .io_next_bits_wen(cores_65_io_next_bits_wen),
    .io_next_bits_id(cores_65_io_next_bits_id)
  );
  RingCore_66 cores_66 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_66_clock),
    .reset(cores_66_reset),
    .io_prev_ready(cores_66_io_prev_ready),
    .io_prev_valid(cores_66_io_prev_valid),
    .io_prev_bits_address(cores_66_io_prev_bits_address),
    .io_prev_bits_data(cores_66_io_prev_bits_data),
    .io_prev_bits_wen(cores_66_io_prev_bits_wen),
    .io_prev_bits_id(cores_66_io_prev_bits_id),
    .io_next_ready(cores_66_io_next_ready),
    .io_next_valid(cores_66_io_next_valid),
    .io_next_bits_address(cores_66_io_next_bits_address),
    .io_next_bits_data(cores_66_io_next_bits_data),
    .io_next_bits_wen(cores_66_io_next_bits_wen),
    .io_next_bits_id(cores_66_io_next_bits_id)
  );
  RingCore_67 cores_67 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_67_clock),
    .reset(cores_67_reset),
    .io_prev_ready(cores_67_io_prev_ready),
    .io_prev_valid(cores_67_io_prev_valid),
    .io_prev_bits_address(cores_67_io_prev_bits_address),
    .io_prev_bits_data(cores_67_io_prev_bits_data),
    .io_prev_bits_wen(cores_67_io_prev_bits_wen),
    .io_prev_bits_id(cores_67_io_prev_bits_id),
    .io_next_ready(cores_67_io_next_ready),
    .io_next_valid(cores_67_io_next_valid),
    .io_next_bits_address(cores_67_io_next_bits_address),
    .io_next_bits_data(cores_67_io_next_bits_data),
    .io_next_bits_wen(cores_67_io_next_bits_wen),
    .io_next_bits_id(cores_67_io_next_bits_id)
  );
  RingCore_68 cores_68 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_68_clock),
    .reset(cores_68_reset),
    .io_prev_ready(cores_68_io_prev_ready),
    .io_prev_valid(cores_68_io_prev_valid),
    .io_prev_bits_address(cores_68_io_prev_bits_address),
    .io_prev_bits_data(cores_68_io_prev_bits_data),
    .io_prev_bits_wen(cores_68_io_prev_bits_wen),
    .io_prev_bits_id(cores_68_io_prev_bits_id),
    .io_next_ready(cores_68_io_next_ready),
    .io_next_valid(cores_68_io_next_valid),
    .io_next_bits_address(cores_68_io_next_bits_address),
    .io_next_bits_data(cores_68_io_next_bits_data),
    .io_next_bits_wen(cores_68_io_next_bits_wen),
    .io_next_bits_id(cores_68_io_next_bits_id)
  );
  RingCore_69 cores_69 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_69_clock),
    .reset(cores_69_reset),
    .io_prev_ready(cores_69_io_prev_ready),
    .io_prev_valid(cores_69_io_prev_valid),
    .io_prev_bits_address(cores_69_io_prev_bits_address),
    .io_prev_bits_data(cores_69_io_prev_bits_data),
    .io_prev_bits_wen(cores_69_io_prev_bits_wen),
    .io_prev_bits_id(cores_69_io_prev_bits_id),
    .io_next_ready(cores_69_io_next_ready),
    .io_next_valid(cores_69_io_next_valid),
    .io_next_bits_address(cores_69_io_next_bits_address),
    .io_next_bits_data(cores_69_io_next_bits_data),
    .io_next_bits_wen(cores_69_io_next_bits_wen),
    .io_next_bits_id(cores_69_io_next_bits_id)
  );
  RingCore_70 cores_70 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_70_clock),
    .reset(cores_70_reset),
    .io_prev_ready(cores_70_io_prev_ready),
    .io_prev_valid(cores_70_io_prev_valid),
    .io_prev_bits_address(cores_70_io_prev_bits_address),
    .io_prev_bits_data(cores_70_io_prev_bits_data),
    .io_prev_bits_wen(cores_70_io_prev_bits_wen),
    .io_prev_bits_id(cores_70_io_prev_bits_id),
    .io_next_ready(cores_70_io_next_ready),
    .io_next_valid(cores_70_io_next_valid),
    .io_next_bits_address(cores_70_io_next_bits_address),
    .io_next_bits_data(cores_70_io_next_bits_data),
    .io_next_bits_wen(cores_70_io_next_bits_wen),
    .io_next_bits_id(cores_70_io_next_bits_id)
  );
  RingCore_71 cores_71 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_71_clock),
    .reset(cores_71_reset),
    .io_prev_ready(cores_71_io_prev_ready),
    .io_prev_valid(cores_71_io_prev_valid),
    .io_prev_bits_address(cores_71_io_prev_bits_address),
    .io_prev_bits_data(cores_71_io_prev_bits_data),
    .io_prev_bits_wen(cores_71_io_prev_bits_wen),
    .io_prev_bits_id(cores_71_io_prev_bits_id),
    .io_next_ready(cores_71_io_next_ready),
    .io_next_valid(cores_71_io_next_valid),
    .io_next_bits_address(cores_71_io_next_bits_address),
    .io_next_bits_data(cores_71_io_next_bits_data),
    .io_next_bits_wen(cores_71_io_next_bits_wen),
    .io_next_bits_id(cores_71_io_next_bits_id)
  );
  RingCore_72 cores_72 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_72_clock),
    .reset(cores_72_reset),
    .io_prev_ready(cores_72_io_prev_ready),
    .io_prev_valid(cores_72_io_prev_valid),
    .io_prev_bits_address(cores_72_io_prev_bits_address),
    .io_prev_bits_data(cores_72_io_prev_bits_data),
    .io_prev_bits_wen(cores_72_io_prev_bits_wen),
    .io_prev_bits_id(cores_72_io_prev_bits_id),
    .io_next_ready(cores_72_io_next_ready),
    .io_next_valid(cores_72_io_next_valid),
    .io_next_bits_address(cores_72_io_next_bits_address),
    .io_next_bits_data(cores_72_io_next_bits_data),
    .io_next_bits_wen(cores_72_io_next_bits_wen),
    .io_next_bits_id(cores_72_io_next_bits_id)
  );
  RingCore_73 cores_73 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_73_clock),
    .reset(cores_73_reset),
    .io_prev_ready(cores_73_io_prev_ready),
    .io_prev_valid(cores_73_io_prev_valid),
    .io_prev_bits_address(cores_73_io_prev_bits_address),
    .io_prev_bits_data(cores_73_io_prev_bits_data),
    .io_prev_bits_wen(cores_73_io_prev_bits_wen),
    .io_prev_bits_id(cores_73_io_prev_bits_id),
    .io_next_ready(cores_73_io_next_ready),
    .io_next_valid(cores_73_io_next_valid),
    .io_next_bits_address(cores_73_io_next_bits_address),
    .io_next_bits_data(cores_73_io_next_bits_data),
    .io_next_bits_wen(cores_73_io_next_bits_wen),
    .io_next_bits_id(cores_73_io_next_bits_id)
  );
  RingCore_74 cores_74 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_74_clock),
    .reset(cores_74_reset),
    .io_prev_ready(cores_74_io_prev_ready),
    .io_prev_valid(cores_74_io_prev_valid),
    .io_prev_bits_address(cores_74_io_prev_bits_address),
    .io_prev_bits_data(cores_74_io_prev_bits_data),
    .io_prev_bits_wen(cores_74_io_prev_bits_wen),
    .io_prev_bits_id(cores_74_io_prev_bits_id),
    .io_next_ready(cores_74_io_next_ready),
    .io_next_valid(cores_74_io_next_valid),
    .io_next_bits_address(cores_74_io_next_bits_address),
    .io_next_bits_data(cores_74_io_next_bits_data),
    .io_next_bits_wen(cores_74_io_next_bits_wen),
    .io_next_bits_id(cores_74_io_next_bits_id)
  );
  RingCore_75 cores_75 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_75_clock),
    .reset(cores_75_reset),
    .io_prev_ready(cores_75_io_prev_ready),
    .io_prev_valid(cores_75_io_prev_valid),
    .io_prev_bits_address(cores_75_io_prev_bits_address),
    .io_prev_bits_data(cores_75_io_prev_bits_data),
    .io_prev_bits_wen(cores_75_io_prev_bits_wen),
    .io_prev_bits_id(cores_75_io_prev_bits_id),
    .io_next_ready(cores_75_io_next_ready),
    .io_next_valid(cores_75_io_next_valid),
    .io_next_bits_address(cores_75_io_next_bits_address),
    .io_next_bits_data(cores_75_io_next_bits_data),
    .io_next_bits_wen(cores_75_io_next_bits_wen),
    .io_next_bits_id(cores_75_io_next_bits_id)
  );
  RingCore_76 cores_76 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_76_clock),
    .reset(cores_76_reset),
    .io_prev_ready(cores_76_io_prev_ready),
    .io_prev_valid(cores_76_io_prev_valid),
    .io_prev_bits_address(cores_76_io_prev_bits_address),
    .io_prev_bits_data(cores_76_io_prev_bits_data),
    .io_prev_bits_wen(cores_76_io_prev_bits_wen),
    .io_prev_bits_id(cores_76_io_prev_bits_id),
    .io_next_ready(cores_76_io_next_ready),
    .io_next_valid(cores_76_io_next_valid),
    .io_next_bits_address(cores_76_io_next_bits_address),
    .io_next_bits_data(cores_76_io_next_bits_data),
    .io_next_bits_wen(cores_76_io_next_bits_wen),
    .io_next_bits_id(cores_76_io_next_bits_id)
  );
  RingCore_77 cores_77 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_77_clock),
    .reset(cores_77_reset),
    .io_prev_ready(cores_77_io_prev_ready),
    .io_prev_valid(cores_77_io_prev_valid),
    .io_prev_bits_address(cores_77_io_prev_bits_address),
    .io_prev_bits_data(cores_77_io_prev_bits_data),
    .io_prev_bits_wen(cores_77_io_prev_bits_wen),
    .io_prev_bits_id(cores_77_io_prev_bits_id),
    .io_next_ready(cores_77_io_next_ready),
    .io_next_valid(cores_77_io_next_valid),
    .io_next_bits_address(cores_77_io_next_bits_address),
    .io_next_bits_data(cores_77_io_next_bits_data),
    .io_next_bits_wen(cores_77_io_next_bits_wen),
    .io_next_bits_id(cores_77_io_next_bits_id)
  );
  RingCore_78 cores_78 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_78_clock),
    .reset(cores_78_reset),
    .io_prev_ready(cores_78_io_prev_ready),
    .io_prev_valid(cores_78_io_prev_valid),
    .io_prev_bits_address(cores_78_io_prev_bits_address),
    .io_prev_bits_data(cores_78_io_prev_bits_data),
    .io_prev_bits_wen(cores_78_io_prev_bits_wen),
    .io_prev_bits_id(cores_78_io_prev_bits_id),
    .io_next_ready(cores_78_io_next_ready),
    .io_next_valid(cores_78_io_next_valid),
    .io_next_bits_address(cores_78_io_next_bits_address),
    .io_next_bits_data(cores_78_io_next_bits_data),
    .io_next_bits_wen(cores_78_io_next_bits_wen),
    .io_next_bits_id(cores_78_io_next_bits_id)
  );
  RingCore_79 cores_79 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_79_clock),
    .reset(cores_79_reset),
    .io_prev_ready(cores_79_io_prev_ready),
    .io_prev_valid(cores_79_io_prev_valid),
    .io_prev_bits_address(cores_79_io_prev_bits_address),
    .io_prev_bits_data(cores_79_io_prev_bits_data),
    .io_prev_bits_wen(cores_79_io_prev_bits_wen),
    .io_prev_bits_id(cores_79_io_prev_bits_id),
    .io_next_ready(cores_79_io_next_ready),
    .io_next_valid(cores_79_io_next_valid),
    .io_next_bits_address(cores_79_io_next_bits_address),
    .io_next_bits_data(cores_79_io_next_bits_data),
    .io_next_bits_wen(cores_79_io_next_bits_wen),
    .io_next_bits_id(cores_79_io_next_bits_id)
  );
  RingCore_80 cores_80 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_80_clock),
    .reset(cores_80_reset),
    .io_prev_ready(cores_80_io_prev_ready),
    .io_prev_valid(cores_80_io_prev_valid),
    .io_prev_bits_address(cores_80_io_prev_bits_address),
    .io_prev_bits_data(cores_80_io_prev_bits_data),
    .io_prev_bits_wen(cores_80_io_prev_bits_wen),
    .io_prev_bits_id(cores_80_io_prev_bits_id),
    .io_next_ready(cores_80_io_next_ready),
    .io_next_valid(cores_80_io_next_valid),
    .io_next_bits_address(cores_80_io_next_bits_address),
    .io_next_bits_data(cores_80_io_next_bits_data),
    .io_next_bits_wen(cores_80_io_next_bits_wen),
    .io_next_bits_id(cores_80_io_next_bits_id)
  );
  RingCore_81 cores_81 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_81_clock),
    .reset(cores_81_reset),
    .io_prev_ready(cores_81_io_prev_ready),
    .io_prev_valid(cores_81_io_prev_valid),
    .io_prev_bits_address(cores_81_io_prev_bits_address),
    .io_prev_bits_data(cores_81_io_prev_bits_data),
    .io_prev_bits_wen(cores_81_io_prev_bits_wen),
    .io_prev_bits_id(cores_81_io_prev_bits_id),
    .io_next_ready(cores_81_io_next_ready),
    .io_next_valid(cores_81_io_next_valid),
    .io_next_bits_address(cores_81_io_next_bits_address),
    .io_next_bits_data(cores_81_io_next_bits_data),
    .io_next_bits_wen(cores_81_io_next_bits_wen),
    .io_next_bits_id(cores_81_io_next_bits_id)
  );
  RingCore_82 cores_82 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_82_clock),
    .reset(cores_82_reset),
    .io_prev_ready(cores_82_io_prev_ready),
    .io_prev_valid(cores_82_io_prev_valid),
    .io_prev_bits_address(cores_82_io_prev_bits_address),
    .io_prev_bits_data(cores_82_io_prev_bits_data),
    .io_prev_bits_wen(cores_82_io_prev_bits_wen),
    .io_prev_bits_id(cores_82_io_prev_bits_id),
    .io_next_ready(cores_82_io_next_ready),
    .io_next_valid(cores_82_io_next_valid),
    .io_next_bits_address(cores_82_io_next_bits_address),
    .io_next_bits_data(cores_82_io_next_bits_data),
    .io_next_bits_wen(cores_82_io_next_bits_wen),
    .io_next_bits_id(cores_82_io_next_bits_id)
  );
  RingCore_83 cores_83 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_83_clock),
    .reset(cores_83_reset),
    .io_prev_ready(cores_83_io_prev_ready),
    .io_prev_valid(cores_83_io_prev_valid),
    .io_prev_bits_address(cores_83_io_prev_bits_address),
    .io_prev_bits_data(cores_83_io_prev_bits_data),
    .io_prev_bits_wen(cores_83_io_prev_bits_wen),
    .io_prev_bits_id(cores_83_io_prev_bits_id),
    .io_next_ready(cores_83_io_next_ready),
    .io_next_valid(cores_83_io_next_valid),
    .io_next_bits_address(cores_83_io_next_bits_address),
    .io_next_bits_data(cores_83_io_next_bits_data),
    .io_next_bits_wen(cores_83_io_next_bits_wen),
    .io_next_bits_id(cores_83_io_next_bits_id)
  );
  RingCore_84 cores_84 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_84_clock),
    .reset(cores_84_reset),
    .io_prev_ready(cores_84_io_prev_ready),
    .io_prev_valid(cores_84_io_prev_valid),
    .io_prev_bits_address(cores_84_io_prev_bits_address),
    .io_prev_bits_data(cores_84_io_prev_bits_data),
    .io_prev_bits_wen(cores_84_io_prev_bits_wen),
    .io_prev_bits_id(cores_84_io_prev_bits_id),
    .io_next_ready(cores_84_io_next_ready),
    .io_next_valid(cores_84_io_next_valid),
    .io_next_bits_address(cores_84_io_next_bits_address),
    .io_next_bits_data(cores_84_io_next_bits_data),
    .io_next_bits_wen(cores_84_io_next_bits_wen),
    .io_next_bits_id(cores_84_io_next_bits_id)
  );
  RingCore_85 cores_85 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_85_clock),
    .reset(cores_85_reset),
    .io_prev_ready(cores_85_io_prev_ready),
    .io_prev_valid(cores_85_io_prev_valid),
    .io_prev_bits_address(cores_85_io_prev_bits_address),
    .io_prev_bits_data(cores_85_io_prev_bits_data),
    .io_prev_bits_wen(cores_85_io_prev_bits_wen),
    .io_prev_bits_id(cores_85_io_prev_bits_id),
    .io_next_ready(cores_85_io_next_ready),
    .io_next_valid(cores_85_io_next_valid),
    .io_next_bits_address(cores_85_io_next_bits_address),
    .io_next_bits_data(cores_85_io_next_bits_data),
    .io_next_bits_wen(cores_85_io_next_bits_wen),
    .io_next_bits_id(cores_85_io_next_bits_id)
  );
  RingCore_86 cores_86 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_86_clock),
    .reset(cores_86_reset),
    .io_prev_ready(cores_86_io_prev_ready),
    .io_prev_valid(cores_86_io_prev_valid),
    .io_prev_bits_address(cores_86_io_prev_bits_address),
    .io_prev_bits_data(cores_86_io_prev_bits_data),
    .io_prev_bits_wen(cores_86_io_prev_bits_wen),
    .io_prev_bits_id(cores_86_io_prev_bits_id),
    .io_next_ready(cores_86_io_next_ready),
    .io_next_valid(cores_86_io_next_valid),
    .io_next_bits_address(cores_86_io_next_bits_address),
    .io_next_bits_data(cores_86_io_next_bits_data),
    .io_next_bits_wen(cores_86_io_next_bits_wen),
    .io_next_bits_id(cores_86_io_next_bits_id)
  );
  RingCore_87 cores_87 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_87_clock),
    .reset(cores_87_reset),
    .io_prev_ready(cores_87_io_prev_ready),
    .io_prev_valid(cores_87_io_prev_valid),
    .io_prev_bits_address(cores_87_io_prev_bits_address),
    .io_prev_bits_data(cores_87_io_prev_bits_data),
    .io_prev_bits_wen(cores_87_io_prev_bits_wen),
    .io_prev_bits_id(cores_87_io_prev_bits_id),
    .io_next_ready(cores_87_io_next_ready),
    .io_next_valid(cores_87_io_next_valid),
    .io_next_bits_address(cores_87_io_next_bits_address),
    .io_next_bits_data(cores_87_io_next_bits_data),
    .io_next_bits_wen(cores_87_io_next_bits_wen),
    .io_next_bits_id(cores_87_io_next_bits_id)
  );
  RingCore_88 cores_88 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_88_clock),
    .reset(cores_88_reset),
    .io_prev_ready(cores_88_io_prev_ready),
    .io_prev_valid(cores_88_io_prev_valid),
    .io_prev_bits_address(cores_88_io_prev_bits_address),
    .io_prev_bits_data(cores_88_io_prev_bits_data),
    .io_prev_bits_wen(cores_88_io_prev_bits_wen),
    .io_prev_bits_id(cores_88_io_prev_bits_id),
    .io_next_ready(cores_88_io_next_ready),
    .io_next_valid(cores_88_io_next_valid),
    .io_next_bits_address(cores_88_io_next_bits_address),
    .io_next_bits_data(cores_88_io_next_bits_data),
    .io_next_bits_wen(cores_88_io_next_bits_wen),
    .io_next_bits_id(cores_88_io_next_bits_id)
  );
  RingCore_89 cores_89 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_89_clock),
    .reset(cores_89_reset),
    .io_prev_ready(cores_89_io_prev_ready),
    .io_prev_valid(cores_89_io_prev_valid),
    .io_prev_bits_address(cores_89_io_prev_bits_address),
    .io_prev_bits_data(cores_89_io_prev_bits_data),
    .io_prev_bits_wen(cores_89_io_prev_bits_wen),
    .io_prev_bits_id(cores_89_io_prev_bits_id),
    .io_next_ready(cores_89_io_next_ready),
    .io_next_valid(cores_89_io_next_valid),
    .io_next_bits_address(cores_89_io_next_bits_address),
    .io_next_bits_data(cores_89_io_next_bits_data),
    .io_next_bits_wen(cores_89_io_next_bits_wen),
    .io_next_bits_id(cores_89_io_next_bits_id)
  );
  RingCore_90 cores_90 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_90_clock),
    .reset(cores_90_reset),
    .io_prev_ready(cores_90_io_prev_ready),
    .io_prev_valid(cores_90_io_prev_valid),
    .io_prev_bits_address(cores_90_io_prev_bits_address),
    .io_prev_bits_data(cores_90_io_prev_bits_data),
    .io_prev_bits_wen(cores_90_io_prev_bits_wen),
    .io_prev_bits_id(cores_90_io_prev_bits_id),
    .io_next_ready(cores_90_io_next_ready),
    .io_next_valid(cores_90_io_next_valid),
    .io_next_bits_address(cores_90_io_next_bits_address),
    .io_next_bits_data(cores_90_io_next_bits_data),
    .io_next_bits_wen(cores_90_io_next_bits_wen),
    .io_next_bits_id(cores_90_io_next_bits_id)
  );
  RingCore_91 cores_91 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_91_clock),
    .reset(cores_91_reset),
    .io_prev_ready(cores_91_io_prev_ready),
    .io_prev_valid(cores_91_io_prev_valid),
    .io_prev_bits_address(cores_91_io_prev_bits_address),
    .io_prev_bits_data(cores_91_io_prev_bits_data),
    .io_prev_bits_wen(cores_91_io_prev_bits_wen),
    .io_prev_bits_id(cores_91_io_prev_bits_id),
    .io_next_ready(cores_91_io_next_ready),
    .io_next_valid(cores_91_io_next_valid),
    .io_next_bits_address(cores_91_io_next_bits_address),
    .io_next_bits_data(cores_91_io_next_bits_data),
    .io_next_bits_wen(cores_91_io_next_bits_wen),
    .io_next_bits_id(cores_91_io_next_bits_id)
  );
  RingCore_92 cores_92 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_92_clock),
    .reset(cores_92_reset),
    .io_prev_ready(cores_92_io_prev_ready),
    .io_prev_valid(cores_92_io_prev_valid),
    .io_prev_bits_address(cores_92_io_prev_bits_address),
    .io_prev_bits_data(cores_92_io_prev_bits_data),
    .io_prev_bits_wen(cores_92_io_prev_bits_wen),
    .io_prev_bits_id(cores_92_io_prev_bits_id),
    .io_next_ready(cores_92_io_next_ready),
    .io_next_valid(cores_92_io_next_valid),
    .io_next_bits_address(cores_92_io_next_bits_address),
    .io_next_bits_data(cores_92_io_next_bits_data),
    .io_next_bits_wen(cores_92_io_next_bits_wen),
    .io_next_bits_id(cores_92_io_next_bits_id)
  );
  RingCore_93 cores_93 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_93_clock),
    .reset(cores_93_reset),
    .io_prev_ready(cores_93_io_prev_ready),
    .io_prev_valid(cores_93_io_prev_valid),
    .io_prev_bits_address(cores_93_io_prev_bits_address),
    .io_prev_bits_data(cores_93_io_prev_bits_data),
    .io_prev_bits_wen(cores_93_io_prev_bits_wen),
    .io_prev_bits_id(cores_93_io_prev_bits_id),
    .io_next_ready(cores_93_io_next_ready),
    .io_next_valid(cores_93_io_next_valid),
    .io_next_bits_address(cores_93_io_next_bits_address),
    .io_next_bits_data(cores_93_io_next_bits_data),
    .io_next_bits_wen(cores_93_io_next_bits_wen),
    .io_next_bits_id(cores_93_io_next_bits_id)
  );
  RingCore_94 cores_94 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_94_clock),
    .reset(cores_94_reset),
    .io_prev_ready(cores_94_io_prev_ready),
    .io_prev_valid(cores_94_io_prev_valid),
    .io_prev_bits_address(cores_94_io_prev_bits_address),
    .io_prev_bits_data(cores_94_io_prev_bits_data),
    .io_prev_bits_wen(cores_94_io_prev_bits_wen),
    .io_prev_bits_id(cores_94_io_prev_bits_id),
    .io_next_ready(cores_94_io_next_ready),
    .io_next_valid(cores_94_io_next_valid),
    .io_next_bits_address(cores_94_io_next_bits_address),
    .io_next_bits_data(cores_94_io_next_bits_data),
    .io_next_bits_wen(cores_94_io_next_bits_wen),
    .io_next_bits_id(cores_94_io_next_bits_id)
  );
  RingCore_95 cores_95 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_95_clock),
    .reset(cores_95_reset),
    .io_prev_ready(cores_95_io_prev_ready),
    .io_prev_valid(cores_95_io_prev_valid),
    .io_prev_bits_address(cores_95_io_prev_bits_address),
    .io_prev_bits_data(cores_95_io_prev_bits_data),
    .io_prev_bits_wen(cores_95_io_prev_bits_wen),
    .io_prev_bits_id(cores_95_io_prev_bits_id),
    .io_next_ready(cores_95_io_next_ready),
    .io_next_valid(cores_95_io_next_valid),
    .io_next_bits_address(cores_95_io_next_bits_address),
    .io_next_bits_data(cores_95_io_next_bits_data),
    .io_next_bits_wen(cores_95_io_next_bits_wen),
    .io_next_bits_id(cores_95_io_next_bits_id)
  );
  RingCore_96 cores_96 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_96_clock),
    .reset(cores_96_reset),
    .io_prev_ready(cores_96_io_prev_ready),
    .io_prev_valid(cores_96_io_prev_valid),
    .io_prev_bits_address(cores_96_io_prev_bits_address),
    .io_prev_bits_data(cores_96_io_prev_bits_data),
    .io_prev_bits_wen(cores_96_io_prev_bits_wen),
    .io_prev_bits_id(cores_96_io_prev_bits_id),
    .io_next_ready(cores_96_io_next_ready),
    .io_next_valid(cores_96_io_next_valid),
    .io_next_bits_address(cores_96_io_next_bits_address),
    .io_next_bits_data(cores_96_io_next_bits_data),
    .io_next_bits_wen(cores_96_io_next_bits_wen),
    .io_next_bits_id(cores_96_io_next_bits_id)
  );
  RingCore_97 cores_97 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_97_clock),
    .reset(cores_97_reset),
    .io_prev_ready(cores_97_io_prev_ready),
    .io_prev_valid(cores_97_io_prev_valid),
    .io_prev_bits_address(cores_97_io_prev_bits_address),
    .io_prev_bits_data(cores_97_io_prev_bits_data),
    .io_prev_bits_wen(cores_97_io_prev_bits_wen),
    .io_prev_bits_id(cores_97_io_prev_bits_id),
    .io_next_ready(cores_97_io_next_ready),
    .io_next_valid(cores_97_io_next_valid),
    .io_next_bits_address(cores_97_io_next_bits_address),
    .io_next_bits_data(cores_97_io_next_bits_data),
    .io_next_bits_wen(cores_97_io_next_bits_wen),
    .io_next_bits_id(cores_97_io_next_bits_id)
  );
  RingCore_98 cores_98 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_98_clock),
    .reset(cores_98_reset),
    .io_prev_ready(cores_98_io_prev_ready),
    .io_prev_valid(cores_98_io_prev_valid),
    .io_prev_bits_address(cores_98_io_prev_bits_address),
    .io_prev_bits_data(cores_98_io_prev_bits_data),
    .io_prev_bits_wen(cores_98_io_prev_bits_wen),
    .io_prev_bits_id(cores_98_io_prev_bits_id),
    .io_next_ready(cores_98_io_next_ready),
    .io_next_valid(cores_98_io_next_valid),
    .io_next_bits_address(cores_98_io_next_bits_address),
    .io_next_bits_data(cores_98_io_next_bits_data),
    .io_next_bits_wen(cores_98_io_next_bits_wen),
    .io_next_bits_id(cores_98_io_next_bits_id)
  );
  RingCore_99 cores_99 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_99_clock),
    .reset(cores_99_reset),
    .io_prev_ready(cores_99_io_prev_ready),
    .io_prev_valid(cores_99_io_prev_valid),
    .io_prev_bits_address(cores_99_io_prev_bits_address),
    .io_prev_bits_data(cores_99_io_prev_bits_data),
    .io_prev_bits_wen(cores_99_io_prev_bits_wen),
    .io_prev_bits_id(cores_99_io_prev_bits_id),
    .io_next_ready(cores_99_io_next_ready),
    .io_next_valid(cores_99_io_next_valid),
    .io_next_bits_address(cores_99_io_next_bits_address),
    .io_next_bits_data(cores_99_io_next_bits_data),
    .io_next_bits_wen(cores_99_io_next_bits_wen),
    .io_next_bits_id(cores_99_io_next_bits_id)
  );
  RingCore_100 cores_100 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_100_clock),
    .reset(cores_100_reset),
    .io_prev_ready(cores_100_io_prev_ready),
    .io_prev_valid(cores_100_io_prev_valid),
    .io_prev_bits_address(cores_100_io_prev_bits_address),
    .io_prev_bits_data(cores_100_io_prev_bits_data),
    .io_prev_bits_wen(cores_100_io_prev_bits_wen),
    .io_prev_bits_id(cores_100_io_prev_bits_id),
    .io_next_ready(cores_100_io_next_ready),
    .io_next_valid(cores_100_io_next_valid),
    .io_next_bits_address(cores_100_io_next_bits_address),
    .io_next_bits_data(cores_100_io_next_bits_data),
    .io_next_bits_wen(cores_100_io_next_bits_wen),
    .io_next_bits_id(cores_100_io_next_bits_id)
  );
  RingCore_101 cores_101 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_101_clock),
    .reset(cores_101_reset),
    .io_prev_ready(cores_101_io_prev_ready),
    .io_prev_valid(cores_101_io_prev_valid),
    .io_prev_bits_address(cores_101_io_prev_bits_address),
    .io_prev_bits_data(cores_101_io_prev_bits_data),
    .io_prev_bits_wen(cores_101_io_prev_bits_wen),
    .io_prev_bits_id(cores_101_io_prev_bits_id),
    .io_next_ready(cores_101_io_next_ready),
    .io_next_valid(cores_101_io_next_valid),
    .io_next_bits_address(cores_101_io_next_bits_address),
    .io_next_bits_data(cores_101_io_next_bits_data),
    .io_next_bits_wen(cores_101_io_next_bits_wen),
    .io_next_bits_id(cores_101_io_next_bits_id)
  );
  RingCore_102 cores_102 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_102_clock),
    .reset(cores_102_reset),
    .io_prev_ready(cores_102_io_prev_ready),
    .io_prev_valid(cores_102_io_prev_valid),
    .io_prev_bits_address(cores_102_io_prev_bits_address),
    .io_prev_bits_data(cores_102_io_prev_bits_data),
    .io_prev_bits_wen(cores_102_io_prev_bits_wen),
    .io_prev_bits_id(cores_102_io_prev_bits_id),
    .io_next_ready(cores_102_io_next_ready),
    .io_next_valid(cores_102_io_next_valid),
    .io_next_bits_address(cores_102_io_next_bits_address),
    .io_next_bits_data(cores_102_io_next_bits_data),
    .io_next_bits_wen(cores_102_io_next_bits_wen),
    .io_next_bits_id(cores_102_io_next_bits_id)
  );
  RingCore_103 cores_103 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_103_clock),
    .reset(cores_103_reset),
    .io_prev_ready(cores_103_io_prev_ready),
    .io_prev_valid(cores_103_io_prev_valid),
    .io_prev_bits_address(cores_103_io_prev_bits_address),
    .io_prev_bits_data(cores_103_io_prev_bits_data),
    .io_prev_bits_wen(cores_103_io_prev_bits_wen),
    .io_prev_bits_id(cores_103_io_prev_bits_id),
    .io_next_ready(cores_103_io_next_ready),
    .io_next_valid(cores_103_io_next_valid),
    .io_next_bits_address(cores_103_io_next_bits_address),
    .io_next_bits_data(cores_103_io_next_bits_data),
    .io_next_bits_wen(cores_103_io_next_bits_wen),
    .io_next_bits_id(cores_103_io_next_bits_id)
  );
  RingCore_104 cores_104 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_104_clock),
    .reset(cores_104_reset),
    .io_prev_ready(cores_104_io_prev_ready),
    .io_prev_valid(cores_104_io_prev_valid),
    .io_prev_bits_address(cores_104_io_prev_bits_address),
    .io_prev_bits_data(cores_104_io_prev_bits_data),
    .io_prev_bits_wen(cores_104_io_prev_bits_wen),
    .io_prev_bits_id(cores_104_io_prev_bits_id),
    .io_next_ready(cores_104_io_next_ready),
    .io_next_valid(cores_104_io_next_valid),
    .io_next_bits_address(cores_104_io_next_bits_address),
    .io_next_bits_data(cores_104_io_next_bits_data),
    .io_next_bits_wen(cores_104_io_next_bits_wen),
    .io_next_bits_id(cores_104_io_next_bits_id)
  );
  RingCore_105 cores_105 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_105_clock),
    .reset(cores_105_reset),
    .io_prev_ready(cores_105_io_prev_ready),
    .io_prev_valid(cores_105_io_prev_valid),
    .io_prev_bits_address(cores_105_io_prev_bits_address),
    .io_prev_bits_data(cores_105_io_prev_bits_data),
    .io_prev_bits_wen(cores_105_io_prev_bits_wen),
    .io_prev_bits_id(cores_105_io_prev_bits_id),
    .io_next_ready(cores_105_io_next_ready),
    .io_next_valid(cores_105_io_next_valid),
    .io_next_bits_address(cores_105_io_next_bits_address),
    .io_next_bits_data(cores_105_io_next_bits_data),
    .io_next_bits_wen(cores_105_io_next_bits_wen),
    .io_next_bits_id(cores_105_io_next_bits_id)
  );
  RingCore_106 cores_106 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_106_clock),
    .reset(cores_106_reset),
    .io_prev_ready(cores_106_io_prev_ready),
    .io_prev_valid(cores_106_io_prev_valid),
    .io_prev_bits_address(cores_106_io_prev_bits_address),
    .io_prev_bits_data(cores_106_io_prev_bits_data),
    .io_prev_bits_wen(cores_106_io_prev_bits_wen),
    .io_prev_bits_id(cores_106_io_prev_bits_id),
    .io_next_ready(cores_106_io_next_ready),
    .io_next_valid(cores_106_io_next_valid),
    .io_next_bits_address(cores_106_io_next_bits_address),
    .io_next_bits_data(cores_106_io_next_bits_data),
    .io_next_bits_wen(cores_106_io_next_bits_wen),
    .io_next_bits_id(cores_106_io_next_bits_id)
  );
  RingCore_107 cores_107 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_107_clock),
    .reset(cores_107_reset),
    .io_prev_ready(cores_107_io_prev_ready),
    .io_prev_valid(cores_107_io_prev_valid),
    .io_prev_bits_address(cores_107_io_prev_bits_address),
    .io_prev_bits_data(cores_107_io_prev_bits_data),
    .io_prev_bits_wen(cores_107_io_prev_bits_wen),
    .io_prev_bits_id(cores_107_io_prev_bits_id),
    .io_next_ready(cores_107_io_next_ready),
    .io_next_valid(cores_107_io_next_valid),
    .io_next_bits_address(cores_107_io_next_bits_address),
    .io_next_bits_data(cores_107_io_next_bits_data),
    .io_next_bits_wen(cores_107_io_next_bits_wen),
    .io_next_bits_id(cores_107_io_next_bits_id)
  );
  RingCore_108 cores_108 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_108_clock),
    .reset(cores_108_reset),
    .io_prev_ready(cores_108_io_prev_ready),
    .io_prev_valid(cores_108_io_prev_valid),
    .io_prev_bits_address(cores_108_io_prev_bits_address),
    .io_prev_bits_data(cores_108_io_prev_bits_data),
    .io_prev_bits_wen(cores_108_io_prev_bits_wen),
    .io_prev_bits_id(cores_108_io_prev_bits_id),
    .io_next_ready(cores_108_io_next_ready),
    .io_next_valid(cores_108_io_next_valid),
    .io_next_bits_address(cores_108_io_next_bits_address),
    .io_next_bits_data(cores_108_io_next_bits_data),
    .io_next_bits_wen(cores_108_io_next_bits_wen),
    .io_next_bits_id(cores_108_io_next_bits_id)
  );
  RingCore_109 cores_109 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_109_clock),
    .reset(cores_109_reset),
    .io_prev_ready(cores_109_io_prev_ready),
    .io_prev_valid(cores_109_io_prev_valid),
    .io_prev_bits_address(cores_109_io_prev_bits_address),
    .io_prev_bits_data(cores_109_io_prev_bits_data),
    .io_prev_bits_wen(cores_109_io_prev_bits_wen),
    .io_prev_bits_id(cores_109_io_prev_bits_id),
    .io_next_ready(cores_109_io_next_ready),
    .io_next_valid(cores_109_io_next_valid),
    .io_next_bits_address(cores_109_io_next_bits_address),
    .io_next_bits_data(cores_109_io_next_bits_data),
    .io_next_bits_wen(cores_109_io_next_bits_wen),
    .io_next_bits_id(cores_109_io_next_bits_id)
  );
  RingCore_110 cores_110 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_110_clock),
    .reset(cores_110_reset),
    .io_prev_ready(cores_110_io_prev_ready),
    .io_prev_valid(cores_110_io_prev_valid),
    .io_prev_bits_address(cores_110_io_prev_bits_address),
    .io_prev_bits_data(cores_110_io_prev_bits_data),
    .io_prev_bits_wen(cores_110_io_prev_bits_wen),
    .io_prev_bits_id(cores_110_io_prev_bits_id),
    .io_next_ready(cores_110_io_next_ready),
    .io_next_valid(cores_110_io_next_valid),
    .io_next_bits_address(cores_110_io_next_bits_address),
    .io_next_bits_data(cores_110_io_next_bits_data),
    .io_next_bits_wen(cores_110_io_next_bits_wen),
    .io_next_bits_id(cores_110_io_next_bits_id)
  );
  RingCore_111 cores_111 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_111_clock),
    .reset(cores_111_reset),
    .io_prev_ready(cores_111_io_prev_ready),
    .io_prev_valid(cores_111_io_prev_valid),
    .io_prev_bits_address(cores_111_io_prev_bits_address),
    .io_prev_bits_data(cores_111_io_prev_bits_data),
    .io_prev_bits_wen(cores_111_io_prev_bits_wen),
    .io_prev_bits_id(cores_111_io_prev_bits_id),
    .io_next_ready(cores_111_io_next_ready),
    .io_next_valid(cores_111_io_next_valid),
    .io_next_bits_address(cores_111_io_next_bits_address),
    .io_next_bits_data(cores_111_io_next_bits_data),
    .io_next_bits_wen(cores_111_io_next_bits_wen),
    .io_next_bits_id(cores_111_io_next_bits_id)
  );
  RingCore_112 cores_112 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_112_clock),
    .reset(cores_112_reset),
    .io_prev_ready(cores_112_io_prev_ready),
    .io_prev_valid(cores_112_io_prev_valid),
    .io_prev_bits_address(cores_112_io_prev_bits_address),
    .io_prev_bits_data(cores_112_io_prev_bits_data),
    .io_prev_bits_wen(cores_112_io_prev_bits_wen),
    .io_prev_bits_id(cores_112_io_prev_bits_id),
    .io_next_ready(cores_112_io_next_ready),
    .io_next_valid(cores_112_io_next_valid),
    .io_next_bits_address(cores_112_io_next_bits_address),
    .io_next_bits_data(cores_112_io_next_bits_data),
    .io_next_bits_wen(cores_112_io_next_bits_wen),
    .io_next_bits_id(cores_112_io_next_bits_id)
  );
  RingCore_113 cores_113 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_113_clock),
    .reset(cores_113_reset),
    .io_prev_ready(cores_113_io_prev_ready),
    .io_prev_valid(cores_113_io_prev_valid),
    .io_prev_bits_address(cores_113_io_prev_bits_address),
    .io_prev_bits_data(cores_113_io_prev_bits_data),
    .io_prev_bits_wen(cores_113_io_prev_bits_wen),
    .io_prev_bits_id(cores_113_io_prev_bits_id),
    .io_next_ready(cores_113_io_next_ready),
    .io_next_valid(cores_113_io_next_valid),
    .io_next_bits_address(cores_113_io_next_bits_address),
    .io_next_bits_data(cores_113_io_next_bits_data),
    .io_next_bits_wen(cores_113_io_next_bits_wen),
    .io_next_bits_id(cores_113_io_next_bits_id)
  );
  RingCore_114 cores_114 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_114_clock),
    .reset(cores_114_reset),
    .io_prev_ready(cores_114_io_prev_ready),
    .io_prev_valid(cores_114_io_prev_valid),
    .io_prev_bits_address(cores_114_io_prev_bits_address),
    .io_prev_bits_data(cores_114_io_prev_bits_data),
    .io_prev_bits_wen(cores_114_io_prev_bits_wen),
    .io_prev_bits_id(cores_114_io_prev_bits_id),
    .io_next_ready(cores_114_io_next_ready),
    .io_next_valid(cores_114_io_next_valid),
    .io_next_bits_address(cores_114_io_next_bits_address),
    .io_next_bits_data(cores_114_io_next_bits_data),
    .io_next_bits_wen(cores_114_io_next_bits_wen),
    .io_next_bits_id(cores_114_io_next_bits_id)
  );
  RingCore_115 cores_115 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_115_clock),
    .reset(cores_115_reset),
    .io_prev_ready(cores_115_io_prev_ready),
    .io_prev_valid(cores_115_io_prev_valid),
    .io_prev_bits_address(cores_115_io_prev_bits_address),
    .io_prev_bits_data(cores_115_io_prev_bits_data),
    .io_prev_bits_wen(cores_115_io_prev_bits_wen),
    .io_prev_bits_id(cores_115_io_prev_bits_id),
    .io_next_ready(cores_115_io_next_ready),
    .io_next_valid(cores_115_io_next_valid),
    .io_next_bits_address(cores_115_io_next_bits_address),
    .io_next_bits_data(cores_115_io_next_bits_data),
    .io_next_bits_wen(cores_115_io_next_bits_wen),
    .io_next_bits_id(cores_115_io_next_bits_id)
  );
  RingCore_116 cores_116 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_116_clock),
    .reset(cores_116_reset),
    .io_prev_ready(cores_116_io_prev_ready),
    .io_prev_valid(cores_116_io_prev_valid),
    .io_prev_bits_address(cores_116_io_prev_bits_address),
    .io_prev_bits_data(cores_116_io_prev_bits_data),
    .io_prev_bits_wen(cores_116_io_prev_bits_wen),
    .io_prev_bits_id(cores_116_io_prev_bits_id),
    .io_next_ready(cores_116_io_next_ready),
    .io_next_valid(cores_116_io_next_valid),
    .io_next_bits_address(cores_116_io_next_bits_address),
    .io_next_bits_data(cores_116_io_next_bits_data),
    .io_next_bits_wen(cores_116_io_next_bits_wen),
    .io_next_bits_id(cores_116_io_next_bits_id)
  );
  RingCore_117 cores_117 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_117_clock),
    .reset(cores_117_reset),
    .io_prev_ready(cores_117_io_prev_ready),
    .io_prev_valid(cores_117_io_prev_valid),
    .io_prev_bits_address(cores_117_io_prev_bits_address),
    .io_prev_bits_data(cores_117_io_prev_bits_data),
    .io_prev_bits_wen(cores_117_io_prev_bits_wen),
    .io_prev_bits_id(cores_117_io_prev_bits_id),
    .io_next_ready(cores_117_io_next_ready),
    .io_next_valid(cores_117_io_next_valid),
    .io_next_bits_address(cores_117_io_next_bits_address),
    .io_next_bits_data(cores_117_io_next_bits_data),
    .io_next_bits_wen(cores_117_io_next_bits_wen),
    .io_next_bits_id(cores_117_io_next_bits_id)
  );
  RingCore_118 cores_118 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_118_clock),
    .reset(cores_118_reset),
    .io_prev_ready(cores_118_io_prev_ready),
    .io_prev_valid(cores_118_io_prev_valid),
    .io_prev_bits_address(cores_118_io_prev_bits_address),
    .io_prev_bits_data(cores_118_io_prev_bits_data),
    .io_prev_bits_wen(cores_118_io_prev_bits_wen),
    .io_prev_bits_id(cores_118_io_prev_bits_id),
    .io_next_ready(cores_118_io_next_ready),
    .io_next_valid(cores_118_io_next_valid),
    .io_next_bits_address(cores_118_io_next_bits_address),
    .io_next_bits_data(cores_118_io_next_bits_data),
    .io_next_bits_wen(cores_118_io_next_bits_wen),
    .io_next_bits_id(cores_118_io_next_bits_id)
  );
  RingCore_119 cores_119 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_119_clock),
    .reset(cores_119_reset),
    .io_prev_ready(cores_119_io_prev_ready),
    .io_prev_valid(cores_119_io_prev_valid),
    .io_prev_bits_address(cores_119_io_prev_bits_address),
    .io_prev_bits_data(cores_119_io_prev_bits_data),
    .io_prev_bits_wen(cores_119_io_prev_bits_wen),
    .io_prev_bits_id(cores_119_io_prev_bits_id),
    .io_next_ready(cores_119_io_next_ready),
    .io_next_valid(cores_119_io_next_valid),
    .io_next_bits_address(cores_119_io_next_bits_address),
    .io_next_bits_data(cores_119_io_next_bits_data),
    .io_next_bits_wen(cores_119_io_next_bits_wen),
    .io_next_bits_id(cores_119_io_next_bits_id)
  );
  RingCore_120 cores_120 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_120_clock),
    .reset(cores_120_reset),
    .io_prev_ready(cores_120_io_prev_ready),
    .io_prev_valid(cores_120_io_prev_valid),
    .io_prev_bits_address(cores_120_io_prev_bits_address),
    .io_prev_bits_data(cores_120_io_prev_bits_data),
    .io_prev_bits_wen(cores_120_io_prev_bits_wen),
    .io_prev_bits_id(cores_120_io_prev_bits_id),
    .io_next_ready(cores_120_io_next_ready),
    .io_next_valid(cores_120_io_next_valid),
    .io_next_bits_address(cores_120_io_next_bits_address),
    .io_next_bits_data(cores_120_io_next_bits_data),
    .io_next_bits_wen(cores_120_io_next_bits_wen),
    .io_next_bits_id(cores_120_io_next_bits_id)
  );
  RingCore_121 cores_121 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_121_clock),
    .reset(cores_121_reset),
    .io_prev_ready(cores_121_io_prev_ready),
    .io_prev_valid(cores_121_io_prev_valid),
    .io_prev_bits_address(cores_121_io_prev_bits_address),
    .io_prev_bits_data(cores_121_io_prev_bits_data),
    .io_prev_bits_wen(cores_121_io_prev_bits_wen),
    .io_prev_bits_id(cores_121_io_prev_bits_id),
    .io_next_ready(cores_121_io_next_ready),
    .io_next_valid(cores_121_io_next_valid),
    .io_next_bits_address(cores_121_io_next_bits_address),
    .io_next_bits_data(cores_121_io_next_bits_data),
    .io_next_bits_wen(cores_121_io_next_bits_wen),
    .io_next_bits_id(cores_121_io_next_bits_id)
  );
  RingCore_122 cores_122 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_122_clock),
    .reset(cores_122_reset),
    .io_prev_ready(cores_122_io_prev_ready),
    .io_prev_valid(cores_122_io_prev_valid),
    .io_prev_bits_address(cores_122_io_prev_bits_address),
    .io_prev_bits_data(cores_122_io_prev_bits_data),
    .io_prev_bits_wen(cores_122_io_prev_bits_wen),
    .io_prev_bits_id(cores_122_io_prev_bits_id),
    .io_next_ready(cores_122_io_next_ready),
    .io_next_valid(cores_122_io_next_valid),
    .io_next_bits_address(cores_122_io_next_bits_address),
    .io_next_bits_data(cores_122_io_next_bits_data),
    .io_next_bits_wen(cores_122_io_next_bits_wen),
    .io_next_bits_id(cores_122_io_next_bits_id)
  );
  RingCore_123 cores_123 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_123_clock),
    .reset(cores_123_reset),
    .io_prev_ready(cores_123_io_prev_ready),
    .io_prev_valid(cores_123_io_prev_valid),
    .io_prev_bits_address(cores_123_io_prev_bits_address),
    .io_prev_bits_data(cores_123_io_prev_bits_data),
    .io_prev_bits_wen(cores_123_io_prev_bits_wen),
    .io_prev_bits_id(cores_123_io_prev_bits_id),
    .io_next_ready(cores_123_io_next_ready),
    .io_next_valid(cores_123_io_next_valid),
    .io_next_bits_address(cores_123_io_next_bits_address),
    .io_next_bits_data(cores_123_io_next_bits_data),
    .io_next_bits_wen(cores_123_io_next_bits_wen),
    .io_next_bits_id(cores_123_io_next_bits_id)
  );
  RingCore_124 cores_124 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_124_clock),
    .reset(cores_124_reset),
    .io_prev_ready(cores_124_io_prev_ready),
    .io_prev_valid(cores_124_io_prev_valid),
    .io_prev_bits_address(cores_124_io_prev_bits_address),
    .io_prev_bits_data(cores_124_io_prev_bits_data),
    .io_prev_bits_wen(cores_124_io_prev_bits_wen),
    .io_prev_bits_id(cores_124_io_prev_bits_id),
    .io_next_ready(cores_124_io_next_ready),
    .io_next_valid(cores_124_io_next_valid),
    .io_next_bits_address(cores_124_io_next_bits_address),
    .io_next_bits_data(cores_124_io_next_bits_data),
    .io_next_bits_wen(cores_124_io_next_bits_wen),
    .io_next_bits_id(cores_124_io_next_bits_id)
  );
  RingCore_125 cores_125 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_125_clock),
    .reset(cores_125_reset),
    .io_prev_ready(cores_125_io_prev_ready),
    .io_prev_valid(cores_125_io_prev_valid),
    .io_prev_bits_address(cores_125_io_prev_bits_address),
    .io_prev_bits_data(cores_125_io_prev_bits_data),
    .io_prev_bits_wen(cores_125_io_prev_bits_wen),
    .io_prev_bits_id(cores_125_io_prev_bits_id),
    .io_next_ready(cores_125_io_next_ready),
    .io_next_valid(cores_125_io_next_valid),
    .io_next_bits_address(cores_125_io_next_bits_address),
    .io_next_bits_data(cores_125_io_next_bits_data),
    .io_next_bits_wen(cores_125_io_next_bits_wen),
    .io_next_bits_id(cores_125_io_next_bits_id)
  );
  RingCore_126 cores_126 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_126_clock),
    .reset(cores_126_reset),
    .io_prev_ready(cores_126_io_prev_ready),
    .io_prev_valid(cores_126_io_prev_valid),
    .io_prev_bits_address(cores_126_io_prev_bits_address),
    .io_prev_bits_data(cores_126_io_prev_bits_data),
    .io_prev_bits_wen(cores_126_io_prev_bits_wen),
    .io_prev_bits_id(cores_126_io_prev_bits_id),
    .io_next_ready(cores_126_io_next_ready),
    .io_next_valid(cores_126_io_next_valid),
    .io_next_bits_address(cores_126_io_next_bits_address),
    .io_next_bits_data(cores_126_io_next_bits_data),
    .io_next_bits_wen(cores_126_io_next_bits_wen),
    .io_next_bits_id(cores_126_io_next_bits_id)
  );
  RingCore_127 cores_127 ( // @[FemtoMips32.scala 470:51]
    .clock(cores_127_clock),
    .reset(cores_127_reset),
    .io_prev_ready(cores_127_io_prev_ready),
    .io_prev_valid(cores_127_io_prev_valid),
    .io_prev_bits_address(cores_127_io_prev_bits_address),
    .io_prev_bits_data(cores_127_io_prev_bits_data),
    .io_prev_bits_wen(cores_127_io_prev_bits_wen),
    .io_prev_bits_id(cores_127_io_prev_bits_id),
    .io_next_ready(cores_127_io_next_ready),
    .io_next_valid(cores_127_io_next_valid),
    .io_next_bits_address(cores_127_io_next_bits_address),
    .io_next_bits_data(cores_127_io_next_bits_data),
    .io_next_bits_wen(cores_127_io_next_bits_wen),
    .io_next_bits_id(cores_127_io_next_bits_id)
  );
  assign io_prev_ready = cores_0_io_prev_ready; // @[FemtoMips32.scala 477:11]
  assign io_next_valid = cores_127_io_next_valid; // @[FemtoMips32.scala 478:22]
  assign io_next_bits_address = cores_127_io_next_bits_address; // @[FemtoMips32.scala 478:22]
  assign io_next_bits_data = cores_127_io_next_bits_data; // @[FemtoMips32.scala 478:22]
  assign io_next_bits_wen = cores_127_io_next_bits_wen; // @[FemtoMips32.scala 478:22]
  assign io_next_bits_id = cores_127_io_next_bits_id; // @[FemtoMips32.scala 478:22]
  assign io_halted = 1'h0; // @[FemtoMips32.scala 476:13]
  assign cores_0_clock = clock;
  assign cores_0_reset = reset;
  assign cores_0_io_prev_valid = io_prev_valid; // @[FemtoMips32.scala 477:11]
  assign cores_0_io_prev_bits_address = io_prev_bits_address; // @[FemtoMips32.scala 477:11]
  assign cores_0_io_prev_bits_data = io_prev_bits_data; // @[FemtoMips32.scala 477:11]
  assign cores_0_io_prev_bits_wen = io_prev_bits_wen; // @[FemtoMips32.scala 477:11]
  assign cores_0_io_prev_bits_id = io_prev_bits_id; // @[FemtoMips32.scala 477:11]
  assign cores_0_io_next_ready = cores_1_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_1_clock = clock;
  assign cores_1_reset = reset;
  assign cores_1_io_prev_valid = cores_0_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_1_io_prev_bits_address = cores_0_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_1_io_prev_bits_data = cores_0_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_1_io_prev_bits_wen = cores_0_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_1_io_prev_bits_id = cores_0_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_1_io_next_ready = cores_2_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_2_clock = clock;
  assign cores_2_reset = reset;
  assign cores_2_io_prev_valid = cores_1_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_2_io_prev_bits_address = cores_1_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_2_io_prev_bits_data = cores_1_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_2_io_prev_bits_wen = cores_1_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_2_io_prev_bits_id = cores_1_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_2_io_next_ready = cores_3_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_3_clock = clock;
  assign cores_3_reset = reset;
  assign cores_3_io_prev_valid = cores_2_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_3_io_prev_bits_address = cores_2_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_3_io_prev_bits_data = cores_2_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_3_io_prev_bits_wen = cores_2_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_3_io_prev_bits_id = cores_2_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_3_io_next_ready = cores_4_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_4_clock = clock;
  assign cores_4_reset = reset;
  assign cores_4_io_prev_valid = cores_3_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_4_io_prev_bits_address = cores_3_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_4_io_prev_bits_data = cores_3_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_4_io_prev_bits_wen = cores_3_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_4_io_prev_bits_id = cores_3_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_4_io_next_ready = cores_5_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_5_clock = clock;
  assign cores_5_reset = reset;
  assign cores_5_io_prev_valid = cores_4_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_5_io_prev_bits_address = cores_4_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_5_io_prev_bits_data = cores_4_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_5_io_prev_bits_wen = cores_4_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_5_io_prev_bits_id = cores_4_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_5_io_next_ready = cores_6_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_6_clock = clock;
  assign cores_6_reset = reset;
  assign cores_6_io_prev_valid = cores_5_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_6_io_prev_bits_address = cores_5_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_6_io_prev_bits_data = cores_5_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_6_io_prev_bits_wen = cores_5_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_6_io_prev_bits_id = cores_5_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_6_io_next_ready = cores_7_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_7_clock = clock;
  assign cores_7_reset = reset;
  assign cores_7_io_prev_valid = cores_6_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_7_io_prev_bits_address = cores_6_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_7_io_prev_bits_data = cores_6_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_7_io_prev_bits_wen = cores_6_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_7_io_prev_bits_id = cores_6_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_7_io_next_ready = cores_8_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_8_clock = clock;
  assign cores_8_reset = reset;
  assign cores_8_io_prev_valid = cores_7_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_8_io_prev_bits_address = cores_7_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_8_io_prev_bits_data = cores_7_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_8_io_prev_bits_wen = cores_7_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_8_io_prev_bits_id = cores_7_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_8_io_next_ready = cores_9_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_9_clock = clock;
  assign cores_9_reset = reset;
  assign cores_9_io_prev_valid = cores_8_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_9_io_prev_bits_address = cores_8_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_9_io_prev_bits_data = cores_8_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_9_io_prev_bits_wen = cores_8_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_9_io_prev_bits_id = cores_8_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_9_io_next_ready = cores_10_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_10_clock = clock;
  assign cores_10_reset = reset;
  assign cores_10_io_prev_valid = cores_9_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_10_io_prev_bits_address = cores_9_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_10_io_prev_bits_data = cores_9_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_10_io_prev_bits_wen = cores_9_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_10_io_prev_bits_id = cores_9_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_10_io_next_ready = cores_11_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_11_clock = clock;
  assign cores_11_reset = reset;
  assign cores_11_io_prev_valid = cores_10_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_11_io_prev_bits_address = cores_10_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_11_io_prev_bits_data = cores_10_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_11_io_prev_bits_wen = cores_10_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_11_io_prev_bits_id = cores_10_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_11_io_next_ready = cores_12_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_12_clock = clock;
  assign cores_12_reset = reset;
  assign cores_12_io_prev_valid = cores_11_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_12_io_prev_bits_address = cores_11_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_12_io_prev_bits_data = cores_11_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_12_io_prev_bits_wen = cores_11_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_12_io_prev_bits_id = cores_11_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_12_io_next_ready = cores_13_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_13_clock = clock;
  assign cores_13_reset = reset;
  assign cores_13_io_prev_valid = cores_12_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_13_io_prev_bits_address = cores_12_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_13_io_prev_bits_data = cores_12_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_13_io_prev_bits_wen = cores_12_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_13_io_prev_bits_id = cores_12_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_13_io_next_ready = cores_14_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_14_clock = clock;
  assign cores_14_reset = reset;
  assign cores_14_io_prev_valid = cores_13_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_14_io_prev_bits_address = cores_13_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_14_io_prev_bits_data = cores_13_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_14_io_prev_bits_wen = cores_13_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_14_io_prev_bits_id = cores_13_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_14_io_next_ready = cores_15_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_15_clock = clock;
  assign cores_15_reset = reset;
  assign cores_15_io_prev_valid = cores_14_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_15_io_prev_bits_address = cores_14_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_15_io_prev_bits_data = cores_14_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_15_io_prev_bits_wen = cores_14_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_15_io_prev_bits_id = cores_14_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_15_io_next_ready = cores_16_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_16_clock = clock;
  assign cores_16_reset = reset;
  assign cores_16_io_prev_valid = cores_15_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_16_io_prev_bits_address = cores_15_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_16_io_prev_bits_data = cores_15_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_16_io_prev_bits_wen = cores_15_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_16_io_prev_bits_id = cores_15_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_16_io_next_ready = cores_17_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_17_clock = clock;
  assign cores_17_reset = reset;
  assign cores_17_io_prev_valid = cores_16_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_17_io_prev_bits_address = cores_16_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_17_io_prev_bits_data = cores_16_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_17_io_prev_bits_wen = cores_16_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_17_io_prev_bits_id = cores_16_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_17_io_next_ready = cores_18_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_18_clock = clock;
  assign cores_18_reset = reset;
  assign cores_18_io_prev_valid = cores_17_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_18_io_prev_bits_address = cores_17_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_18_io_prev_bits_data = cores_17_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_18_io_prev_bits_wen = cores_17_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_18_io_prev_bits_id = cores_17_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_18_io_next_ready = cores_19_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_19_clock = clock;
  assign cores_19_reset = reset;
  assign cores_19_io_prev_valid = cores_18_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_19_io_prev_bits_address = cores_18_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_19_io_prev_bits_data = cores_18_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_19_io_prev_bits_wen = cores_18_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_19_io_prev_bits_id = cores_18_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_19_io_next_ready = cores_20_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_20_clock = clock;
  assign cores_20_reset = reset;
  assign cores_20_io_prev_valid = cores_19_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_20_io_prev_bits_address = cores_19_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_20_io_prev_bits_data = cores_19_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_20_io_prev_bits_wen = cores_19_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_20_io_prev_bits_id = cores_19_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_20_io_next_ready = cores_21_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_21_clock = clock;
  assign cores_21_reset = reset;
  assign cores_21_io_prev_valid = cores_20_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_21_io_prev_bits_address = cores_20_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_21_io_prev_bits_data = cores_20_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_21_io_prev_bits_wen = cores_20_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_21_io_prev_bits_id = cores_20_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_21_io_next_ready = cores_22_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_22_clock = clock;
  assign cores_22_reset = reset;
  assign cores_22_io_prev_valid = cores_21_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_22_io_prev_bits_address = cores_21_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_22_io_prev_bits_data = cores_21_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_22_io_prev_bits_wen = cores_21_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_22_io_prev_bits_id = cores_21_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_22_io_next_ready = cores_23_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_23_clock = clock;
  assign cores_23_reset = reset;
  assign cores_23_io_prev_valid = cores_22_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_23_io_prev_bits_address = cores_22_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_23_io_prev_bits_data = cores_22_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_23_io_prev_bits_wen = cores_22_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_23_io_prev_bits_id = cores_22_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_23_io_next_ready = cores_24_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_24_clock = clock;
  assign cores_24_reset = reset;
  assign cores_24_io_prev_valid = cores_23_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_24_io_prev_bits_address = cores_23_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_24_io_prev_bits_data = cores_23_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_24_io_prev_bits_wen = cores_23_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_24_io_prev_bits_id = cores_23_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_24_io_next_ready = cores_25_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_25_clock = clock;
  assign cores_25_reset = reset;
  assign cores_25_io_prev_valid = cores_24_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_25_io_prev_bits_address = cores_24_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_25_io_prev_bits_data = cores_24_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_25_io_prev_bits_wen = cores_24_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_25_io_prev_bits_id = cores_24_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_25_io_next_ready = cores_26_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_26_clock = clock;
  assign cores_26_reset = reset;
  assign cores_26_io_prev_valid = cores_25_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_26_io_prev_bits_address = cores_25_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_26_io_prev_bits_data = cores_25_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_26_io_prev_bits_wen = cores_25_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_26_io_prev_bits_id = cores_25_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_26_io_next_ready = cores_27_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_27_clock = clock;
  assign cores_27_reset = reset;
  assign cores_27_io_prev_valid = cores_26_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_27_io_prev_bits_address = cores_26_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_27_io_prev_bits_data = cores_26_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_27_io_prev_bits_wen = cores_26_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_27_io_prev_bits_id = cores_26_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_27_io_next_ready = cores_28_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_28_clock = clock;
  assign cores_28_reset = reset;
  assign cores_28_io_prev_valid = cores_27_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_28_io_prev_bits_address = cores_27_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_28_io_prev_bits_data = cores_27_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_28_io_prev_bits_wen = cores_27_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_28_io_prev_bits_id = cores_27_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_28_io_next_ready = cores_29_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_29_clock = clock;
  assign cores_29_reset = reset;
  assign cores_29_io_prev_valid = cores_28_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_29_io_prev_bits_address = cores_28_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_29_io_prev_bits_data = cores_28_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_29_io_prev_bits_wen = cores_28_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_29_io_prev_bits_id = cores_28_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_29_io_next_ready = cores_30_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_30_clock = clock;
  assign cores_30_reset = reset;
  assign cores_30_io_prev_valid = cores_29_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_30_io_prev_bits_address = cores_29_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_30_io_prev_bits_data = cores_29_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_30_io_prev_bits_wen = cores_29_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_30_io_prev_bits_id = cores_29_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_30_io_next_ready = cores_31_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_31_clock = clock;
  assign cores_31_reset = reset;
  assign cores_31_io_prev_valid = cores_30_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_31_io_prev_bits_address = cores_30_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_31_io_prev_bits_data = cores_30_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_31_io_prev_bits_wen = cores_30_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_31_io_prev_bits_id = cores_30_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_31_io_next_ready = cores_32_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_32_clock = clock;
  assign cores_32_reset = reset;
  assign cores_32_io_prev_valid = cores_31_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_32_io_prev_bits_address = cores_31_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_32_io_prev_bits_data = cores_31_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_32_io_prev_bits_wen = cores_31_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_32_io_prev_bits_id = cores_31_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_32_io_next_ready = cores_33_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_33_clock = clock;
  assign cores_33_reset = reset;
  assign cores_33_io_prev_valid = cores_32_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_33_io_prev_bits_address = cores_32_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_33_io_prev_bits_data = cores_32_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_33_io_prev_bits_wen = cores_32_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_33_io_prev_bits_id = cores_32_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_33_io_next_ready = cores_34_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_34_clock = clock;
  assign cores_34_reset = reset;
  assign cores_34_io_prev_valid = cores_33_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_34_io_prev_bits_address = cores_33_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_34_io_prev_bits_data = cores_33_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_34_io_prev_bits_wen = cores_33_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_34_io_prev_bits_id = cores_33_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_34_io_next_ready = cores_35_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_35_clock = clock;
  assign cores_35_reset = reset;
  assign cores_35_io_prev_valid = cores_34_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_35_io_prev_bits_address = cores_34_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_35_io_prev_bits_data = cores_34_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_35_io_prev_bits_wen = cores_34_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_35_io_prev_bits_id = cores_34_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_35_io_next_ready = cores_36_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_36_clock = clock;
  assign cores_36_reset = reset;
  assign cores_36_io_prev_valid = cores_35_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_36_io_prev_bits_address = cores_35_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_36_io_prev_bits_data = cores_35_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_36_io_prev_bits_wen = cores_35_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_36_io_prev_bits_id = cores_35_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_36_io_next_ready = cores_37_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_37_clock = clock;
  assign cores_37_reset = reset;
  assign cores_37_io_prev_valid = cores_36_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_37_io_prev_bits_address = cores_36_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_37_io_prev_bits_data = cores_36_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_37_io_prev_bits_wen = cores_36_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_37_io_prev_bits_id = cores_36_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_37_io_next_ready = cores_38_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_38_clock = clock;
  assign cores_38_reset = reset;
  assign cores_38_io_prev_valid = cores_37_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_38_io_prev_bits_address = cores_37_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_38_io_prev_bits_data = cores_37_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_38_io_prev_bits_wen = cores_37_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_38_io_prev_bits_id = cores_37_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_38_io_next_ready = cores_39_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_39_clock = clock;
  assign cores_39_reset = reset;
  assign cores_39_io_prev_valid = cores_38_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_39_io_prev_bits_address = cores_38_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_39_io_prev_bits_data = cores_38_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_39_io_prev_bits_wen = cores_38_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_39_io_prev_bits_id = cores_38_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_39_io_next_ready = cores_40_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_40_clock = clock;
  assign cores_40_reset = reset;
  assign cores_40_io_prev_valid = cores_39_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_40_io_prev_bits_address = cores_39_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_40_io_prev_bits_data = cores_39_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_40_io_prev_bits_wen = cores_39_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_40_io_prev_bits_id = cores_39_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_40_io_next_ready = cores_41_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_41_clock = clock;
  assign cores_41_reset = reset;
  assign cores_41_io_prev_valid = cores_40_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_41_io_prev_bits_address = cores_40_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_41_io_prev_bits_data = cores_40_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_41_io_prev_bits_wen = cores_40_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_41_io_prev_bits_id = cores_40_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_41_io_next_ready = cores_42_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_42_clock = clock;
  assign cores_42_reset = reset;
  assign cores_42_io_prev_valid = cores_41_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_42_io_prev_bits_address = cores_41_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_42_io_prev_bits_data = cores_41_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_42_io_prev_bits_wen = cores_41_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_42_io_prev_bits_id = cores_41_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_42_io_next_ready = cores_43_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_43_clock = clock;
  assign cores_43_reset = reset;
  assign cores_43_io_prev_valid = cores_42_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_43_io_prev_bits_address = cores_42_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_43_io_prev_bits_data = cores_42_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_43_io_prev_bits_wen = cores_42_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_43_io_prev_bits_id = cores_42_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_43_io_next_ready = cores_44_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_44_clock = clock;
  assign cores_44_reset = reset;
  assign cores_44_io_prev_valid = cores_43_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_44_io_prev_bits_address = cores_43_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_44_io_prev_bits_data = cores_43_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_44_io_prev_bits_wen = cores_43_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_44_io_prev_bits_id = cores_43_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_44_io_next_ready = cores_45_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_45_clock = clock;
  assign cores_45_reset = reset;
  assign cores_45_io_prev_valid = cores_44_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_45_io_prev_bits_address = cores_44_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_45_io_prev_bits_data = cores_44_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_45_io_prev_bits_wen = cores_44_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_45_io_prev_bits_id = cores_44_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_45_io_next_ready = cores_46_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_46_clock = clock;
  assign cores_46_reset = reset;
  assign cores_46_io_prev_valid = cores_45_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_46_io_prev_bits_address = cores_45_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_46_io_prev_bits_data = cores_45_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_46_io_prev_bits_wen = cores_45_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_46_io_prev_bits_id = cores_45_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_46_io_next_ready = cores_47_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_47_clock = clock;
  assign cores_47_reset = reset;
  assign cores_47_io_prev_valid = cores_46_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_47_io_prev_bits_address = cores_46_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_47_io_prev_bits_data = cores_46_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_47_io_prev_bits_wen = cores_46_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_47_io_prev_bits_id = cores_46_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_47_io_next_ready = cores_48_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_48_clock = clock;
  assign cores_48_reset = reset;
  assign cores_48_io_prev_valid = cores_47_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_48_io_prev_bits_address = cores_47_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_48_io_prev_bits_data = cores_47_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_48_io_prev_bits_wen = cores_47_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_48_io_prev_bits_id = cores_47_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_48_io_next_ready = cores_49_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_49_clock = clock;
  assign cores_49_reset = reset;
  assign cores_49_io_prev_valid = cores_48_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_49_io_prev_bits_address = cores_48_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_49_io_prev_bits_data = cores_48_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_49_io_prev_bits_wen = cores_48_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_49_io_prev_bits_id = cores_48_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_49_io_next_ready = cores_50_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_50_clock = clock;
  assign cores_50_reset = reset;
  assign cores_50_io_prev_valid = cores_49_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_50_io_prev_bits_address = cores_49_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_50_io_prev_bits_data = cores_49_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_50_io_prev_bits_wen = cores_49_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_50_io_prev_bits_id = cores_49_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_50_io_next_ready = cores_51_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_51_clock = clock;
  assign cores_51_reset = reset;
  assign cores_51_io_prev_valid = cores_50_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_51_io_prev_bits_address = cores_50_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_51_io_prev_bits_data = cores_50_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_51_io_prev_bits_wen = cores_50_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_51_io_prev_bits_id = cores_50_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_51_io_next_ready = cores_52_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_52_clock = clock;
  assign cores_52_reset = reset;
  assign cores_52_io_prev_valid = cores_51_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_52_io_prev_bits_address = cores_51_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_52_io_prev_bits_data = cores_51_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_52_io_prev_bits_wen = cores_51_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_52_io_prev_bits_id = cores_51_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_52_io_next_ready = cores_53_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_53_clock = clock;
  assign cores_53_reset = reset;
  assign cores_53_io_prev_valid = cores_52_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_53_io_prev_bits_address = cores_52_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_53_io_prev_bits_data = cores_52_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_53_io_prev_bits_wen = cores_52_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_53_io_prev_bits_id = cores_52_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_53_io_next_ready = cores_54_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_54_clock = clock;
  assign cores_54_reset = reset;
  assign cores_54_io_prev_valid = cores_53_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_54_io_prev_bits_address = cores_53_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_54_io_prev_bits_data = cores_53_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_54_io_prev_bits_wen = cores_53_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_54_io_prev_bits_id = cores_53_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_54_io_next_ready = cores_55_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_55_clock = clock;
  assign cores_55_reset = reset;
  assign cores_55_io_prev_valid = cores_54_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_55_io_prev_bits_address = cores_54_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_55_io_prev_bits_data = cores_54_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_55_io_prev_bits_wen = cores_54_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_55_io_prev_bits_id = cores_54_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_55_io_next_ready = cores_56_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_56_clock = clock;
  assign cores_56_reset = reset;
  assign cores_56_io_prev_valid = cores_55_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_56_io_prev_bits_address = cores_55_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_56_io_prev_bits_data = cores_55_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_56_io_prev_bits_wen = cores_55_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_56_io_prev_bits_id = cores_55_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_56_io_next_ready = cores_57_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_57_clock = clock;
  assign cores_57_reset = reset;
  assign cores_57_io_prev_valid = cores_56_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_57_io_prev_bits_address = cores_56_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_57_io_prev_bits_data = cores_56_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_57_io_prev_bits_wen = cores_56_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_57_io_prev_bits_id = cores_56_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_57_io_next_ready = cores_58_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_58_clock = clock;
  assign cores_58_reset = reset;
  assign cores_58_io_prev_valid = cores_57_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_58_io_prev_bits_address = cores_57_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_58_io_prev_bits_data = cores_57_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_58_io_prev_bits_wen = cores_57_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_58_io_prev_bits_id = cores_57_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_58_io_next_ready = cores_59_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_59_clock = clock;
  assign cores_59_reset = reset;
  assign cores_59_io_prev_valid = cores_58_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_59_io_prev_bits_address = cores_58_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_59_io_prev_bits_data = cores_58_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_59_io_prev_bits_wen = cores_58_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_59_io_prev_bits_id = cores_58_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_59_io_next_ready = cores_60_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_60_clock = clock;
  assign cores_60_reset = reset;
  assign cores_60_io_prev_valid = cores_59_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_60_io_prev_bits_address = cores_59_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_60_io_prev_bits_data = cores_59_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_60_io_prev_bits_wen = cores_59_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_60_io_prev_bits_id = cores_59_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_60_io_next_ready = cores_61_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_61_clock = clock;
  assign cores_61_reset = reset;
  assign cores_61_io_prev_valid = cores_60_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_61_io_prev_bits_address = cores_60_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_61_io_prev_bits_data = cores_60_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_61_io_prev_bits_wen = cores_60_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_61_io_prev_bits_id = cores_60_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_61_io_next_ready = cores_62_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_62_clock = clock;
  assign cores_62_reset = reset;
  assign cores_62_io_prev_valid = cores_61_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_62_io_prev_bits_address = cores_61_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_62_io_prev_bits_data = cores_61_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_62_io_prev_bits_wen = cores_61_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_62_io_prev_bits_id = cores_61_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_62_io_next_ready = cores_63_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_63_clock = clock;
  assign cores_63_reset = reset;
  assign cores_63_io_prev_valid = cores_62_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_63_io_prev_bits_address = cores_62_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_63_io_prev_bits_data = cores_62_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_63_io_prev_bits_wen = cores_62_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_63_io_prev_bits_id = cores_62_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_63_io_next_ready = cores_64_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_64_clock = clock;
  assign cores_64_reset = reset;
  assign cores_64_io_prev_valid = cores_63_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_64_io_prev_bits_address = cores_63_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_64_io_prev_bits_data = cores_63_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_64_io_prev_bits_wen = cores_63_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_64_io_prev_bits_id = cores_63_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_64_io_next_ready = cores_65_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_65_clock = clock;
  assign cores_65_reset = reset;
  assign cores_65_io_prev_valid = cores_64_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_65_io_prev_bits_address = cores_64_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_65_io_prev_bits_data = cores_64_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_65_io_prev_bits_wen = cores_64_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_65_io_prev_bits_id = cores_64_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_65_io_next_ready = cores_66_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_66_clock = clock;
  assign cores_66_reset = reset;
  assign cores_66_io_prev_valid = cores_65_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_66_io_prev_bits_address = cores_65_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_66_io_prev_bits_data = cores_65_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_66_io_prev_bits_wen = cores_65_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_66_io_prev_bits_id = cores_65_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_66_io_next_ready = cores_67_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_67_clock = clock;
  assign cores_67_reset = reset;
  assign cores_67_io_prev_valid = cores_66_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_67_io_prev_bits_address = cores_66_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_67_io_prev_bits_data = cores_66_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_67_io_prev_bits_wen = cores_66_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_67_io_prev_bits_id = cores_66_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_67_io_next_ready = cores_68_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_68_clock = clock;
  assign cores_68_reset = reset;
  assign cores_68_io_prev_valid = cores_67_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_68_io_prev_bits_address = cores_67_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_68_io_prev_bits_data = cores_67_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_68_io_prev_bits_wen = cores_67_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_68_io_prev_bits_id = cores_67_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_68_io_next_ready = cores_69_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_69_clock = clock;
  assign cores_69_reset = reset;
  assign cores_69_io_prev_valid = cores_68_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_69_io_prev_bits_address = cores_68_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_69_io_prev_bits_data = cores_68_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_69_io_prev_bits_wen = cores_68_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_69_io_prev_bits_id = cores_68_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_69_io_next_ready = cores_70_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_70_clock = clock;
  assign cores_70_reset = reset;
  assign cores_70_io_prev_valid = cores_69_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_70_io_prev_bits_address = cores_69_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_70_io_prev_bits_data = cores_69_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_70_io_prev_bits_wen = cores_69_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_70_io_prev_bits_id = cores_69_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_70_io_next_ready = cores_71_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_71_clock = clock;
  assign cores_71_reset = reset;
  assign cores_71_io_prev_valid = cores_70_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_71_io_prev_bits_address = cores_70_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_71_io_prev_bits_data = cores_70_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_71_io_prev_bits_wen = cores_70_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_71_io_prev_bits_id = cores_70_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_71_io_next_ready = cores_72_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_72_clock = clock;
  assign cores_72_reset = reset;
  assign cores_72_io_prev_valid = cores_71_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_72_io_prev_bits_address = cores_71_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_72_io_prev_bits_data = cores_71_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_72_io_prev_bits_wen = cores_71_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_72_io_prev_bits_id = cores_71_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_72_io_next_ready = cores_73_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_73_clock = clock;
  assign cores_73_reset = reset;
  assign cores_73_io_prev_valid = cores_72_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_73_io_prev_bits_address = cores_72_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_73_io_prev_bits_data = cores_72_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_73_io_prev_bits_wen = cores_72_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_73_io_prev_bits_id = cores_72_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_73_io_next_ready = cores_74_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_74_clock = clock;
  assign cores_74_reset = reset;
  assign cores_74_io_prev_valid = cores_73_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_74_io_prev_bits_address = cores_73_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_74_io_prev_bits_data = cores_73_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_74_io_prev_bits_wen = cores_73_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_74_io_prev_bits_id = cores_73_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_74_io_next_ready = cores_75_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_75_clock = clock;
  assign cores_75_reset = reset;
  assign cores_75_io_prev_valid = cores_74_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_75_io_prev_bits_address = cores_74_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_75_io_prev_bits_data = cores_74_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_75_io_prev_bits_wen = cores_74_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_75_io_prev_bits_id = cores_74_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_75_io_next_ready = cores_76_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_76_clock = clock;
  assign cores_76_reset = reset;
  assign cores_76_io_prev_valid = cores_75_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_76_io_prev_bits_address = cores_75_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_76_io_prev_bits_data = cores_75_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_76_io_prev_bits_wen = cores_75_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_76_io_prev_bits_id = cores_75_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_76_io_next_ready = cores_77_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_77_clock = clock;
  assign cores_77_reset = reset;
  assign cores_77_io_prev_valid = cores_76_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_77_io_prev_bits_address = cores_76_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_77_io_prev_bits_data = cores_76_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_77_io_prev_bits_wen = cores_76_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_77_io_prev_bits_id = cores_76_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_77_io_next_ready = cores_78_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_78_clock = clock;
  assign cores_78_reset = reset;
  assign cores_78_io_prev_valid = cores_77_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_78_io_prev_bits_address = cores_77_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_78_io_prev_bits_data = cores_77_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_78_io_prev_bits_wen = cores_77_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_78_io_prev_bits_id = cores_77_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_78_io_next_ready = cores_79_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_79_clock = clock;
  assign cores_79_reset = reset;
  assign cores_79_io_prev_valid = cores_78_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_79_io_prev_bits_address = cores_78_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_79_io_prev_bits_data = cores_78_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_79_io_prev_bits_wen = cores_78_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_79_io_prev_bits_id = cores_78_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_79_io_next_ready = cores_80_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_80_clock = clock;
  assign cores_80_reset = reset;
  assign cores_80_io_prev_valid = cores_79_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_80_io_prev_bits_address = cores_79_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_80_io_prev_bits_data = cores_79_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_80_io_prev_bits_wen = cores_79_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_80_io_prev_bits_id = cores_79_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_80_io_next_ready = cores_81_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_81_clock = clock;
  assign cores_81_reset = reset;
  assign cores_81_io_prev_valid = cores_80_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_81_io_prev_bits_address = cores_80_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_81_io_prev_bits_data = cores_80_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_81_io_prev_bits_wen = cores_80_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_81_io_prev_bits_id = cores_80_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_81_io_next_ready = cores_82_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_82_clock = clock;
  assign cores_82_reset = reset;
  assign cores_82_io_prev_valid = cores_81_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_82_io_prev_bits_address = cores_81_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_82_io_prev_bits_data = cores_81_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_82_io_prev_bits_wen = cores_81_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_82_io_prev_bits_id = cores_81_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_82_io_next_ready = cores_83_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_83_clock = clock;
  assign cores_83_reset = reset;
  assign cores_83_io_prev_valid = cores_82_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_83_io_prev_bits_address = cores_82_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_83_io_prev_bits_data = cores_82_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_83_io_prev_bits_wen = cores_82_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_83_io_prev_bits_id = cores_82_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_83_io_next_ready = cores_84_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_84_clock = clock;
  assign cores_84_reset = reset;
  assign cores_84_io_prev_valid = cores_83_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_84_io_prev_bits_address = cores_83_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_84_io_prev_bits_data = cores_83_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_84_io_prev_bits_wen = cores_83_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_84_io_prev_bits_id = cores_83_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_84_io_next_ready = cores_85_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_85_clock = clock;
  assign cores_85_reset = reset;
  assign cores_85_io_prev_valid = cores_84_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_85_io_prev_bits_address = cores_84_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_85_io_prev_bits_data = cores_84_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_85_io_prev_bits_wen = cores_84_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_85_io_prev_bits_id = cores_84_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_85_io_next_ready = cores_86_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_86_clock = clock;
  assign cores_86_reset = reset;
  assign cores_86_io_prev_valid = cores_85_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_86_io_prev_bits_address = cores_85_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_86_io_prev_bits_data = cores_85_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_86_io_prev_bits_wen = cores_85_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_86_io_prev_bits_id = cores_85_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_86_io_next_ready = cores_87_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_87_clock = clock;
  assign cores_87_reset = reset;
  assign cores_87_io_prev_valid = cores_86_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_87_io_prev_bits_address = cores_86_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_87_io_prev_bits_data = cores_86_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_87_io_prev_bits_wen = cores_86_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_87_io_prev_bits_id = cores_86_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_87_io_next_ready = cores_88_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_88_clock = clock;
  assign cores_88_reset = reset;
  assign cores_88_io_prev_valid = cores_87_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_88_io_prev_bits_address = cores_87_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_88_io_prev_bits_data = cores_87_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_88_io_prev_bits_wen = cores_87_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_88_io_prev_bits_id = cores_87_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_88_io_next_ready = cores_89_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_89_clock = clock;
  assign cores_89_reset = reset;
  assign cores_89_io_prev_valid = cores_88_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_89_io_prev_bits_address = cores_88_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_89_io_prev_bits_data = cores_88_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_89_io_prev_bits_wen = cores_88_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_89_io_prev_bits_id = cores_88_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_89_io_next_ready = cores_90_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_90_clock = clock;
  assign cores_90_reset = reset;
  assign cores_90_io_prev_valid = cores_89_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_90_io_prev_bits_address = cores_89_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_90_io_prev_bits_data = cores_89_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_90_io_prev_bits_wen = cores_89_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_90_io_prev_bits_id = cores_89_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_90_io_next_ready = cores_91_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_91_clock = clock;
  assign cores_91_reset = reset;
  assign cores_91_io_prev_valid = cores_90_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_91_io_prev_bits_address = cores_90_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_91_io_prev_bits_data = cores_90_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_91_io_prev_bits_wen = cores_90_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_91_io_prev_bits_id = cores_90_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_91_io_next_ready = cores_92_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_92_clock = clock;
  assign cores_92_reset = reset;
  assign cores_92_io_prev_valid = cores_91_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_92_io_prev_bits_address = cores_91_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_92_io_prev_bits_data = cores_91_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_92_io_prev_bits_wen = cores_91_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_92_io_prev_bits_id = cores_91_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_92_io_next_ready = cores_93_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_93_clock = clock;
  assign cores_93_reset = reset;
  assign cores_93_io_prev_valid = cores_92_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_93_io_prev_bits_address = cores_92_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_93_io_prev_bits_data = cores_92_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_93_io_prev_bits_wen = cores_92_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_93_io_prev_bits_id = cores_92_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_93_io_next_ready = cores_94_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_94_clock = clock;
  assign cores_94_reset = reset;
  assign cores_94_io_prev_valid = cores_93_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_94_io_prev_bits_address = cores_93_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_94_io_prev_bits_data = cores_93_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_94_io_prev_bits_wen = cores_93_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_94_io_prev_bits_id = cores_93_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_94_io_next_ready = cores_95_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_95_clock = clock;
  assign cores_95_reset = reset;
  assign cores_95_io_prev_valid = cores_94_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_95_io_prev_bits_address = cores_94_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_95_io_prev_bits_data = cores_94_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_95_io_prev_bits_wen = cores_94_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_95_io_prev_bits_id = cores_94_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_95_io_next_ready = cores_96_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_96_clock = clock;
  assign cores_96_reset = reset;
  assign cores_96_io_prev_valid = cores_95_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_96_io_prev_bits_address = cores_95_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_96_io_prev_bits_data = cores_95_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_96_io_prev_bits_wen = cores_95_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_96_io_prev_bits_id = cores_95_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_96_io_next_ready = cores_97_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_97_clock = clock;
  assign cores_97_reset = reset;
  assign cores_97_io_prev_valid = cores_96_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_97_io_prev_bits_address = cores_96_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_97_io_prev_bits_data = cores_96_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_97_io_prev_bits_wen = cores_96_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_97_io_prev_bits_id = cores_96_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_97_io_next_ready = cores_98_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_98_clock = clock;
  assign cores_98_reset = reset;
  assign cores_98_io_prev_valid = cores_97_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_98_io_prev_bits_address = cores_97_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_98_io_prev_bits_data = cores_97_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_98_io_prev_bits_wen = cores_97_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_98_io_prev_bits_id = cores_97_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_98_io_next_ready = cores_99_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_99_clock = clock;
  assign cores_99_reset = reset;
  assign cores_99_io_prev_valid = cores_98_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_99_io_prev_bits_address = cores_98_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_99_io_prev_bits_data = cores_98_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_99_io_prev_bits_wen = cores_98_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_99_io_prev_bits_id = cores_98_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_99_io_next_ready = cores_100_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_100_clock = clock;
  assign cores_100_reset = reset;
  assign cores_100_io_prev_valid = cores_99_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_100_io_prev_bits_address = cores_99_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_100_io_prev_bits_data = cores_99_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_100_io_prev_bits_wen = cores_99_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_100_io_prev_bits_id = cores_99_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_100_io_next_ready = cores_101_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_101_clock = clock;
  assign cores_101_reset = reset;
  assign cores_101_io_prev_valid = cores_100_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_101_io_prev_bits_address = cores_100_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_101_io_prev_bits_data = cores_100_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_101_io_prev_bits_wen = cores_100_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_101_io_prev_bits_id = cores_100_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_101_io_next_ready = cores_102_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_102_clock = clock;
  assign cores_102_reset = reset;
  assign cores_102_io_prev_valid = cores_101_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_102_io_prev_bits_address = cores_101_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_102_io_prev_bits_data = cores_101_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_102_io_prev_bits_wen = cores_101_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_102_io_prev_bits_id = cores_101_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_102_io_next_ready = cores_103_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_103_clock = clock;
  assign cores_103_reset = reset;
  assign cores_103_io_prev_valid = cores_102_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_103_io_prev_bits_address = cores_102_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_103_io_prev_bits_data = cores_102_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_103_io_prev_bits_wen = cores_102_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_103_io_prev_bits_id = cores_102_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_103_io_next_ready = cores_104_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_104_clock = clock;
  assign cores_104_reset = reset;
  assign cores_104_io_prev_valid = cores_103_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_104_io_prev_bits_address = cores_103_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_104_io_prev_bits_data = cores_103_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_104_io_prev_bits_wen = cores_103_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_104_io_prev_bits_id = cores_103_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_104_io_next_ready = cores_105_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_105_clock = clock;
  assign cores_105_reset = reset;
  assign cores_105_io_prev_valid = cores_104_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_105_io_prev_bits_address = cores_104_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_105_io_prev_bits_data = cores_104_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_105_io_prev_bits_wen = cores_104_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_105_io_prev_bits_id = cores_104_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_105_io_next_ready = cores_106_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_106_clock = clock;
  assign cores_106_reset = reset;
  assign cores_106_io_prev_valid = cores_105_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_106_io_prev_bits_address = cores_105_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_106_io_prev_bits_data = cores_105_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_106_io_prev_bits_wen = cores_105_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_106_io_prev_bits_id = cores_105_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_106_io_next_ready = cores_107_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_107_clock = clock;
  assign cores_107_reset = reset;
  assign cores_107_io_prev_valid = cores_106_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_107_io_prev_bits_address = cores_106_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_107_io_prev_bits_data = cores_106_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_107_io_prev_bits_wen = cores_106_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_107_io_prev_bits_id = cores_106_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_107_io_next_ready = cores_108_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_108_clock = clock;
  assign cores_108_reset = reset;
  assign cores_108_io_prev_valid = cores_107_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_108_io_prev_bits_address = cores_107_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_108_io_prev_bits_data = cores_107_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_108_io_prev_bits_wen = cores_107_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_108_io_prev_bits_id = cores_107_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_108_io_next_ready = cores_109_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_109_clock = clock;
  assign cores_109_reset = reset;
  assign cores_109_io_prev_valid = cores_108_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_109_io_prev_bits_address = cores_108_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_109_io_prev_bits_data = cores_108_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_109_io_prev_bits_wen = cores_108_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_109_io_prev_bits_id = cores_108_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_109_io_next_ready = cores_110_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_110_clock = clock;
  assign cores_110_reset = reset;
  assign cores_110_io_prev_valid = cores_109_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_110_io_prev_bits_address = cores_109_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_110_io_prev_bits_data = cores_109_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_110_io_prev_bits_wen = cores_109_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_110_io_prev_bits_id = cores_109_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_110_io_next_ready = cores_111_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_111_clock = clock;
  assign cores_111_reset = reset;
  assign cores_111_io_prev_valid = cores_110_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_111_io_prev_bits_address = cores_110_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_111_io_prev_bits_data = cores_110_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_111_io_prev_bits_wen = cores_110_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_111_io_prev_bits_id = cores_110_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_111_io_next_ready = cores_112_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_112_clock = clock;
  assign cores_112_reset = reset;
  assign cores_112_io_prev_valid = cores_111_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_112_io_prev_bits_address = cores_111_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_112_io_prev_bits_data = cores_111_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_112_io_prev_bits_wen = cores_111_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_112_io_prev_bits_id = cores_111_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_112_io_next_ready = cores_113_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_113_clock = clock;
  assign cores_113_reset = reset;
  assign cores_113_io_prev_valid = cores_112_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_113_io_prev_bits_address = cores_112_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_113_io_prev_bits_data = cores_112_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_113_io_prev_bits_wen = cores_112_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_113_io_prev_bits_id = cores_112_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_113_io_next_ready = cores_114_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_114_clock = clock;
  assign cores_114_reset = reset;
  assign cores_114_io_prev_valid = cores_113_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_114_io_prev_bits_address = cores_113_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_114_io_prev_bits_data = cores_113_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_114_io_prev_bits_wen = cores_113_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_114_io_prev_bits_id = cores_113_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_114_io_next_ready = cores_115_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_115_clock = clock;
  assign cores_115_reset = reset;
  assign cores_115_io_prev_valid = cores_114_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_115_io_prev_bits_address = cores_114_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_115_io_prev_bits_data = cores_114_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_115_io_prev_bits_wen = cores_114_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_115_io_prev_bits_id = cores_114_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_115_io_next_ready = cores_116_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_116_clock = clock;
  assign cores_116_reset = reset;
  assign cores_116_io_prev_valid = cores_115_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_116_io_prev_bits_address = cores_115_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_116_io_prev_bits_data = cores_115_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_116_io_prev_bits_wen = cores_115_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_116_io_prev_bits_id = cores_115_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_116_io_next_ready = cores_117_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_117_clock = clock;
  assign cores_117_reset = reset;
  assign cores_117_io_prev_valid = cores_116_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_117_io_prev_bits_address = cores_116_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_117_io_prev_bits_data = cores_116_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_117_io_prev_bits_wen = cores_116_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_117_io_prev_bits_id = cores_116_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_117_io_next_ready = cores_118_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_118_clock = clock;
  assign cores_118_reset = reset;
  assign cores_118_io_prev_valid = cores_117_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_118_io_prev_bits_address = cores_117_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_118_io_prev_bits_data = cores_117_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_118_io_prev_bits_wen = cores_117_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_118_io_prev_bits_id = cores_117_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_118_io_next_ready = cores_119_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_119_clock = clock;
  assign cores_119_reset = reset;
  assign cores_119_io_prev_valid = cores_118_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_119_io_prev_bits_address = cores_118_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_119_io_prev_bits_data = cores_118_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_119_io_prev_bits_wen = cores_118_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_119_io_prev_bits_id = cores_118_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_119_io_next_ready = cores_120_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_120_clock = clock;
  assign cores_120_reset = reset;
  assign cores_120_io_prev_valid = cores_119_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_120_io_prev_bits_address = cores_119_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_120_io_prev_bits_data = cores_119_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_120_io_prev_bits_wen = cores_119_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_120_io_prev_bits_id = cores_119_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_120_io_next_ready = cores_121_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_121_clock = clock;
  assign cores_121_reset = reset;
  assign cores_121_io_prev_valid = cores_120_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_121_io_prev_bits_address = cores_120_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_121_io_prev_bits_data = cores_120_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_121_io_prev_bits_wen = cores_120_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_121_io_prev_bits_id = cores_120_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_121_io_next_ready = cores_122_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_122_clock = clock;
  assign cores_122_reset = reset;
  assign cores_122_io_prev_valid = cores_121_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_122_io_prev_bits_address = cores_121_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_122_io_prev_bits_data = cores_121_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_122_io_prev_bits_wen = cores_121_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_122_io_prev_bits_id = cores_121_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_122_io_next_ready = cores_123_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_123_clock = clock;
  assign cores_123_reset = reset;
  assign cores_123_io_prev_valid = cores_122_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_123_io_prev_bits_address = cores_122_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_123_io_prev_bits_data = cores_122_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_123_io_prev_bits_wen = cores_122_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_123_io_prev_bits_id = cores_122_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_123_io_next_ready = cores_124_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_124_clock = clock;
  assign cores_124_reset = reset;
  assign cores_124_io_prev_valid = cores_123_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_124_io_prev_bits_address = cores_123_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_124_io_prev_bits_data = cores_123_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_124_io_prev_bits_wen = cores_123_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_124_io_prev_bits_id = cores_123_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_124_io_next_ready = cores_125_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_125_clock = clock;
  assign cores_125_reset = reset;
  assign cores_125_io_prev_valid = cores_124_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_125_io_prev_bits_address = cores_124_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_125_io_prev_bits_data = cores_124_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_125_io_prev_bits_wen = cores_124_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_125_io_prev_bits_id = cores_124_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_125_io_next_ready = cores_126_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_126_clock = clock;
  assign cores_126_reset = reset;
  assign cores_126_io_prev_valid = cores_125_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_126_io_prev_bits_address = cores_125_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_126_io_prev_bits_data = cores_125_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_126_io_prev_bits_wen = cores_125_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_126_io_prev_bits_id = cores_125_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_126_io_next_ready = cores_127_io_prev_ready; // @[FemtoMips32.scala 473:21]
  assign cores_127_clock = clock;
  assign cores_127_reset = reset;
  assign cores_127_io_prev_valid = cores_126_io_next_valid; // @[FemtoMips32.scala 473:21]
  assign cores_127_io_prev_bits_address = cores_126_io_next_bits_address; // @[FemtoMips32.scala 473:21]
  assign cores_127_io_prev_bits_data = cores_126_io_next_bits_data; // @[FemtoMips32.scala 473:21]
  assign cores_127_io_prev_bits_wen = cores_126_io_next_bits_wen; // @[FemtoMips32.scala 473:21]
  assign cores_127_io_prev_bits_id = cores_126_io_next_bits_id; // @[FemtoMips32.scala 473:21]
  assign cores_127_io_next_ready = io_next_ready; // @[FemtoMips32.scala 478:22]
endmodule
